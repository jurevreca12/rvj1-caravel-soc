magic
tech sky130A
magscale 1 2
timestamp 1653848533
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 219342 700408 219348 700460
rect 219400 700448 219406 700460
rect 267642 700448 267648 700460
rect 219400 700420 267648 700448
rect 219400 700408 219406 700420
rect 267642 700408 267648 700420
rect 267700 700408 267706 700460
rect 8110 700340 8116 700392
rect 8168 700380 8174 700392
rect 13078 700380 13084 700392
rect 8168 700352 13084 700380
rect 8168 700340 8174 700352
rect 13078 700340 13084 700352
rect 13136 700340 13142 700392
rect 137830 700340 137836 700392
rect 137888 700380 137894 700392
rect 138658 700380 138664 700392
rect 137888 700352 138664 700380
rect 137888 700340 137894 700352
rect 138658 700340 138664 700352
rect 138716 700340 138722 700392
rect 217962 700340 217968 700392
rect 218020 700380 218026 700392
rect 283834 700380 283840 700392
rect 218020 700352 283840 700380
rect 218020 700340 218026 700352
rect 283834 700340 283840 700352
rect 283892 700340 283898 700392
rect 348786 700340 348792 700392
rect 348844 700380 348850 700392
rect 357434 700380 357440 700392
rect 348844 700352 357440 700380
rect 348844 700340 348850 700352
rect 357434 700340 357440 700352
rect 357492 700340 357498 700392
rect 105446 700272 105452 700324
rect 105504 700312 105510 700324
rect 206278 700312 206284 700324
rect 105504 700284 206284 700312
rect 105504 700272 105510 700284
rect 206278 700272 206284 700284
rect 206336 700272 206342 700324
rect 219250 700272 219256 700324
rect 219308 700312 219314 700324
rect 300118 700312 300124 700324
rect 219308 700284 300124 700312
rect 219308 700272 219314 700284
rect 300118 700272 300124 700284
rect 300176 700272 300182 700324
rect 332502 700272 332508 700324
rect 332560 700312 332566 700324
rect 358814 700312 358820 700324
rect 332560 700284 358820 700312
rect 332560 700272 332566 700284
rect 358814 700272 358820 700284
rect 358872 700272 358878 700324
rect 367738 700272 367744 700324
rect 367796 700312 367802 700324
rect 559650 700312 559656 700324
rect 367796 700284 559656 700312
rect 367796 700272 367802 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 25498 699700 25504 699712
rect 24360 699672 25504 699700
rect 24360 699660 24366 699672
rect 25498 699660 25504 699672
rect 25556 699660 25562 699712
rect 396718 699660 396724 699712
rect 396776 699700 396782 699712
rect 397454 699700 397460 699712
rect 396776 699672 397460 699700
rect 396776 699660 396782 699672
rect 397454 699660 397460 699672
rect 397512 699660 397518 699712
rect 428458 699660 428464 699712
rect 428516 699700 428522 699712
rect 429838 699700 429844 699712
rect 428516 699672 429844 699700
rect 428516 699660 428522 699672
rect 429838 699660 429844 699672
rect 429896 699660 429902 699712
rect 371878 696940 371884 696992
rect 371936 696980 371942 696992
rect 580166 696980 580172 696992
rect 371936 696952 580172 696980
rect 371936 696940 371942 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 10318 683176 10324 683188
rect 3476 683148 10324 683176
rect 3476 683136 3482 683148
rect 10318 683136 10324 683148
rect 10376 683136 10382 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 180058 670732 180064 670744
rect 3568 670704 180064 670732
rect 3568 670692 3574 670704
rect 180058 670692 180064 670704
rect 180116 670692 180122 670744
rect 360838 670692 360844 670744
rect 360896 670732 360902 670744
rect 580166 670732 580172 670744
rect 360896 670704 580172 670732
rect 360896 670692 360902 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 14458 656928 14464 656940
rect 3476 656900 14464 656928
rect 3476 656888 3482 656900
rect 14458 656888 14464 656900
rect 14516 656888 14522 656940
rect 369118 643084 369124 643136
rect 369176 643124 369182 643136
rect 580166 643124 580172 643136
rect 369176 643096 580172 643124
rect 369176 643084 369182 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 8938 632108 8944 632120
rect 3476 632080 8944 632108
rect 3476 632068 3482 632080
rect 8938 632068 8944 632080
rect 8996 632068 9002 632120
rect 377398 630640 377404 630692
rect 377456 630680 377462 630692
rect 579982 630680 579988 630692
rect 377456 630652 579988 630680
rect 377456 630640 377462 630652
rect 579982 630640 579988 630652
rect 580040 630640 580046 630692
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 182818 618304 182824 618316
rect 3200 618276 182824 618304
rect 3200 618264 3206 618276
rect 182818 618264 182824 618276
rect 182876 618264 182882 618316
rect 432598 616836 432604 616888
rect 432656 616876 432662 616888
rect 580166 616876 580172 616888
rect 432656 616848 580172 616876
rect 432656 616836 432662 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3418 606024 3424 606076
rect 3476 606064 3482 606076
rect 7558 606064 7564 606076
rect 3476 606036 7564 606064
rect 3476 606024 3482 606036
rect 7558 606024 7564 606036
rect 7616 606024 7622 606076
rect 363598 590656 363604 590708
rect 363656 590696 363662 590708
rect 580166 590696 580172 590708
rect 363656 590668 580172 590696
rect 363656 590656 363662 590668
rect 580166 590656 580172 590668
rect 580224 590656 580230 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 32398 579680 32404 579692
rect 3384 579652 32404 579680
rect 3384 579640 3390 579652
rect 32398 579640 32404 579652
rect 32456 579640 32462 579692
rect 373258 576852 373264 576904
rect 373316 576892 373322 576904
rect 580166 576892 580172 576904
rect 373316 576864 580172 576892
rect 373316 576852 373322 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 21358 565876 21364 565888
rect 3476 565848 21364 565876
rect 3476 565836 3482 565848
rect 21358 565836 21364 565848
rect 21416 565836 21422 565888
rect 217870 565088 217876 565140
rect 217928 565128 217934 565140
rect 234614 565128 234620 565140
rect 217928 565100 234620 565128
rect 217928 565088 217934 565100
rect 234614 565088 234620 565100
rect 234672 565088 234678 565140
rect 359458 563048 359464 563100
rect 359516 563088 359522 563100
rect 580166 563088 580172 563100
rect 359516 563060 580172 563088
rect 359516 563048 359522 563060
rect 580166 563048 580172 563060
rect 580224 563048 580230 563100
rect 3418 553392 3424 553444
rect 3476 553432 3482 553444
rect 17218 553432 17224 553444
rect 3476 553404 17224 553432
rect 3476 553392 3482 553404
rect 17218 553392 17224 553404
rect 17276 553392 17282 553444
rect 576118 536800 576124 536852
rect 576176 536840 576182 536852
rect 579890 536840 579896 536852
rect 576176 536812 579896 536840
rect 576176 536800 576182 536812
rect 579890 536800 579896 536812
rect 579948 536800 579954 536852
rect 2774 527144 2780 527196
rect 2832 527184 2838 527196
rect 4798 527184 4804 527196
rect 2832 527156 4804 527184
rect 2832 527144 2838 527156
rect 4798 527144 4804 527156
rect 4856 527144 4862 527196
rect 570598 524424 570604 524476
rect 570656 524464 570662 524476
rect 580166 524464 580172 524476
rect 570656 524436 580172 524464
rect 570656 524424 570662 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 18598 501004 18604 501016
rect 3108 500976 18604 501004
rect 3108 500964 3114 500976
rect 18598 500964 18604 500976
rect 18656 500964 18662 501016
rect 574738 484372 574744 484424
rect 574796 484412 574802 484424
rect 580166 484412 580172 484424
rect 574796 484384 580172 484412
rect 574796 484372 574802 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 219250 478524 219256 478576
rect 219308 478564 219314 478576
rect 266446 478564 266452 478576
rect 219308 478536 266452 478564
rect 219308 478524 219314 478536
rect 266446 478524 266452 478536
rect 266504 478524 266510 478576
rect 217962 478456 217968 478508
rect 218020 478496 218026 478508
rect 267734 478496 267740 478508
rect 218020 478468 267740 478496
rect 218020 478456 218026 478468
rect 267734 478456 267740 478468
rect 267792 478456 267798 478508
rect 217410 478388 217416 478440
rect 217468 478428 217474 478440
rect 302234 478428 302240 478440
rect 217468 478400 302240 478428
rect 217468 478388 217474 478400
rect 302234 478388 302240 478400
rect 302292 478388 302298 478440
rect 266354 478320 266360 478372
rect 266412 478360 266418 478372
rect 357434 478360 357440 478372
rect 266412 478332 357440 478360
rect 266412 478320 266418 478332
rect 357434 478320 357440 478332
rect 357492 478320 357498 478372
rect 218882 478252 218888 478304
rect 218940 478292 218946 478304
rect 310514 478292 310520 478304
rect 218940 478264 310520 478292
rect 218940 478252 218946 478264
rect 310514 478252 310520 478264
rect 310572 478252 310578 478304
rect 264974 478184 264980 478236
rect 265032 478224 265038 478236
rect 358814 478224 358820 478236
rect 265032 478196 358820 478224
rect 265032 478184 265038 478196
rect 358814 478184 358820 478196
rect 358872 478184 358878 478236
rect 18598 478116 18604 478168
rect 18656 478156 18662 478168
rect 281534 478156 281540 478168
rect 18656 478128 281540 478156
rect 18656 478116 18662 478128
rect 281534 478116 281540 478128
rect 281592 478116 281598 478168
rect 241422 476756 241428 476808
rect 241480 476796 241486 476808
rect 309134 476796 309140 476808
rect 241480 476768 309140 476796
rect 241480 476756 241486 476768
rect 309134 476756 309140 476768
rect 309192 476756 309198 476808
rect 242802 476688 242808 476740
rect 242860 476728 242866 476740
rect 311894 476728 311900 476740
rect 242860 476700 311900 476728
rect 242860 476688 242866 476700
rect 311894 476688 311900 476700
rect 311952 476688 311958 476740
rect 238478 476620 238484 476672
rect 238536 476660 238542 476672
rect 304994 476660 305000 476672
rect 238536 476632 305000 476660
rect 238536 476620 238542 476632
rect 304994 476620 305000 476632
rect 305052 476620 305058 476672
rect 306098 476620 306104 476672
rect 306156 476660 306162 476672
rect 322198 476660 322204 476672
rect 306156 476632 322204 476660
rect 306156 476620 306162 476632
rect 322198 476620 322204 476632
rect 322256 476620 322262 476672
rect 264882 476552 264888 476604
rect 264940 476592 264946 476604
rect 317414 476592 317420 476604
rect 264940 476564 317420 476592
rect 264940 476552 264946 476564
rect 317414 476552 317420 476564
rect 317472 476552 317478 476604
rect 269022 476484 269028 476536
rect 269080 476524 269086 476536
rect 321554 476524 321560 476536
rect 269080 476496 321560 476524
rect 269080 476484 269086 476496
rect 321554 476484 321560 476496
rect 321612 476484 321618 476536
rect 259362 476416 259368 476468
rect 259420 476456 259426 476468
rect 314654 476456 314660 476468
rect 259420 476428 314660 476456
rect 259420 476416 259426 476428
rect 314654 476416 314660 476428
rect 314712 476416 314718 476468
rect 253842 476348 253848 476400
rect 253900 476388 253906 476400
rect 309226 476388 309232 476400
rect 253900 476360 309232 476388
rect 253900 476348 253906 476360
rect 309226 476348 309232 476360
rect 309284 476348 309290 476400
rect 318702 476348 318708 476400
rect 318760 476388 318766 476400
rect 327718 476388 327724 476400
rect 318760 476360 327724 476388
rect 318760 476348 318766 476360
rect 327718 476348 327724 476360
rect 327776 476348 327782 476400
rect 303522 476280 303528 476332
rect 303580 476320 303586 476332
rect 320818 476320 320824 476332
rect 303580 476292 320824 476320
rect 303580 476280 303586 476292
rect 320818 476280 320824 476292
rect 320876 476280 320882 476332
rect 321462 476280 321468 476332
rect 321520 476320 321526 476332
rect 329098 476320 329104 476332
rect 321520 476292 329104 476320
rect 321520 476280 321526 476292
rect 329098 476280 329104 476292
rect 329156 476280 329162 476332
rect 309042 476212 309048 476264
rect 309100 476252 309106 476264
rect 323578 476252 323584 476264
rect 309100 476224 323584 476252
rect 309100 476212 309106 476224
rect 323578 476212 323584 476224
rect 323636 476212 323642 476264
rect 324222 476212 324228 476264
rect 324280 476252 324286 476264
rect 338758 476252 338764 476264
rect 324280 476224 338764 476252
rect 324280 476212 324286 476224
rect 338758 476212 338764 476224
rect 338816 476212 338822 476264
rect 240042 476144 240048 476196
rect 240100 476184 240106 476196
rect 307754 476184 307760 476196
rect 240100 476156 307760 476184
rect 240100 476144 240106 476156
rect 307754 476144 307760 476156
rect 307812 476144 307818 476196
rect 311802 476076 311808 476128
rect 311860 476116 311866 476128
rect 324958 476116 324964 476128
rect 311860 476088 324964 476116
rect 311860 476076 311866 476088
rect 324958 476076 324964 476088
rect 325016 476076 325022 476128
rect 326982 476076 326988 476128
rect 327040 476116 327046 476128
rect 331858 476116 331864 476128
rect 327040 476088 331864 476116
rect 327040 476076 327046 476088
rect 331858 476076 331864 476088
rect 331916 476076 331922 476128
rect 302142 475532 302148 475584
rect 302200 475572 302206 475584
rect 336734 475572 336740 475584
rect 302200 475544 336740 475572
rect 302200 475532 302206 475544
rect 336734 475532 336740 475544
rect 336792 475532 336798 475584
rect 281442 475464 281448 475516
rect 281500 475504 281506 475516
rect 327074 475504 327080 475516
rect 281500 475476 327080 475504
rect 281500 475464 281506 475476
rect 327074 475464 327080 475476
rect 327132 475464 327138 475516
rect 237282 475396 237288 475448
rect 237340 475436 237346 475448
rect 305086 475436 305092 475448
rect 237340 475408 305092 475436
rect 237340 475396 237346 475408
rect 305086 475396 305092 475408
rect 305144 475396 305150 475448
rect 217594 475328 217600 475380
rect 217652 475368 217658 475380
rect 316126 475368 316132 475380
rect 217652 475340 316132 475368
rect 217652 475328 217658 475340
rect 316126 475328 316132 475340
rect 316184 475328 316190 475380
rect 3418 474716 3424 474768
rect 3476 474756 3482 474768
rect 282914 474756 282920 474768
rect 3476 474728 282920 474756
rect 3476 474716 3482 474728
rect 282914 474716 282920 474728
rect 282972 474716 282978 474768
rect 274542 474172 274548 474224
rect 274600 474212 274606 474224
rect 324314 474212 324320 474224
rect 274600 474184 324320 474212
rect 274600 474172 274606 474184
rect 324314 474172 324320 474184
rect 324372 474172 324378 474224
rect 237374 474104 237380 474156
rect 237432 474144 237438 474156
rect 303614 474144 303620 474156
rect 237432 474116 303620 474144
rect 237432 474104 237438 474116
rect 303614 474104 303620 474116
rect 303672 474104 303678 474156
rect 255222 474036 255228 474088
rect 255280 474076 255286 474088
rect 323026 474076 323032 474088
rect 255280 474048 323032 474076
rect 255280 474036 255286 474048
rect 323026 474036 323032 474048
rect 323084 474036 323090 474088
rect 17218 473968 17224 474020
rect 17276 474008 17282 474020
rect 280154 474008 280160 474020
rect 17276 473980 280160 474008
rect 17276 473968 17282 473980
rect 280154 473968 280160 473980
rect 280212 473968 280218 474020
rect 314562 473968 314568 474020
rect 314620 474008 314626 474020
rect 343634 474008 343640 474020
rect 314620 473980 343640 474008
rect 314620 473968 314626 473980
rect 343634 473968 343640 473980
rect 343692 473968 343698 474020
rect 252370 472744 252376 472796
rect 252428 472784 252434 472796
rect 318794 472784 318800 472796
rect 252428 472756 318800 472784
rect 252428 472744 252434 472756
rect 318794 472744 318800 472756
rect 318852 472744 318858 472796
rect 218974 472676 218980 472728
rect 219032 472716 219038 472728
rect 307846 472716 307852 472728
rect 219032 472688 307852 472716
rect 219032 472676 219038 472688
rect 307846 472676 307852 472688
rect 307904 472676 307910 472728
rect 315942 472676 315948 472728
rect 316000 472716 316006 472728
rect 345198 472716 345204 472728
rect 316000 472688 345204 472716
rect 316000 472676 316006 472688
rect 345198 472676 345204 472688
rect 345256 472676 345262 472728
rect 255314 472608 255320 472660
rect 255372 472648 255378 472660
rect 373258 472648 373264 472660
rect 255372 472620 373264 472648
rect 255372 472608 255378 472620
rect 373258 472608 373264 472620
rect 373316 472608 373322 472660
rect 217502 471316 217508 471368
rect 217560 471356 217566 471368
rect 300854 471356 300860 471368
rect 217560 471328 300860 471356
rect 217560 471316 217566 471328
rect 300854 471316 300860 471328
rect 300912 471316 300918 471368
rect 3510 471248 3516 471300
rect 3568 471288 3574 471300
rect 283006 471288 283012 471300
rect 3568 471260 283012 471288
rect 3568 471248 3574 471260
rect 283006 471248 283012 471260
rect 283064 471248 283070 471300
rect 284202 471248 284208 471300
rect 284260 471288 284266 471300
rect 328454 471288 328460 471300
rect 284260 471260 328460 471288
rect 284260 471248 284266 471260
rect 328454 471248 328460 471260
rect 328512 471248 328518 471300
rect 251818 470568 251824 470620
rect 251876 470608 251882 470620
rect 580166 470608 580172 470620
rect 251876 470580 580172 470608
rect 251876 470568 251882 470580
rect 580166 470568 580172 470580
rect 580224 470568 580230 470620
rect 274450 469956 274456 470008
rect 274508 469996 274514 470008
rect 342346 469996 342352 470008
rect 274508 469968 342352 469996
rect 274508 469956 274514 469968
rect 342346 469956 342352 469968
rect 342404 469956 342410 470008
rect 219066 469888 219072 469940
rect 219124 469928 219130 469940
rect 313274 469928 313280 469940
rect 219124 469900 313280 469928
rect 219124 469888 219130 469900
rect 313274 469888 313280 469900
rect 313332 469888 313338 469940
rect 25498 469820 25504 469872
rect 25556 469860 25562 469872
rect 274634 469860 274640 469872
rect 25556 469832 274640 469860
rect 25556 469820 25562 469832
rect 274634 469820 274640 469832
rect 274692 469820 274698 469872
rect 299382 469820 299388 469872
rect 299440 469860 299446 469872
rect 335354 469860 335360 469872
rect 299440 469832 335360 469860
rect 299440 469820 299446 469832
rect 335354 469820 335360 469832
rect 335412 469820 335418 469872
rect 218054 468596 218060 468648
rect 218112 468636 218118 468648
rect 269298 468636 269304 468648
rect 218112 468608 269304 468636
rect 218112 468596 218118 468608
rect 269298 468596 269304 468608
rect 269356 468596 269362 468648
rect 271690 468596 271696 468648
rect 271748 468636 271754 468648
rect 289078 468636 289084 468648
rect 271748 468608 289084 468636
rect 271748 468596 271754 468608
rect 289078 468596 289084 468608
rect 289136 468596 289142 468648
rect 291102 468596 291108 468648
rect 291160 468636 291166 468648
rect 332594 468636 332600 468648
rect 291160 468608 332600 468636
rect 291160 468596 291166 468608
rect 332594 468596 332600 468608
rect 332652 468596 332658 468648
rect 217686 468528 217692 468580
rect 217744 468568 217750 468580
rect 318886 468568 318892 468580
rect 217744 468540 318892 468568
rect 217744 468528 217750 468540
rect 318886 468528 318892 468540
rect 318944 468528 318950 468580
rect 263594 468460 263600 468512
rect 263652 468500 263658 468512
rect 396718 468500 396724 468512
rect 263652 468472 396724 468500
rect 263652 468460 263658 468472
rect 396718 468460 396724 468472
rect 396776 468460 396782 468512
rect 270402 467236 270408 467288
rect 270460 467276 270466 467288
rect 339586 467276 339592 467288
rect 270460 467248 339592 467276
rect 270460 467236 270466 467248
rect 339586 467236 339592 467248
rect 339644 467236 339650 467288
rect 21358 467168 21364 467220
rect 21416 467208 21422 467220
rect 280246 467208 280252 467220
rect 21416 467180 280252 467208
rect 21416 467168 21422 467180
rect 280246 467168 280252 467180
rect 280304 467168 280310 467220
rect 252554 467100 252560 467152
rect 252612 467140 252618 467152
rect 576118 467140 576124 467152
rect 252612 467112 576124 467140
rect 252612 467100 252618 467112
rect 576118 467100 576124 467112
rect 576176 467100 576182 467152
rect 266170 465876 266176 465928
rect 266228 465916 266234 465928
rect 297358 465916 297364 465928
rect 266228 465888 297364 465916
rect 266228 465876 266234 465888
rect 297358 465876 297364 465888
rect 297416 465876 297422 465928
rect 217778 465808 217784 465860
rect 217836 465848 217842 465860
rect 320358 465848 320364 465860
rect 217836 465820 320364 465848
rect 217836 465808 217842 465820
rect 320358 465808 320364 465820
rect 320416 465808 320422 465860
rect 88334 465740 88340 465792
rect 88392 465780 88398 465792
rect 273254 465780 273260 465792
rect 88392 465752 273260 465780
rect 88392 465740 88398 465752
rect 273254 465740 273260 465752
rect 273312 465740 273318 465792
rect 259454 465672 259460 465724
rect 259512 465712 259518 465724
rect 527174 465712 527180 465724
rect 259512 465684 527180 465712
rect 259512 465672 259518 465684
rect 527174 465672 527180 465684
rect 527232 465672 527238 465724
rect 267550 464448 267556 464500
rect 267608 464488 267614 464500
rect 335446 464488 335452 464500
rect 267608 464460 335452 464488
rect 267608 464448 267614 464460
rect 335446 464448 335452 464460
rect 335504 464448 335510 464500
rect 180058 464380 180064 464432
rect 180116 464420 180122 464432
rect 277394 464420 277400 464432
rect 180116 464392 277400 464420
rect 180116 464380 180122 464392
rect 277394 464380 277400 464392
rect 277452 464380 277458 464432
rect 251174 464312 251180 464364
rect 251232 464352 251238 464364
rect 574738 464352 574744 464364
rect 251232 464324 574744 464352
rect 251232 464312 251238 464324
rect 574738 464312 574744 464324
rect 574796 464312 574802 464364
rect 259270 462952 259276 463004
rect 259328 462992 259334 463004
rect 327166 462992 327172 463004
rect 259328 462964 327172 462992
rect 259328 462952 259334 462964
rect 327166 462952 327172 462964
rect 327224 462952 327230 463004
rect 3234 462340 3240 462392
rect 3292 462380 3298 462392
rect 284478 462380 284484 462392
rect 3292 462352 284484 462380
rect 3292 462340 3298 462352
rect 284478 462340 284484 462352
rect 284536 462340 284542 462392
rect 256510 461796 256516 461848
rect 256568 461836 256574 461848
rect 311986 461836 311992 461848
rect 256568 461808 311992 461836
rect 256568 461796 256574 461808
rect 311986 461796 311992 461808
rect 312044 461796 312050 461848
rect 278590 461728 278596 461780
rect 278648 461768 278654 461780
rect 347774 461768 347780 461780
rect 278648 461740 347780 461768
rect 278648 461728 278654 461740
rect 347774 461728 347780 461740
rect 347832 461728 347838 461780
rect 4798 461660 4804 461712
rect 4856 461700 4862 461712
rect 281626 461700 281632 461712
rect 4856 461672 281632 461700
rect 4856 461660 4862 461672
rect 281626 461660 281632 461672
rect 281684 461660 281690 461712
rect 258074 461592 258080 461644
rect 258132 461632 258138 461644
rect 580258 461632 580264 461644
rect 258132 461604 580264 461632
rect 258132 461592 258138 461604
rect 580258 461592 580264 461604
rect 580316 461592 580322 461644
rect 250990 460368 250996 460420
rect 251048 460408 251054 460420
rect 306374 460408 306380 460420
rect 251048 460380 306380 460408
rect 251048 460368 251054 460380
rect 306374 460368 306380 460380
rect 306432 460368 306438 460420
rect 277210 460300 277216 460352
rect 277268 460340 277274 460352
rect 346486 460340 346492 460352
rect 277268 460312 346492 460340
rect 277268 460300 277274 460312
rect 346486 460300 346492 460312
rect 346544 460300 346550 460352
rect 256694 460232 256700 460284
rect 256752 460272 256758 460284
rect 377398 460272 377404 460284
rect 256752 460244 377404 460272
rect 256752 460232 256758 460244
rect 377398 460232 377404 460244
rect 377456 460232 377462 460284
rect 32398 460164 32404 460216
rect 32456 460204 32462 460216
rect 278774 460204 278780 460216
rect 32456 460176 278780 460204
rect 32456 460164 32462 460176
rect 278774 460164 278780 460176
rect 278832 460164 278838 460216
rect 262030 459008 262036 459060
rect 262088 459048 262094 459060
rect 298738 459048 298744 459060
rect 262088 459020 298744 459048
rect 262088 459008 262094 459020
rect 298738 459008 298744 459020
rect 298796 459008 298802 459060
rect 273162 458940 273168 458992
rect 273220 458980 273226 458992
rect 341058 458980 341064 458992
rect 273220 458952 341064 458980
rect 273220 458940 273226 458952
rect 341058 458940 341064 458952
rect 341116 458940 341122 458992
rect 8938 458872 8944 458924
rect 8996 458912 9002 458924
rect 277486 458912 277492 458924
rect 8996 458884 277492 458912
rect 8996 458872 9002 458884
rect 277486 458872 277492 458884
rect 277544 458872 277550 458924
rect 253934 458804 253940 458856
rect 253992 458844 253998 458856
rect 570598 458844 570604 458856
rect 253992 458816 570604 458844
rect 253992 458804 253998 458816
rect 570598 458804 570604 458816
rect 570656 458804 570662 458856
rect 260650 457512 260656 457564
rect 260708 457552 260714 457564
rect 328546 457552 328552 457564
rect 260708 457524 328552 457552
rect 260708 457512 260714 457524
rect 328546 457512 328552 457524
rect 328604 457512 328610 457564
rect 153194 457444 153200 457496
rect 153252 457484 153258 457496
rect 271874 457484 271880 457496
rect 153252 457456 271880 457484
rect 153252 457444 153258 457456
rect 271874 457444 271880 457456
rect 271932 457444 271938 457496
rect 249794 456764 249800 456816
rect 249852 456804 249858 456816
rect 580166 456804 580172 456816
rect 249852 456776 580172 456804
rect 249852 456764 249858 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 251082 456152 251088 456204
rect 251140 456192 251146 456204
rect 317506 456192 317512 456204
rect 251140 456164 317512 456192
rect 251140 456152 251146 456164
rect 317506 456152 317512 456164
rect 317564 456152 317570 456204
rect 262214 456084 262220 456136
rect 262272 456124 262278 456136
rect 462314 456124 462320 456136
rect 262272 456096 462320 456124
rect 262272 456084 262278 456096
rect 462314 456084 462320 456096
rect 462372 456084 462378 456136
rect 10318 456016 10324 456068
rect 10376 456056 10382 456068
rect 276014 456056 276020 456068
rect 10376 456028 276020 456056
rect 10376 456016 10382 456028
rect 276014 456016 276020 456028
rect 276072 456016 276078 456068
rect 280062 456016 280068 456068
rect 280120 456056 280126 456068
rect 349246 456056 349252 456068
rect 280120 456028 349252 456056
rect 280120 456016 280126 456028
rect 349246 456016 349252 456028
rect 349304 456016 349310 456068
rect 252462 454792 252468 454844
rect 252520 454832 252526 454844
rect 320266 454832 320272 454844
rect 252520 454804 320272 454832
rect 252520 454792 252526 454804
rect 320266 454792 320272 454804
rect 320324 454792 320330 454844
rect 256786 454724 256792 454776
rect 256844 454764 256850 454776
rect 369118 454764 369124 454776
rect 256844 454736 369124 454764
rect 256844 454724 256850 454736
rect 369118 454724 369124 454736
rect 369176 454724 369182 454776
rect 40034 454656 40040 454708
rect 40092 454696 40098 454708
rect 274726 454696 274732 454708
rect 40092 454668 274732 454696
rect 40092 454656 40098 454668
rect 274726 454656 274732 454668
rect 274784 454656 274790 454708
rect 275922 454656 275928 454708
rect 275980 454696 275986 454708
rect 345106 454696 345112 454708
rect 275980 454668 345112 454696
rect 275980 454656 275986 454668
rect 345106 454656 345112 454668
rect 345164 454656 345170 454708
rect 249058 453432 249064 453484
rect 249116 453472 249122 453484
rect 305178 453472 305184 453484
rect 249116 453444 305184 453472
rect 249116 453432 249122 453444
rect 305178 453432 305184 453444
rect 305236 453432 305242 453484
rect 169754 453364 169760 453416
rect 169812 453404 169818 453416
rect 270494 453404 270500 453416
rect 169812 453376 270500 453404
rect 169812 453364 169818 453376
rect 270494 453364 270500 453376
rect 270552 453364 270558 453416
rect 271782 453364 271788 453416
rect 271840 453404 271846 453416
rect 340966 453404 340972 453416
rect 271840 453376 340972 453404
rect 271840 453364 271846 453376
rect 340966 453364 340972 453376
rect 341024 453364 341030 453416
rect 254026 453296 254032 453348
rect 254084 453336 254090 453348
rect 363598 453336 363604 453348
rect 254084 453308 363604 453336
rect 254084 453296 254090 453308
rect 363598 453296 363604 453308
rect 363656 453296 363662 453348
rect 246298 452004 246304 452056
rect 246356 452044 246362 452056
rect 309318 452044 309324 452056
rect 246356 452016 309324 452044
rect 246356 452004 246362 452016
rect 309318 452004 309324 452016
rect 309376 452004 309382 452056
rect 265066 451936 265072 451988
rect 265124 451976 265130 451988
rect 364334 451976 364340 451988
rect 265124 451948 364340 451976
rect 265124 451936 265130 451948
rect 364334 451936 364340 451948
rect 364392 451936 364398 451988
rect 7558 451868 7564 451920
rect 7616 451908 7622 451920
rect 278866 451908 278872 451920
rect 7616 451880 278872 451908
rect 7616 451868 7622 451880
rect 278866 451868 278872 451880
rect 278924 451868 278930 451920
rect 288342 451868 288348 451920
rect 288400 451908 288406 451920
rect 331214 451908 331220 451920
rect 288400 451880 331220 451908
rect 288400 451868 288406 451880
rect 331214 451868 331220 451880
rect 331272 451868 331278 451920
rect 253750 450712 253756 450764
rect 253808 450752 253814 450764
rect 321646 450752 321652 450764
rect 253808 450724 321652 450752
rect 253808 450712 253814 450724
rect 321646 450712 321652 450724
rect 321704 450712 321710 450764
rect 217318 450644 217324 450696
rect 217376 450684 217382 450696
rect 302326 450684 302332 450696
rect 217376 450656 302332 450684
rect 217376 450644 217382 450656
rect 302326 450644 302332 450656
rect 302384 450644 302390 450696
rect 263686 450576 263692 450628
rect 263744 450616 263750 450628
rect 428458 450616 428464 450628
rect 263744 450588 428464 450616
rect 263744 450576 263750 450588
rect 428458 450576 428464 450588
rect 428516 450576 428522 450628
rect 13078 450508 13084 450560
rect 13136 450548 13142 450560
rect 274818 450548 274824 450560
rect 13136 450520 274824 450548
rect 13136 450508 13142 450520
rect 274818 450508 274824 450520
rect 274876 450508 274882 450560
rect 293862 449284 293868 449336
rect 293920 449324 293926 449336
rect 333974 449324 333980 449336
rect 293920 449296 333980 449324
rect 293920 449284 293926 449296
rect 333974 449284 333980 449296
rect 334032 449284 334038 449336
rect 247678 449216 247684 449268
rect 247736 449256 247742 449268
rect 310606 449256 310612 449268
rect 247736 449228 310612 449256
rect 247736 449216 247742 449228
rect 310606 449216 310612 449228
rect 310664 449216 310670 449268
rect 258166 449148 258172 449200
rect 258224 449188 258230 449200
rect 371878 449188 371884 449200
rect 258224 449160 371884 449188
rect 258224 449148 258230 449160
rect 371878 449148 371884 449160
rect 371936 449148 371942 449200
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 284386 448576 284392 448588
rect 3200 448548 284392 448576
rect 3200 448536 3206 448548
rect 284386 448536 284392 448548
rect 284444 448536 284450 448588
rect 256602 447924 256608 447976
rect 256660 447964 256666 447976
rect 324406 447964 324412 447976
rect 256660 447936 324412 447964
rect 256660 447924 256666 447936
rect 324406 447924 324412 447936
rect 324464 447924 324470 447976
rect 71774 447856 71780 447908
rect 71832 447896 71838 447908
rect 273346 447896 273352 447908
rect 71832 447868 273352 447896
rect 71832 447856 71838 447868
rect 273346 447856 273352 447868
rect 273404 447856 273410 447908
rect 296622 447856 296628 447908
rect 296680 447896 296686 447908
rect 335538 447896 335544 447908
rect 296680 447868 335544 447896
rect 296680 447856 296686 447868
rect 335538 447856 335544 447868
rect 335596 447856 335602 447908
rect 260834 447788 260840 447840
rect 260892 447828 260898 447840
rect 494054 447828 494060 447840
rect 260892 447800 494060 447828
rect 260892 447788 260898 447800
rect 494054 447788 494060 447800
rect 494112 447788 494118 447840
rect 260742 446496 260748 446548
rect 260800 446536 260806 446548
rect 330018 446536 330024 446548
rect 260800 446508 330024 446536
rect 260800 446496 260806 446508
rect 330018 446496 330024 446508
rect 330076 446496 330082 446548
rect 259546 446428 259552 446480
rect 259604 446468 259610 446480
rect 367738 446468 367744 446480
rect 259604 446440 367744 446468
rect 259604 446428 259610 446440
rect 367738 446428 367744 446440
rect 367796 446428 367802 446480
rect 138658 446360 138664 446412
rect 138716 446400 138722 446412
rect 270586 446400 270592 446412
rect 138716 446372 270592 446400
rect 138716 446360 138722 446372
rect 270586 446360 270592 446372
rect 270644 446360 270650 446412
rect 206278 445136 206284 445188
rect 206336 445176 206342 445188
rect 271966 445176 271972 445188
rect 206336 445148 271972 445176
rect 206336 445136 206342 445148
rect 271966 445136 271972 445148
rect 272024 445136 272030 445188
rect 257982 445068 257988 445120
rect 258040 445108 258046 445120
rect 325694 445108 325700 445120
rect 258040 445080 325700 445108
rect 258040 445068 258046 445080
rect 325694 445068 325700 445080
rect 325752 445068 325758 445120
rect 258258 445000 258264 445052
rect 258316 445040 258322 445052
rect 360838 445040 360844 445052
rect 258316 445012 360844 445040
rect 258316 445000 258322 445012
rect 360838 445000 360844 445012
rect 360896 445000 360902 445052
rect 201494 443776 201500 443828
rect 201552 443816 201558 443828
rect 269206 443816 269212 443828
rect 201552 443788 269212 443816
rect 201552 443776 201558 443788
rect 269206 443776 269212 443788
rect 269264 443776 269270 443828
rect 278682 443776 278688 443828
rect 278740 443816 278746 443828
rect 325786 443816 325792 443828
rect 278740 443788 325792 443816
rect 278740 443776 278746 443788
rect 325786 443776 325792 443788
rect 325844 443776 325850 443828
rect 219158 443708 219164 443760
rect 219216 443748 219222 443760
rect 314746 443748 314752 443760
rect 219216 443720 314752 443748
rect 219216 443708 219222 443720
rect 314746 443708 314752 443720
rect 314804 443708 314810 443760
rect 255406 443640 255412 443692
rect 255464 443680 255470 443692
rect 432598 443680 432604 443692
rect 255464 443652 432604 443680
rect 255464 443640 255470 443652
rect 432598 443640 432604 443652
rect 432656 443640 432662 443692
rect 277302 442416 277308 442468
rect 277360 442456 277366 442468
rect 325878 442456 325884 442468
rect 277360 442428 325884 442456
rect 277360 442416 277366 442428
rect 325878 442416 325884 442428
rect 325936 442416 325942 442468
rect 249702 442348 249708 442400
rect 249760 442388 249766 442400
rect 314838 442388 314844 442400
rect 249760 442360 314844 442388
rect 249760 442348 249766 442360
rect 314838 442348 314844 442360
rect 314896 442348 314902 442400
rect 182818 442280 182824 442332
rect 182876 442320 182882 442332
rect 278958 442320 278964 442332
rect 182876 442292 278964 442320
rect 182876 442280 182882 442292
rect 278958 442280 278964 442292
rect 279016 442280 279022 442332
rect 254118 442212 254124 442264
rect 254176 442252 254182 442264
rect 359458 442252 359464 442264
rect 254176 442224 359464 442252
rect 254176 442212 254182 442224
rect 359458 442212 359464 442224
rect 359516 442212 359522 442264
rect 248230 440988 248236 441040
rect 248288 441028 248294 441040
rect 314102 441028 314108 441040
rect 248288 441000 314108 441028
rect 248288 440988 248294 441000
rect 314102 440988 314108 441000
rect 314160 440988 314166 441040
rect 14458 440920 14464 440972
rect 14516 440960 14522 440972
rect 277026 440960 277032 440972
rect 14516 440932 277032 440960
rect 14516 440920 14522 440932
rect 277026 440920 277032 440932
rect 277084 440920 277090 440972
rect 286962 440920 286968 440972
rect 287020 440960 287026 440972
rect 330570 440960 330576 440972
rect 287020 440932 330576 440960
rect 287020 440920 287026 440932
rect 330570 440920 330576 440932
rect 330628 440920 330634 440972
rect 252738 440852 252744 440904
rect 252796 440892 252802 440904
rect 578878 440892 578884 440904
rect 252796 440864 578884 440892
rect 252796 440852 252802 440864
rect 578878 440852 578884 440864
rect 578936 440852 578942 440904
rect 245470 439832 245476 439884
rect 245528 439872 245534 439884
rect 306834 439872 306840 439884
rect 245528 439844 306840 439872
rect 245528 439832 245534 439844
rect 306834 439832 306840 439844
rect 306892 439832 306898 439884
rect 266262 439764 266268 439816
rect 266320 439804 266326 439816
rect 334802 439804 334808 439816
rect 266320 439776 334808 439804
rect 266320 439764 266326 439776
rect 334802 439764 334808 439776
rect 334860 439764 334866 439816
rect 264790 439696 264796 439748
rect 264848 439736 264854 439748
rect 333606 439736 333612 439748
rect 264848 439708 333612 439736
rect 264848 439696 264854 439708
rect 333606 439696 333612 439708
rect 333664 439696 333670 439748
rect 263502 439628 263508 439680
rect 263560 439668 263566 439680
rect 332318 439668 332324 439680
rect 263560 439640 332324 439668
rect 263560 439628 263566 439640
rect 332318 439628 332324 439640
rect 332376 439628 332382 439680
rect 268930 439560 268936 439612
rect 268988 439600 268994 439612
rect 338390 439600 338396 439612
rect 268988 439572 338396 439600
rect 268988 439560 268994 439572
rect 338390 439560 338396 439572
rect 338448 439560 338454 439612
rect 267642 439492 267648 439544
rect 267700 439532 267706 439544
rect 337194 439532 337200 439544
rect 267700 439504 337200 439532
rect 267700 439492 267706 439504
rect 337194 439492 337200 439504
rect 337252 439492 337258 439544
rect 338758 439492 338764 439544
rect 338816 439532 338822 439544
rect 348786 439532 348792 439544
rect 338816 439504 348792 439532
rect 338816 439492 338822 439504
rect 348786 439492 348792 439504
rect 348844 439492 348850 439544
rect 244182 438268 244188 438320
rect 244240 438308 244246 438320
rect 304350 438308 304356 438320
rect 244240 438280 304356 438308
rect 244240 438268 244246 438280
rect 304350 438268 304356 438280
rect 304408 438268 304414 438320
rect 262122 438200 262128 438252
rect 262180 438240 262186 438252
rect 331122 438240 331128 438252
rect 262180 438212 331128 438240
rect 262180 438200 262186 438212
rect 331122 438200 331128 438212
rect 331180 438200 331186 438252
rect 274358 438132 274364 438184
rect 274416 438172 274422 438184
rect 344554 438172 344560 438184
rect 274416 438144 344560 438172
rect 274416 438132 274422 438144
rect 344554 438132 344560 438144
rect 344612 438132 344618 438184
rect 264882 437044 264888 437096
rect 264940 437084 264946 437096
rect 264940 437056 268608 437084
rect 264940 437044 264946 437056
rect 219342 436908 219348 436960
rect 219400 436948 219406 436960
rect 267918 436948 267924 436960
rect 219400 436920 267924 436948
rect 219400 436908 219406 436920
rect 267918 436908 267924 436920
rect 267976 436908 267982 436960
rect 258166 436840 258172 436892
rect 258224 436880 258230 436892
rect 258534 436880 258540 436892
rect 258224 436852 258540 436880
rect 258224 436840 258230 436852
rect 258534 436840 258540 436852
rect 258592 436840 258598 436892
rect 268580 436880 268608 437056
rect 273254 436908 273260 436960
rect 273312 436948 273318 436960
rect 273622 436948 273628 436960
rect 273312 436920 273628 436948
rect 273312 436908 273318 436920
rect 273622 436908 273628 436920
rect 273680 436908 273686 436960
rect 274634 436908 274640 436960
rect 274692 436948 274698 436960
rect 275462 436948 275468 436960
rect 274692 436920 275468 436948
rect 274692 436908 274698 436920
rect 275462 436908 275468 436920
rect 275520 436908 275526 436960
rect 278774 436908 278780 436960
rect 278832 436948 278838 436960
rect 279694 436948 279700 436960
rect 278832 436920 279700 436948
rect 278832 436908 278838 436920
rect 279694 436908 279700 436920
rect 279752 436908 279758 436960
rect 281534 436908 281540 436960
rect 281592 436948 281598 436960
rect 282086 436948 282092 436960
rect 281592 436920 282092 436948
rect 281592 436908 281598 436920
rect 282086 436908 282092 436920
rect 282144 436908 282150 436960
rect 282914 436908 282920 436960
rect 282972 436948 282978 436960
rect 283374 436948 283380 436960
rect 282972 436920 283380 436948
rect 282972 436908 282978 436920
rect 283374 436908 283380 436920
rect 283432 436908 283438 436960
rect 311894 436908 311900 436960
rect 311952 436948 311958 436960
rect 312630 436948 312636 436960
rect 311952 436920 312636 436948
rect 311952 436908 311958 436920
rect 312630 436908 312636 436920
rect 312688 436908 312694 436960
rect 317414 436908 317420 436960
rect 317472 436948 317478 436960
rect 317966 436948 317972 436960
rect 317472 436920 317972 436948
rect 317472 436908 317478 436920
rect 317966 436908 317972 436920
rect 318024 436908 318030 436960
rect 318794 436908 318800 436960
rect 318852 436948 318858 436960
rect 319254 436948 319260 436960
rect 318852 436920 319260 436948
rect 318852 436908 318858 436920
rect 319254 436908 319260 436920
rect 319312 436908 319318 436960
rect 320266 436908 320272 436960
rect 320324 436948 320330 436960
rect 321094 436948 321100 436960
rect 320324 436920 321100 436948
rect 320324 436908 320330 436920
rect 321094 436908 321100 436920
rect 321152 436908 321158 436960
rect 325786 436908 325792 436960
rect 325844 436948 325850 436960
rect 326614 436948 326620 436960
rect 325844 436920 326620 436948
rect 325844 436908 325850 436920
rect 326614 436908 326620 436920
rect 326672 436908 326678 436960
rect 327074 436908 327080 436960
rect 327132 436948 327138 436960
rect 327718 436948 327724 436960
rect 327132 436920 327724 436948
rect 327132 436908 327138 436920
rect 327718 436908 327724 436920
rect 327776 436908 327782 436960
rect 328454 436908 328460 436960
rect 328512 436948 328518 436960
rect 329006 436948 329012 436960
rect 328512 436920 329012 436948
rect 328512 436908 328518 436920
rect 329006 436908 329012 436920
rect 329064 436908 329070 436960
rect 345106 436908 345112 436960
rect 345164 436948 345170 436960
rect 345382 436948 345388 436960
rect 345164 436920 345388 436948
rect 345164 436908 345170 436920
rect 345382 436908 345388 436920
rect 345440 436908 345446 436960
rect 412634 436880 412640 436892
rect 268580 436852 412640 436880
rect 412634 436840 412640 436852
rect 412692 436840 412698 436892
rect 254026 436772 254032 436824
rect 254084 436812 254090 436824
rect 254854 436812 254860 436824
rect 254084 436784 254860 436812
rect 254084 436772 254090 436784
rect 254854 436772 254860 436784
rect 254912 436772 254918 436824
rect 256694 436772 256700 436824
rect 256752 436812 256758 436824
rect 257246 436812 257252 436824
rect 256752 436784 257252 436812
rect 256752 436772 256758 436784
rect 257246 436772 257252 436784
rect 257304 436772 257310 436824
rect 258074 436772 258080 436824
rect 258132 436812 258138 436824
rect 259086 436812 259092 436824
rect 258132 436784 259092 436812
rect 258132 436772 258138 436784
rect 259086 436772 259092 436784
rect 259144 436772 259150 436824
rect 259454 436772 259460 436824
rect 259512 436812 259518 436824
rect 260374 436812 260380 436824
rect 259512 436784 260380 436812
rect 259512 436772 259518 436784
rect 260374 436772 260380 436784
rect 260432 436772 260438 436824
rect 268562 436772 268568 436824
rect 268620 436812 268626 436824
rect 477494 436812 477500 436824
rect 268620 436784 477500 436812
rect 268620 436772 268626 436784
rect 477494 436772 477500 436784
rect 477552 436772 477558 436824
rect 263778 436704 263784 436756
rect 263836 436744 263842 436756
rect 542354 436744 542360 436756
rect 263836 436716 542360 436744
rect 263836 436704 263842 436716
rect 542354 436704 542360 436716
rect 542412 436704 542418 436756
rect 231210 436636 231216 436688
rect 231268 436676 231274 436688
rect 286134 436676 286140 436688
rect 231268 436648 286140 436676
rect 231268 436636 231274 436648
rect 286134 436636 286140 436648
rect 286192 436636 286198 436688
rect 325694 436636 325700 436688
rect 325752 436676 325758 436688
rect 325970 436676 325976 436688
rect 325752 436648 325976 436676
rect 325752 436636 325758 436648
rect 325970 436636 325976 436648
rect 326028 436636 326034 436688
rect 210418 436568 210424 436620
rect 210476 436608 210482 436620
rect 295886 436608 295892 436620
rect 210476 436580 295892 436608
rect 210476 436568 210482 436580
rect 295886 436568 295892 436580
rect 295944 436568 295950 436620
rect 203518 436500 203524 436552
rect 203576 436540 203582 436552
rect 295242 436540 295248 436552
rect 203576 436512 295248 436540
rect 203576 436500 203582 436512
rect 295242 436500 295248 436512
rect 295300 436500 295306 436552
rect 197998 436432 198004 436484
rect 198056 436472 198062 436484
rect 297726 436472 297732 436484
rect 198056 436444 297732 436472
rect 198056 436432 198062 436444
rect 297726 436432 297732 436444
rect 297784 436432 297790 436484
rect 244826 436364 244832 436416
rect 244884 436404 244890 436416
rect 353938 436404 353944 436416
rect 244884 436376 353944 436404
rect 244884 436364 244890 436376
rect 353938 436364 353944 436376
rect 353996 436364 354002 436416
rect 244182 436296 244188 436348
rect 244240 436336 244246 436348
rect 355318 436336 355324 436348
rect 244240 436308 355324 436336
rect 244240 436296 244246 436308
rect 355318 436296 355324 436308
rect 355376 436296 355382 436348
rect 88978 436228 88984 436280
rect 89036 436268 89042 436280
rect 300762 436268 300768 436280
rect 89036 436240 300768 436268
rect 89036 436228 89042 436240
rect 300762 436228 300768 436240
rect 300820 436228 300826 436280
rect 14550 436160 14556 436212
rect 14608 436200 14614 436212
rect 291654 436200 291660 436212
rect 14608 436172 291660 436200
rect 14608 436160 14614 436172
rect 291654 436160 291660 436172
rect 291712 436160 291718 436212
rect 8938 436092 8944 436144
rect 8996 436132 9002 436144
rect 292206 436132 292212 436144
rect 8996 436104 292212 436132
rect 8996 436092 9002 436104
rect 292206 436092 292212 436104
rect 292264 436092 292270 436144
rect 263042 435752 263048 435804
rect 263100 435792 263106 435804
rect 268562 435792 268568 435804
rect 263100 435764 268568 435792
rect 263100 435752 263106 435764
rect 268562 435752 268568 435764
rect 268620 435752 268626 435804
rect 261202 435684 261208 435736
rect 261260 435724 261266 435736
rect 263778 435724 263784 435736
rect 261260 435696 263784 435724
rect 261260 435684 261266 435696
rect 263778 435684 263784 435696
rect 263836 435684 263842 435736
rect 98638 435208 98644 435260
rect 98696 435248 98702 435260
rect 289170 435248 289176 435260
rect 98696 435220 289176 435248
rect 98696 435208 98702 435220
rect 289170 435208 289176 435220
rect 289228 435208 289234 435260
rect 225598 435140 225604 435192
rect 225656 435180 225662 435192
rect 291010 435180 291016 435192
rect 225656 435152 291016 435180
rect 225656 435140 225662 435152
rect 291010 435140 291016 435152
rect 291068 435140 291074 435192
rect 207658 435072 207664 435124
rect 207716 435112 207722 435124
rect 298278 435112 298284 435124
rect 207716 435084 298284 435112
rect 207716 435072 207722 435084
rect 298278 435072 298284 435084
rect 298336 435072 298342 435124
rect 246022 435004 246028 435056
rect 246080 435044 246086 435056
rect 356698 435044 356704 435056
rect 246080 435016 356704 435044
rect 246080 435004 246086 435016
rect 356698 435004 356704 435016
rect 356756 435004 356762 435056
rect 100018 434936 100024 434988
rect 100076 434976 100082 434988
rect 287330 434976 287336 434988
rect 100076 434948 287336 434976
rect 100076 434936 100082 434948
rect 287330 434936 287336 434948
rect 287388 434936 287394 434988
rect 7558 434868 7564 434920
rect 7616 434908 7622 434920
rect 285490 434908 285496 434920
rect 7616 434880 285496 434908
rect 7616 434868 7622 434880
rect 285490 434868 285496 434880
rect 285548 434868 285554 434920
rect 285674 434868 285680 434920
rect 285732 434908 285738 434920
rect 580902 434908 580908 434920
rect 285732 434880 580908 434908
rect 285732 434868 285738 434880
rect 580902 434868 580908 434880
rect 580960 434868 580966 434920
rect 282178 434800 282184 434852
rect 282236 434840 282242 434852
rect 580534 434840 580540 434852
rect 282236 434812 580540 434840
rect 282236 434800 282242 434812
rect 580534 434800 580540 434812
rect 580592 434800 580598 434852
rect 241146 434732 241152 434784
rect 241204 434772 241210 434784
rect 577498 434772 577504 434784
rect 241204 434744 577504 434772
rect 241204 434732 241210 434744
rect 577498 434732 577504 434744
rect 577556 434732 577562 434784
rect 309134 434596 309140 434648
rect 309192 434636 309198 434648
rect 310054 434636 310060 434648
rect 309192 434608 310060 434636
rect 309192 434596 309198 434608
rect 310054 434596 310060 434608
rect 310112 434596 310118 434648
rect 335630 434596 335636 434648
rect 335688 434636 335694 434648
rect 335998 434636 336004 434648
rect 335688 434608 336004 434636
rect 335688 434596 335694 434608
rect 335998 434596 336004 434608
rect 336056 434596 336062 434648
rect 263594 434528 263600 434580
rect 263652 434568 263658 434580
rect 263870 434568 263876 434580
rect 263652 434540 263876 434568
rect 263652 434528 263658 434540
rect 263870 434528 263876 434540
rect 263928 434528 263934 434580
rect 264974 434528 264980 434580
rect 265032 434568 265038 434580
rect 265710 434568 265716 434580
rect 265032 434540 265716 434568
rect 265032 434528 265038 434540
rect 265710 434528 265716 434540
rect 265768 434528 265774 434580
rect 302234 434528 302240 434580
rect 302292 434568 302298 434580
rect 302878 434568 302884 434580
rect 302292 434540 302884 434568
rect 302292 434528 302298 434540
rect 302878 434528 302884 434540
rect 302936 434528 302942 434580
rect 305086 434528 305092 434580
rect 305144 434568 305150 434580
rect 305822 434568 305828 434580
rect 305144 434540 305828 434568
rect 305144 434528 305150 434540
rect 305822 434528 305828 434540
rect 305880 434528 305886 434580
rect 309226 434528 309232 434580
rect 309284 434568 309290 434580
rect 309502 434568 309508 434580
rect 309284 434540 309508 434568
rect 309284 434528 309290 434540
rect 309502 434528 309508 434540
rect 309560 434528 309566 434580
rect 335354 434528 335360 434580
rect 335412 434568 335418 434580
rect 336366 434568 336372 434580
rect 335412 434540 336372 434568
rect 335412 434528 335418 434540
rect 336366 434528 336372 434540
rect 336424 434528 336430 434580
rect 243538 434460 243544 434512
rect 243596 434500 243602 434512
rect 352558 434500 352564 434512
rect 243596 434472 352564 434500
rect 243596 434460 243602 434472
rect 352558 434460 352564 434472
rect 352616 434460 352622 434512
rect 327810 434392 327816 434444
rect 327868 434432 327874 434444
rect 346302 434432 346308 434444
rect 327868 434404 346308 434432
rect 327868 434392 327874 434404
rect 346302 434392 346308 434404
rect 346360 434392 346366 434444
rect 329098 434324 329104 434376
rect 329156 434364 329162 434376
rect 347590 434364 347596 434376
rect 329156 434336 347596 434364
rect 329156 434324 329162 434336
rect 347590 434324 347596 434336
rect 347648 434324 347654 434376
rect 331858 434256 331864 434308
rect 331916 434296 331922 434308
rect 349982 434296 349988 434308
rect 331916 434268 349988 434296
rect 331916 434256 331922 434268
rect 349982 434256 349988 434268
rect 350040 434256 350046 434308
rect 94498 434188 94504 434240
rect 94556 434228 94562 434240
rect 290366 434228 290372 434240
rect 94556 434200 290372 434228
rect 94556 434188 94562 434200
rect 290366 434188 290372 434200
rect 290424 434188 290430 434240
rect 324958 434188 324964 434240
rect 325016 434228 325022 434240
rect 342714 434228 342720 434240
rect 325016 434200 342720 434228
rect 325016 434188 325022 434200
rect 342714 434188 342720 434200
rect 342772 434188 342778 434240
rect 246666 434120 246672 434172
rect 246724 434160 246730 434172
rect 285674 434160 285680 434172
rect 246724 434132 285680 434160
rect 246724 434120 246730 434132
rect 285674 434120 285680 434132
rect 285732 434120 285738 434172
rect 298738 434120 298744 434172
rect 298796 434160 298802 434172
rect 316586 434160 316592 434172
rect 298796 434132 316592 434160
rect 298796 434120 298802 434132
rect 316586 434120 316592 434132
rect 316644 434120 316650 434172
rect 322382 434120 322388 434172
rect 322440 434160 322446 434172
rect 340230 434160 340236 434172
rect 322440 434132 340236 434160
rect 322440 434120 322446 434132
rect 340230 434120 340236 434132
rect 340288 434120 340294 434172
rect 238754 434052 238760 434104
rect 238812 434092 238818 434104
rect 282178 434092 282184 434104
rect 238812 434064 282184 434092
rect 238812 434052 238818 434064
rect 282178 434052 282184 434064
rect 282236 434052 282242 434104
rect 297358 434052 297364 434104
rect 297416 434092 297422 434104
rect 320174 434092 320180 434104
rect 297416 434064 320180 434092
rect 297416 434052 297422 434064
rect 320174 434052 320180 434064
rect 320232 434052 320238 434104
rect 320818 434052 320824 434104
rect 320876 434092 320882 434104
rect 339034 434092 339040 434104
rect 320876 434064 339040 434092
rect 320876 434052 320882 434064
rect 339034 434052 339040 434064
rect 339092 434052 339098 434104
rect 217870 433984 217876 434036
rect 217928 434024 217934 434036
rect 269114 434024 269120 434036
rect 217928 433996 269120 434024
rect 217928 433984 217934 433996
rect 269114 433984 269120 433996
rect 269172 433984 269178 434036
rect 279970 434024 279976 434036
rect 269224 433996 279976 434024
rect 240502 433848 240508 433900
rect 240560 433888 240566 433900
rect 269224 433888 269252 433996
rect 279970 433984 279976 433996
rect 280028 433984 280034 434036
rect 289078 433984 289084 434036
rect 289136 434024 289142 434036
rect 323210 434024 323216 434036
rect 289136 433996 323216 434024
rect 289136 433984 289142 433996
rect 323210 433984 323216 433996
rect 323268 433984 323274 434036
rect 323578 433984 323584 434036
rect 323636 434024 323642 434036
rect 341518 434024 341524 434036
rect 323636 433996 341524 434024
rect 323636 433984 323642 433996
rect 341518 433984 341524 433996
rect 341576 433984 341582 434036
rect 269390 433916 269396 433968
rect 269448 433956 269454 433968
rect 287974 433956 287980 433968
rect 269448 433928 287980 433956
rect 269448 433916 269454 433928
rect 287974 433916 287980 433928
rect 288032 433916 288038 433968
rect 240560 433860 269252 433888
rect 240560 433848 240566 433860
rect 248414 433780 248420 433832
rect 248472 433820 248478 433832
rect 289722 433820 289728 433832
rect 248472 433792 289728 433820
rect 248472 433780 248478 433792
rect 289722 433780 289728 433792
rect 289780 433780 289786 433832
rect 242342 433712 242348 433764
rect 242400 433752 242406 433764
rect 282914 433752 282920 433764
rect 242400 433724 282920 433752
rect 242400 433712 242406 433724
rect 282914 433712 282920 433724
rect 282972 433712 282978 433764
rect 229738 433644 229744 433696
rect 229796 433684 229802 433696
rect 286778 433684 286784 433696
rect 229796 433656 286784 433684
rect 229796 433644 229802 433656
rect 286778 433644 286784 433656
rect 286836 433644 286842 433696
rect 231118 433576 231124 433628
rect 231176 433616 231182 433628
rect 288618 433616 288624 433628
rect 231176 433588 288624 433616
rect 231176 433576 231182 433588
rect 288618 433576 288624 433588
rect 288676 433576 288682 433628
rect 209038 433508 209044 433560
rect 209096 433548 209102 433560
rect 292850 433548 292856 433560
rect 209096 433520 292856 433548
rect 209096 433508 209102 433520
rect 292850 433508 292856 433520
rect 292908 433508 292914 433560
rect 199378 433440 199384 433492
rect 199436 433480 199442 433492
rect 294046 433480 294052 433492
rect 199436 433452 294052 433480
rect 199436 433440 199442 433452
rect 294046 433440 294052 433452
rect 294104 433440 294110 433492
rect 350626 433440 350632 433492
rect 350684 433480 350690 433492
rect 480898 433480 480904 433492
rect 350684 433452 480904 433480
rect 350684 433440 350690 433452
rect 480898 433440 480904 433452
rect 480956 433440 480962 433492
rect 247862 433372 247868 433424
rect 247920 433412 247926 433424
rect 262674 433412 262680 433424
rect 247920 433384 262680 433412
rect 247920 433372 247926 433384
rect 262674 433372 262680 433384
rect 262732 433372 262738 433424
rect 351178 433372 351184 433424
rect 351236 433412 351242 433424
rect 581086 433412 581092 433424
rect 351236 433384 581092 433412
rect 351236 433372 351242 433384
rect 581086 433372 581092 433384
rect 581144 433372 581150 433424
rect 249702 433304 249708 433356
rect 249760 433344 249766 433356
rect 272242 433344 272248 433356
rect 249760 433316 272248 433344
rect 249760 433304 249766 433316
rect 272242 433304 272248 433316
rect 272300 433304 272306 433356
rect 280062 433304 280068 433356
rect 280120 433344 280126 433356
rect 289814 433344 289820 433356
rect 280120 433316 289820 433344
rect 280120 433304 280126 433316
rect 289814 433304 289820 433316
rect 289872 433304 289878 433356
rect 304902 433304 304908 433356
rect 304960 433344 304966 433356
rect 305178 433344 305184 433356
rect 304960 433316 305184 433344
rect 304960 433304 304966 433316
rect 305178 433304 305184 433316
rect 305236 433304 305242 433356
rect 351822 433304 351828 433356
rect 351880 433344 351886 433356
rect 582374 433344 582380 433356
rect 351880 433316 582380 433344
rect 351880 433304 351886 433316
rect 582374 433304 582380 433316
rect 582432 433304 582438 433356
rect 289722 432760 289728 432812
rect 289780 432800 289786 432812
rect 580166 432800 580172 432812
rect 289780 432772 580172 432800
rect 289780 432760 289786 432772
rect 580166 432760 580172 432772
rect 580224 432760 580230 432812
rect 3602 432692 3608 432744
rect 3660 432732 3666 432744
rect 269390 432732 269396 432744
rect 3660 432704 269396 432732
rect 3660 432692 3666 432704
rect 269390 432692 269396 432704
rect 269448 432692 269454 432744
rect 279970 432692 279976 432744
rect 280028 432732 280034 432744
rect 280028 432704 280200 432732
rect 280028 432692 280034 432704
rect 3510 432624 3516 432676
rect 3568 432664 3574 432676
rect 280062 432664 280068 432676
rect 3568 432636 280068 432664
rect 3568 432624 3574 432636
rect 280062 432624 280068 432636
rect 280120 432624 280126 432676
rect 280172 432664 280200 432704
rect 282914 432692 282920 432744
rect 282972 432732 282978 432744
rect 580626 432732 580632 432744
rect 282972 432704 580632 432732
rect 282972 432692 282978 432704
rect 580626 432692 580632 432704
rect 580684 432692 580690 432744
rect 580718 432664 580724 432676
rect 280172 432636 580724 432664
rect 580718 432624 580724 432636
rect 580776 432624 580782 432676
rect 3418 432556 3424 432608
rect 3476 432596 3482 432608
rect 253198 432596 253204 432608
rect 3476 432568 253204 432596
rect 3476 432556 3482 432568
rect 253198 432556 253204 432568
rect 253256 432556 253262 432608
rect 262674 432556 262680 432608
rect 262732 432596 262738 432608
rect 580074 432596 580080 432608
rect 262732 432568 580080 432596
rect 262732 432556 262738 432568
rect 580074 432556 580080 432568
rect 580132 432556 580138 432608
rect 97902 432488 97908 432540
rect 97960 432528 97966 432540
rect 251818 432528 251824 432540
rect 97960 432500 251824 432528
rect 97960 432488 97966 432500
rect 251818 432488 251824 432500
rect 251876 432488 251882 432540
rect 206278 432420 206284 432472
rect 206336 432460 206342 432472
rect 293402 432460 293408 432472
rect 206336 432432 293408 432460
rect 206336 432420 206342 432432
rect 293402 432420 293408 432432
rect 293460 432420 293466 432472
rect 200758 432352 200764 432404
rect 200816 432392 200822 432404
rect 297082 432392 297088 432404
rect 200816 432364 297088 432392
rect 200816 432352 200822 432364
rect 297082 432352 297088 432364
rect 297140 432352 297146 432404
rect 196618 432284 196624 432336
rect 196676 432324 196682 432336
rect 301038 432324 301044 432336
rect 196676 432296 301044 432324
rect 196676 432284 196682 432296
rect 301038 432284 301044 432296
rect 301096 432284 301102 432336
rect 140774 432216 140780 432268
rect 140832 432256 140838 432268
rect 249426 432256 249432 432268
rect 140832 432228 249432 432256
rect 140832 432216 140838 432228
rect 249426 432216 249432 432228
rect 249484 432256 249490 432268
rect 352834 432256 352840 432268
rect 249484 432228 352840 432256
rect 249484 432216 249490 432228
rect 352834 432216 352840 432228
rect 352892 432216 352898 432268
rect 247586 432148 247592 432200
rect 247644 432188 247650 432200
rect 352742 432188 352748 432200
rect 247644 432160 352748 432188
rect 247644 432148 247650 432160
rect 352742 432148 352748 432160
rect 352800 432148 352806 432200
rect 242066 432080 242072 432132
rect 242124 432120 242130 432132
rect 358078 432120 358084 432132
rect 242124 432092 358084 432120
rect 242124 432080 242130 432092
rect 358078 432080 358084 432092
rect 358136 432080 358142 432132
rect 245562 432012 245568 432064
rect 245620 432052 245626 432064
rect 352650 432052 352656 432064
rect 245620 432024 352656 432052
rect 245620 432012 245626 432024
rect 352650 432012 352656 432024
rect 352708 432012 352714 432064
rect 233602 431944 233608 431996
rect 233660 431984 233666 431996
rect 580350 431984 580356 431996
rect 233660 431956 580356 431984
rect 233660 431944 233666 431956
rect 580350 431944 580356 431956
rect 580408 431944 580414 431996
rect 272242 431876 272248 431928
rect 272300 431916 272306 431928
rect 579890 431916 579896 431928
rect 272300 431888 579896 431916
rect 272300 431876 272306 431888
rect 579890 431876 579896 431888
rect 579948 431876 579954 431928
rect 250530 431740 250536 431792
rect 250588 431780 250594 431792
rect 250588 431752 258074 431780
rect 250588 431740 250594 431752
rect 258046 430624 258074 431752
rect 355410 430624 355416 430636
rect 258046 430596 355416 430624
rect 355410 430584 355416 430596
rect 355468 430584 355474 430636
rect 580718 427320 580724 427372
rect 580776 427320 580782 427372
rect 580736 427168 580764 427320
rect 579982 427116 579988 427168
rect 580040 427156 580046 427168
rect 580626 427156 580632 427168
rect 580040 427128 580632 427156
rect 580040 427116 580046 427128
rect 580626 427116 580632 427128
rect 580684 427116 580690 427168
rect 580718 427116 580724 427168
rect 580776 427116 580782 427168
rect 3326 423580 3332 423632
rect 3384 423620 3390 423632
rect 7558 423620 7564 423632
rect 3384 423592 7564 423620
rect 3384 423580 3390 423592
rect 7558 423580 7564 423592
rect 7616 423580 7622 423632
rect 355410 419432 355416 419484
rect 355468 419472 355474 419484
rect 579982 419472 579988 419484
rect 355468 419444 579988 419472
rect 355468 419432 355474 419444
rect 579982 419432 579988 419444
rect 580040 419432 580046 419484
rect 3326 411204 3332 411256
rect 3384 411244 3390 411256
rect 229738 411244 229744 411256
rect 3384 411216 229744 411244
rect 3384 411204 3390 411216
rect 229738 411204 229744 411216
rect 229796 411204 229802 411256
rect 352834 405628 352840 405680
rect 352892 405668 352898 405680
rect 579982 405668 579988 405680
rect 352892 405640 579988 405668
rect 352892 405628 352898 405640
rect 579982 405628 579988 405640
rect 580040 405628 580046 405680
rect 3326 398760 3332 398812
rect 3384 398800 3390 398812
rect 231210 398800 231216 398812
rect 3384 398772 231216 398800
rect 3384 398760 3390 398772
rect 231210 398760 231216 398772
rect 231268 398760 231274 398812
rect 3694 375980 3700 376032
rect 3752 376020 3758 376032
rect 231118 376020 231124 376032
rect 3752 375992 231124 376020
rect 3752 375980 3758 375992
rect 231118 375980 231124 375992
rect 231176 375980 231182 376032
rect 167638 374892 167644 374944
rect 167696 374932 167702 374944
rect 174630 374932 174636 374944
rect 167696 374904 174636 374932
rect 167696 374892 167702 374904
rect 174630 374892 174636 374904
rect 174688 374892 174694 374944
rect 121270 374824 121276 374876
rect 121328 374864 121334 374876
rect 170766 374864 170772 374876
rect 121328 374836 170772 374864
rect 121328 374824 121334 374836
rect 170766 374824 170772 374836
rect 170824 374824 170830 374876
rect 108390 374756 108396 374808
rect 108448 374796 108454 374808
rect 229738 374796 229744 374808
rect 108448 374768 229744 374796
rect 108448 374756 108454 374768
rect 229738 374756 229744 374768
rect 229796 374756 229802 374808
rect 131574 374688 131580 374740
rect 131632 374728 131638 374740
rect 171870 374728 171876 374740
rect 131632 374700 171876 374728
rect 131632 374688 131638 374700
rect 171870 374688 171876 374700
rect 171928 374688 171934 374740
rect 147030 374620 147036 374672
rect 147088 374660 147094 374672
rect 170398 374660 170404 374672
rect 147088 374632 170404 374660
rect 147088 374620 147094 374632
rect 170398 374620 170404 374632
rect 170456 374620 170462 374672
rect 139302 374552 139308 374604
rect 139360 374592 139366 374604
rect 170858 374592 170864 374604
rect 139360 374564 170864 374592
rect 139360 374552 139366 374564
rect 170858 374552 170864 374564
rect 170916 374552 170922 374604
rect 116118 374484 116124 374536
rect 116176 374524 116182 374536
rect 173250 374524 173256 374536
rect 116176 374496 173256 374524
rect 116176 374484 116182 374496
rect 173250 374484 173256 374496
rect 173308 374484 173314 374536
rect 110966 374416 110972 374468
rect 111024 374456 111030 374468
rect 170950 374456 170956 374468
rect 111024 374428 170956 374456
rect 111024 374416 111030 374428
rect 170950 374416 170956 374428
rect 171008 374416 171014 374468
rect 165522 374348 165528 374400
rect 165580 374388 165586 374400
rect 226978 374388 226984 374400
rect 165580 374360 226984 374388
rect 165580 374348 165586 374360
rect 226978 374348 226984 374360
rect 227036 374348 227042 374400
rect 162486 374280 162492 374332
rect 162544 374320 162550 374332
rect 228358 374320 228364 374332
rect 162544 374292 228364 374320
rect 162544 374280 162550 374292
rect 228358 374280 228364 374292
rect 228416 374280 228422 374332
rect 157334 374212 157340 374264
rect 157392 374252 157398 374264
rect 230014 374252 230020 374264
rect 157392 374224 230020 374252
rect 157392 374212 157398 374224
rect 230014 374212 230020 374224
rect 230072 374212 230078 374264
rect 128998 374144 129004 374196
rect 129056 374184 129062 374196
rect 229830 374184 229836 374196
rect 129056 374156 229836 374184
rect 129056 374144 129062 374156
rect 229830 374144 229836 374156
rect 229888 374144 229894 374196
rect 113542 374076 113548 374128
rect 113600 374116 113606 374128
rect 231210 374116 231216 374128
rect 113600 374088 231216 374116
rect 113600 374076 113606 374088
rect 231210 374076 231216 374088
rect 231268 374076 231274 374128
rect 14458 373056 14464 373108
rect 14516 373096 14522 373108
rect 165062 373096 165068 373108
rect 14516 373068 165068 373096
rect 14516 373056 14522 373068
rect 165062 373056 165068 373068
rect 165120 373096 165126 373108
rect 165522 373096 165528 373108
rect 165120 373068 165528 373096
rect 165120 373056 165126 373068
rect 165522 373056 165528 373068
rect 165580 373056 165586 373108
rect 136726 372988 136732 373040
rect 136784 373028 136790 373040
rect 170674 373028 170680 373040
rect 136784 373000 170680 373028
rect 136784 372988 136790 373000
rect 170674 372988 170680 373000
rect 170732 372988 170738 373040
rect 144454 372920 144460 372972
rect 144512 372960 144518 372972
rect 188338 372960 188344 372972
rect 144512 372932 188344 372960
rect 144512 372920 144518 372932
rect 188338 372920 188344 372932
rect 188396 372920 188402 372972
rect 126422 372852 126428 372904
rect 126480 372892 126486 372904
rect 173158 372892 173164 372904
rect 126480 372864 173164 372892
rect 126480 372852 126486 372864
rect 173158 372852 173164 372864
rect 173216 372852 173222 372904
rect 100662 372784 100668 372836
rect 100720 372824 100726 372836
rect 174538 372824 174544 372836
rect 100720 372796 174544 372824
rect 100720 372784 100726 372796
rect 174538 372784 174544 372796
rect 174596 372784 174602 372836
rect 152182 372716 152188 372768
rect 152240 372756 152246 372768
rect 231118 372756 231124 372768
rect 152240 372728 231124 372756
rect 152240 372716 152246 372728
rect 231118 372716 231124 372728
rect 231176 372716 231182 372768
rect 103238 372648 103244 372700
rect 103296 372688 103302 372700
rect 229922 372688 229928 372700
rect 103296 372660 229928 372688
rect 103296 372648 103302 372660
rect 229922 372648 229928 372660
rect 229980 372648 229986 372700
rect 149606 372580 149612 372632
rect 149664 372620 149670 372632
rect 170582 372620 170588 372632
rect 149664 372592 170588 372620
rect 149664 372580 149670 372592
rect 170582 372580 170588 372592
rect 170640 372580 170646 372632
rect 3326 372512 3332 372564
rect 3384 372552 3390 372564
rect 100018 372552 100024 372564
rect 3384 372524 100024 372552
rect 3384 372512 3390 372524
rect 100018 372512 100024 372524
rect 100076 372512 100082 372564
rect 99834 371764 99840 371816
rect 99892 371804 99898 371816
rect 99892 371776 131114 371804
rect 99892 371764 99898 371776
rect 99346 371708 109034 371736
rect 97718 371492 97724 371544
rect 97776 371532 97782 371544
rect 99346 371532 99374 371708
rect 97776 371504 99374 371532
rect 99576 371640 106274 371668
rect 97776 371492 97782 371504
rect 97810 371424 97816 371476
rect 97868 371464 97874 371476
rect 99576 371464 99604 371640
rect 106090 371560 106096 371612
rect 106148 371560 106154 371612
rect 97868 371436 99604 371464
rect 97868 371424 97874 371436
rect 106108 371328 106136 371560
rect 106246 371464 106274 371640
rect 109006 371600 109034 371708
rect 113146 371708 124076 371736
rect 113146 371600 113174 371708
rect 109006 371572 113174 371600
rect 115906 371640 121592 371668
rect 106246 371436 109034 371464
rect 109006 371396 109034 371436
rect 115906 371396 115934 371640
rect 118326 371600 118332 371612
rect 109006 371368 115934 371396
rect 117286 371572 118332 371600
rect 106108 371300 113174 371328
rect 113146 370988 113174 371300
rect 117286 370988 117314 371572
rect 118326 371560 118332 371572
rect 118384 371560 118390 371612
rect 118970 371560 118976 371612
rect 119028 371560 119034 371612
rect 119062 371560 119068 371612
rect 119120 371560 119126 371612
rect 113146 370960 117314 370988
rect 118988 370784 119016 371560
rect 119080 371396 119108 371560
rect 121564 371464 121592 371640
rect 124048 371532 124076 371708
rect 131086 371668 131114 371776
rect 155034 371696 155040 371748
rect 155092 371736 155098 371748
rect 170030 371736 170036 371748
rect 155092 371708 170036 371736
rect 155092 371696 155098 371708
rect 170030 371696 170036 371708
rect 170088 371696 170094 371748
rect 173434 371668 173440 371680
rect 131086 371640 173440 371668
rect 173434 371628 173440 371640
rect 173492 371628 173498 371680
rect 124122 371560 124128 371612
rect 124180 371600 124186 371612
rect 173342 371600 173348 371612
rect 124180 371572 173348 371600
rect 124180 371560 124186 371572
rect 173342 371560 173348 371572
rect 173400 371560 173406 371612
rect 230106 371532 230112 371544
rect 124048 371504 230112 371532
rect 230106 371492 230112 371504
rect 230164 371492 230170 371544
rect 231302 371464 231308 371476
rect 121564 371436 231308 371464
rect 231302 371424 231308 371436
rect 231360 371424 231366 371476
rect 173618 371396 173624 371408
rect 119080 371368 173624 371396
rect 173618 371356 173624 371368
rect 173676 371356 173682 371408
rect 132466 371300 133874 371328
rect 132466 371260 132494 371300
rect 131086 371232 132494 371260
rect 133846 371260 133874 371300
rect 170030 371288 170036 371340
rect 170088 371328 170094 371340
rect 231394 371328 231400 371340
rect 170088 371300 231400 371328
rect 170088 371288 170094 371300
rect 231394 371288 231400 371300
rect 231452 371288 231458 371340
rect 228450 371260 228456 371272
rect 133846 371232 228456 371260
rect 131086 371192 131114 371232
rect 228450 371220 228456 371232
rect 228508 371220 228514 371272
rect 128326 371164 131114 371192
rect 128326 370920 128354 371164
rect 126946 370892 128354 370920
rect 126946 370784 126974 370892
rect 118988 370756 126974 370784
rect 172330 368500 172336 368552
rect 172388 368540 172394 368552
rect 231578 368540 231584 368552
rect 172388 368512 231584 368540
rect 172388 368500 172394 368512
rect 231578 368500 231584 368512
rect 231636 368500 231642 368552
rect 169938 367888 169944 367940
rect 169996 367928 170002 367940
rect 170490 367928 170496 367940
rect 169996 367900 170496 367928
rect 169996 367888 170002 367900
rect 170490 367888 170496 367900
rect 170548 367888 170554 367940
rect 172330 362924 172336 362976
rect 172388 362964 172394 362976
rect 230198 362964 230204 362976
rect 172388 362936 230204 362964
rect 172388 362924 172394 362936
rect 230198 362924 230204 362936
rect 230256 362924 230262 362976
rect 172422 357416 172428 357468
rect 172480 357456 172486 357468
rect 230290 357456 230296 357468
rect 172480 357428 230296 357456
rect 172480 357416 172486 357428
rect 230290 357416 230296 357428
rect 230348 357416 230354 357468
rect 172422 354696 172428 354748
rect 172480 354736 172486 354748
rect 230382 354736 230388 354748
rect 172480 354708 230388 354736
rect 172480 354696 172486 354708
rect 230382 354696 230388 354708
rect 230440 354696 230446 354748
rect 352742 353200 352748 353252
rect 352800 353240 352806 353252
rect 580166 353240 580172 353252
rect 352800 353212 580172 353240
rect 352800 353200 352806 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 172422 351908 172428 351960
rect 172480 351948 172486 351960
rect 220078 351948 220084 351960
rect 172480 351920 220084 351948
rect 172480 351908 172486 351920
rect 220078 351908 220084 351920
rect 220136 351908 220142 351960
rect 172422 346400 172428 346452
rect 172480 346440 172486 346452
rect 224218 346440 224224 346452
rect 172480 346412 224224 346440
rect 172480 346400 172486 346412
rect 224218 346400 224224 346412
rect 224276 346400 224282 346452
rect 172422 342252 172428 342304
rect 172480 342292 172486 342304
rect 232222 342292 232228 342304
rect 172480 342264 232228 342292
rect 172480 342252 172486 342264
rect 232222 342252 232228 342264
rect 232280 342252 232286 342304
rect 172422 339464 172428 339516
rect 172480 339504 172486 339516
rect 231670 339504 231676 339516
rect 172480 339476 231676 339504
rect 172480 339464 172486 339476
rect 231670 339464 231676 339476
rect 231728 339464 231734 339516
rect 172422 336744 172428 336796
rect 172480 336784 172486 336796
rect 182818 336784 182824 336796
rect 172480 336756 182824 336784
rect 172480 336744 172486 336756
rect 182818 336744 182824 336756
rect 182876 336744 182882 336796
rect 172422 331236 172428 331288
rect 172480 331276 172486 331288
rect 231762 331276 231768 331288
rect 172480 331248 231768 331276
rect 172480 331236 172486 331248
rect 231762 331236 231768 331248
rect 231820 331236 231826 331288
rect 172422 328448 172428 328500
rect 172480 328488 172486 328500
rect 227070 328488 227076 328500
rect 172480 328460 227076 328488
rect 172480 328448 172486 328460
rect 227070 328448 227076 328460
rect 227128 328448 227134 328500
rect 356698 325592 356704 325644
rect 356756 325632 356762 325644
rect 580166 325632 580172 325644
rect 356756 325604 580172 325632
rect 356756 325592 356762 325604
rect 580166 325592 580172 325604
rect 580224 325592 580230 325644
rect 171318 322940 171324 322992
rect 171376 322980 171382 322992
rect 228542 322980 228548 322992
rect 171376 322952 228548 322980
rect 171376 322940 171382 322952
rect 228542 322940 228548 322952
rect 228600 322940 228606 322992
rect 171502 320152 171508 320204
rect 171560 320192 171566 320204
rect 231026 320192 231032 320204
rect 171560 320164 231032 320192
rect 171560 320152 171566 320164
rect 231026 320152 231032 320164
rect 231084 320152 231090 320204
rect 3326 320084 3332 320136
rect 3384 320124 3390 320136
rect 98638 320124 98644 320136
rect 3384 320096 98644 320124
rect 3384 320084 3390 320096
rect 98638 320084 98644 320096
rect 98696 320084 98702 320136
rect 171502 317432 171508 317484
rect 171560 317472 171566 317484
rect 231946 317472 231952 317484
rect 171560 317444 231952 317472
rect 171560 317432 171566 317444
rect 231946 317432 231952 317444
rect 232004 317432 232010 317484
rect 172422 314644 172428 314696
rect 172480 314684 172486 314696
rect 232130 314684 232136 314696
rect 172480 314656 232136 314684
rect 172480 314644 172486 314656
rect 232130 314644 232136 314656
rect 232188 314644 232194 314696
rect 231854 313216 231860 313268
rect 231912 313256 231918 313268
rect 232038 313256 232044 313268
rect 231912 313228 232044 313256
rect 231912 313216 231918 313228
rect 232038 313216 232044 313228
rect 232096 313216 232102 313268
rect 172422 311856 172428 311908
rect 172480 311896 172486 311908
rect 232038 311896 232044 311908
rect 172480 311868 232044 311896
rect 172480 311856 172486 311868
rect 232038 311856 232044 311868
rect 232096 311856 232102 311908
rect 172330 311244 172336 311296
rect 172388 311284 172394 311296
rect 230934 311284 230940 311296
rect 172388 311256 230940 311284
rect 172388 311244 172394 311256
rect 230934 311244 230940 311256
rect 230992 311244 230998 311296
rect 172238 311176 172244 311228
rect 172296 311216 172302 311228
rect 232222 311216 232228 311228
rect 172296 311188 232228 311216
rect 172296 311176 172302 311188
rect 232222 311176 232228 311188
rect 232280 311176 232286 311228
rect 170858 311108 170864 311160
rect 170916 311148 170922 311160
rect 232314 311148 232320 311160
rect 170916 311120 232320 311148
rect 170916 311108 170922 311120
rect 232314 311108 232320 311120
rect 232372 311108 232378 311160
rect 219406 310848 224954 310876
rect 172146 310700 172152 310752
rect 172204 310740 172210 310752
rect 219406 310740 219434 310848
rect 172204 310712 219434 310740
rect 224926 310740 224954 310848
rect 224926 310712 233740 310740
rect 172204 310700 172210 310712
rect 171962 310632 171968 310684
rect 172020 310672 172026 310684
rect 222286 310672 222292 310684
rect 172020 310644 222292 310672
rect 172020 310632 172026 310644
rect 222286 310632 222292 310644
rect 222344 310632 222350 310684
rect 225064 310644 233188 310672
rect 172054 310564 172060 310616
rect 172112 310604 172118 310616
rect 225064 310604 225092 310644
rect 233160 310616 233188 310644
rect 233712 310616 233740 310712
rect 172112 310576 225092 310604
rect 172112 310564 172118 310576
rect 232222 310564 232228 310616
rect 232280 310604 232286 310616
rect 232280 310576 233096 310604
rect 232280 310564 232286 310576
rect 231780 310508 232268 310536
rect 230198 310428 230204 310480
rect 230256 310468 230262 310480
rect 231780 310468 231808 310508
rect 230256 310440 231808 310468
rect 232240 310468 232268 310508
rect 232314 310496 232320 310548
rect 232372 310536 232378 310548
rect 232590 310536 232596 310548
rect 232372 310508 232596 310536
rect 232372 310496 232378 310508
rect 232590 310496 232596 310508
rect 232648 310496 232654 310548
rect 232958 310536 232964 310548
rect 232700 310508 232964 310536
rect 232700 310468 232728 310508
rect 232958 310496 232964 310508
rect 233016 310496 233022 310548
rect 232240 310440 232728 310468
rect 233068 310468 233096 310576
rect 233142 310564 233148 310616
rect 233200 310564 233206 310616
rect 233694 310564 233700 310616
rect 233752 310564 233758 310616
rect 233510 310468 233516 310480
rect 233068 310440 233516 310468
rect 230256 310428 230262 310440
rect 233510 310428 233516 310440
rect 233568 310428 233574 310480
rect 232222 310360 232228 310412
rect 232280 310400 232286 310412
rect 232280 310372 244274 310400
rect 232280 310360 232286 310372
rect 222286 310292 222292 310344
rect 222344 310332 222350 310344
rect 231854 310332 231860 310344
rect 222344 310304 231860 310332
rect 222344 310292 222350 310304
rect 231854 310292 231860 310304
rect 231912 310292 231918 310344
rect 232130 310292 232136 310344
rect 232188 310332 232194 310344
rect 235166 310332 235172 310344
rect 232188 310304 235172 310332
rect 232188 310292 232194 310304
rect 235166 310292 235172 310304
rect 235224 310292 235230 310344
rect 244246 310332 244274 310372
rect 248322 310332 248328 310344
rect 244246 310304 248328 310332
rect 248322 310292 248328 310304
rect 248380 310292 248386 310344
rect 232038 310224 232044 310276
rect 232096 310264 232102 310276
rect 235902 310264 235908 310276
rect 232096 310236 235908 310264
rect 232096 310224 232102 310236
rect 235902 310224 235908 310236
rect 235960 310224 235966 310276
rect 230382 310156 230388 310208
rect 230440 310196 230446 310208
rect 238202 310196 238208 310208
rect 230440 310168 238208 310196
rect 230440 310156 230446 310168
rect 238202 310156 238208 310168
rect 238260 310156 238266 310208
rect 230934 310088 230940 310140
rect 230992 310128 230998 310140
rect 232038 310128 232044 310140
rect 230992 310100 232044 310128
rect 230992 310088 230998 310100
rect 232038 310088 232044 310100
rect 232096 310088 232102 310140
rect 231762 310020 231768 310072
rect 231820 310060 231826 310072
rect 241054 310060 241060 310072
rect 231820 310032 241060 310060
rect 231820 310020 231826 310032
rect 241054 310020 241060 310032
rect 241112 310020 241118 310072
rect 172422 309952 172428 310004
rect 172480 309992 172486 310004
rect 235534 309992 235540 310004
rect 172480 309964 235540 309992
rect 172480 309952 172486 309964
rect 235534 309952 235540 309964
rect 235592 309952 235598 310004
rect 231670 309612 231676 309664
rect 231728 309652 231734 309664
rect 244734 309652 244740 309664
rect 231728 309624 244740 309652
rect 231728 309612 231734 309624
rect 244734 309612 244740 309624
rect 244792 309612 244798 309664
rect 228542 309544 228548 309596
rect 228600 309584 228606 309596
rect 238938 309584 238944 309596
rect 228600 309556 238944 309584
rect 228600 309544 228606 309556
rect 238938 309544 238944 309556
rect 238996 309544 239002 309596
rect 356790 309584 356796 309596
rect 331186 309556 356796 309584
rect 230290 309476 230296 309528
rect 230348 309516 230354 309528
rect 242066 309516 242072 309528
rect 230348 309488 242072 309516
rect 230348 309476 230354 309488
rect 242066 309476 242072 309488
rect 242124 309476 242130 309528
rect 297174 309476 297180 309528
rect 297232 309516 297238 309528
rect 331186 309516 331214 309556
rect 356790 309544 356796 309556
rect 356848 309544 356854 309596
rect 297232 309488 331214 309516
rect 297232 309476 297238 309488
rect 231578 309408 231584 309460
rect 231636 309448 231642 309460
rect 247770 309448 247776 309460
rect 231636 309420 247776 309448
rect 231636 309408 231642 309420
rect 247770 309408 247776 309420
rect 247828 309408 247834 309460
rect 297358 309408 297364 309460
rect 297416 309448 297422 309460
rect 356698 309448 356704 309460
rect 297416 309420 356704 309448
rect 297416 309408 297422 309420
rect 356698 309408 356704 309420
rect 356756 309408 356762 309460
rect 231026 309340 231032 309392
rect 231084 309380 231090 309392
rect 248506 309380 248512 309392
rect 231084 309352 248512 309380
rect 231084 309340 231090 309352
rect 248506 309340 248512 309352
rect 248564 309340 248570 309392
rect 298646 309340 298652 309392
rect 298704 309380 298710 309392
rect 358814 309380 358820 309392
rect 298704 309352 358820 309380
rect 298704 309340 298710 309352
rect 358814 309340 358820 309352
rect 358872 309340 358878 309392
rect 231946 309272 231952 309324
rect 232004 309312 232010 309324
rect 251358 309312 251364 309324
rect 232004 309284 251364 309312
rect 232004 309272 232010 309284
rect 251358 309272 251364 309284
rect 251416 309272 251422 309324
rect 298278 309272 298284 309324
rect 298336 309312 298342 309324
rect 361574 309312 361580 309324
rect 298336 309284 361580 309312
rect 298336 309272 298342 309284
rect 361574 309272 361580 309284
rect 361632 309272 361638 309324
rect 182818 309204 182824 309256
rect 182876 309244 182882 309256
rect 238386 309244 238392 309256
rect 182876 309216 238392 309244
rect 182876 309204 182882 309216
rect 238386 309204 238392 309216
rect 238444 309204 238450 309256
rect 297910 309204 297916 309256
rect 297968 309244 297974 309256
rect 360286 309244 360292 309256
rect 297968 309216 360292 309244
rect 297968 309204 297974 309216
rect 360286 309204 360292 309216
rect 360344 309204 360350 309256
rect 170490 309136 170496 309188
rect 170548 309176 170554 309188
rect 233970 309176 233976 309188
rect 170548 309148 233976 309176
rect 170548 309136 170554 309148
rect 233970 309136 233976 309148
rect 234028 309136 234034 309188
rect 299198 309136 299204 309188
rect 299256 309176 299262 309188
rect 367094 309176 367100 309188
rect 299256 309148 367100 309176
rect 299256 309136 299262 309148
rect 367094 309136 367100 309148
rect 367152 309136 367158 309188
rect 171778 309068 171784 309120
rect 171836 309108 171842 309120
rect 232406 309108 232412 309120
rect 171836 309080 232412 309108
rect 171836 309068 171842 309080
rect 232406 309068 232412 309080
rect 232464 309068 232470 309120
rect 233694 309068 233700 309120
rect 233752 309108 233758 309120
rect 238018 309108 238024 309120
rect 233752 309080 238024 309108
rect 233752 309068 233758 309080
rect 238018 309068 238024 309080
rect 238076 309068 238082 309120
rect 347222 309068 347228 309120
rect 347280 309108 347286 309120
rect 363598 309108 363604 309120
rect 347280 309080 363604 309108
rect 347280 309068 347286 309080
rect 363598 309068 363604 309080
rect 363656 309068 363662 309120
rect 230106 309000 230112 309052
rect 230164 309040 230170 309052
rect 233418 309040 233424 309052
rect 230164 309012 233424 309040
rect 230164 309000 230170 309012
rect 233418 309000 233424 309012
rect 233476 309000 233482 309052
rect 346854 309000 346860 309052
rect 346912 309040 346918 309052
rect 364610 309040 364616 309052
rect 346912 309012 364616 309040
rect 346912 309000 346918 309012
rect 364610 309000 364616 309012
rect 364668 309000 364674 309052
rect 233142 308932 233148 308984
rect 233200 308972 233206 308984
rect 240870 308972 240876 308984
rect 233200 308944 240876 308972
rect 233200 308932 233206 308944
rect 240870 308932 240876 308944
rect 240928 308932 240934 308984
rect 261202 308932 261208 308984
rect 261260 308972 261266 308984
rect 261478 308972 261484 308984
rect 261260 308944 261484 308972
rect 261260 308932 261266 308944
rect 261478 308932 261484 308944
rect 261536 308932 261542 308984
rect 346486 308932 346492 308984
rect 346544 308972 346550 308984
rect 364978 308972 364984 308984
rect 346544 308944 364984 308972
rect 346544 308932 346550 308944
rect 364978 308932 364984 308944
rect 365036 308932 365042 308984
rect 229830 308864 229836 308916
rect 229888 308904 229894 308916
rect 241422 308904 241428 308916
rect 229888 308876 241428 308904
rect 229888 308864 229894 308876
rect 241422 308864 241428 308876
rect 241480 308864 241486 308916
rect 345014 308864 345020 308916
rect 345072 308904 345078 308916
rect 364334 308904 364340 308916
rect 345072 308876 364340 308904
rect 345072 308864 345078 308876
rect 364334 308864 364340 308876
rect 364392 308864 364398 308916
rect 231394 308796 231400 308848
rect 231452 308836 231458 308848
rect 239122 308836 239128 308848
rect 231452 308808 239128 308836
rect 231452 308796 231458 308808
rect 239122 308796 239128 308808
rect 239180 308796 239186 308848
rect 249058 308836 249064 308848
rect 239324 308808 249064 308836
rect 188338 308728 188344 308780
rect 188396 308768 188402 308780
rect 237650 308768 237656 308780
rect 188396 308740 237656 308768
rect 188396 308728 188402 308740
rect 237650 308728 237656 308740
rect 237708 308728 237714 308780
rect 228450 308660 228456 308712
rect 228508 308700 228514 308712
rect 239324 308700 239352 308808
rect 249058 308796 249064 308808
rect 249116 308796 249122 308848
rect 345382 308796 345388 308848
rect 345440 308836 345446 308848
rect 364518 308836 364524 308848
rect 345440 308808 364524 308836
rect 345440 308796 345446 308808
rect 364518 308796 364524 308808
rect 364576 308796 364582 308848
rect 228508 308672 239352 308700
rect 239508 308740 241514 308768
rect 228508 308660 228514 308672
rect 170582 308592 170588 308644
rect 170640 308632 170646 308644
rect 239508 308632 239536 308740
rect 170640 308604 239536 308632
rect 241486 308632 241514 308740
rect 246942 308728 246948 308780
rect 247000 308768 247006 308780
rect 258074 308768 258080 308780
rect 247000 308740 258080 308768
rect 247000 308728 247006 308740
rect 258074 308728 258080 308740
rect 258132 308728 258138 308780
rect 346118 308728 346124 308780
rect 346176 308768 346182 308780
rect 364886 308768 364892 308780
rect 346176 308740 364892 308768
rect 346176 308728 346182 308740
rect 364886 308728 364892 308740
rect 364944 308728 364950 308780
rect 250898 308660 250904 308712
rect 250956 308700 250962 308712
rect 250956 308672 253934 308700
rect 250956 308660 250962 308672
rect 245654 308632 245660 308644
rect 241486 308604 245660 308632
rect 170640 308592 170646 308604
rect 245654 308592 245660 308604
rect 245712 308592 245718 308644
rect 253906 308632 253934 308672
rect 305178 308660 305184 308712
rect 305236 308700 305242 308712
rect 305454 308700 305460 308712
rect 305236 308672 305460 308700
rect 305236 308660 305242 308672
rect 305454 308660 305460 308672
rect 305512 308660 305518 308712
rect 348234 308660 348240 308712
rect 348292 308700 348298 308712
rect 352466 308700 352472 308712
rect 348292 308672 352472 308700
rect 348292 308660 348298 308672
rect 352466 308660 352472 308672
rect 352524 308660 352530 308712
rect 352742 308660 352748 308712
rect 352800 308700 352806 308712
rect 364702 308700 364708 308712
rect 352800 308672 364708 308700
rect 352800 308660 352806 308672
rect 364702 308660 364708 308672
rect 364760 308660 364766 308712
rect 267642 308632 267648 308644
rect 253906 308604 267648 308632
rect 267642 308592 267648 308604
rect 267700 308592 267706 308644
rect 314654 308592 314660 308644
rect 314712 308632 314718 308644
rect 315850 308632 315856 308644
rect 314712 308604 315856 308632
rect 314712 308592 314718 308604
rect 315850 308592 315856 308604
rect 315908 308592 315914 308644
rect 316218 308592 316224 308644
rect 316276 308632 316282 308644
rect 318242 308632 318248 308644
rect 316276 308604 318248 308632
rect 316276 308592 316282 308604
rect 318242 308592 318248 308604
rect 318300 308592 318306 308644
rect 320358 308592 320364 308644
rect 320416 308632 320422 308644
rect 320634 308632 320640 308644
rect 320416 308604 320640 308632
rect 320416 308592 320422 308604
rect 320634 308592 320640 308604
rect 320692 308592 320698 308644
rect 344738 308592 344744 308644
rect 344796 308632 344802 308644
rect 364426 308632 364432 308644
rect 344796 308604 364432 308632
rect 344796 308592 344802 308604
rect 364426 308592 364432 308604
rect 364484 308592 364490 308644
rect 173158 308524 173164 308576
rect 173216 308564 173222 308576
rect 243722 308564 243728 308576
rect 173216 308536 243728 308564
rect 173216 308524 173222 308536
rect 243722 308524 243728 308536
rect 243780 308524 243786 308576
rect 252278 308524 252284 308576
rect 252336 308564 252342 308576
rect 252336 308536 253934 308564
rect 252336 308524 252342 308536
rect 236638 308496 236644 308508
rect 219406 308468 236644 308496
rect 170674 308388 170680 308440
rect 170732 308428 170738 308440
rect 219406 308428 219434 308468
rect 236638 308456 236644 308468
rect 236696 308456 236702 308508
rect 253906 308496 253934 308536
rect 270218 308524 270224 308576
rect 270276 308564 270282 308576
rect 275278 308564 275284 308576
rect 270276 308536 275284 308564
rect 270276 308524 270282 308536
rect 275278 308524 275284 308536
rect 275336 308524 275342 308576
rect 294598 308524 294604 308576
rect 294656 308564 294662 308576
rect 294782 308564 294788 308576
rect 294656 308536 294788 308564
rect 294656 308524 294662 308536
rect 294782 308524 294788 308536
rect 294840 308524 294846 308576
rect 313274 308524 313280 308576
rect 313332 308564 313338 308576
rect 314194 308564 314200 308576
rect 313332 308536 314200 308564
rect 313332 308524 313338 308536
rect 314194 308524 314200 308536
rect 314252 308524 314258 308576
rect 314746 308524 314752 308576
rect 314804 308564 314810 308576
rect 315206 308564 315212 308576
rect 314804 308536 315212 308564
rect 314804 308524 314810 308536
rect 315206 308524 315212 308536
rect 315264 308524 315270 308576
rect 316126 308524 316132 308576
rect 316184 308564 316190 308576
rect 316494 308564 316500 308576
rect 316184 308536 316500 308564
rect 316184 308524 316190 308536
rect 316494 308524 316500 308536
rect 316552 308524 316558 308576
rect 317506 308524 317512 308576
rect 317564 308564 317570 308576
rect 317966 308564 317972 308576
rect 317564 308536 317972 308564
rect 317564 308524 317570 308536
rect 317966 308524 317972 308536
rect 318024 308524 318030 308576
rect 339402 308524 339408 308576
rect 339460 308564 339466 308576
rect 364794 308564 364800 308576
rect 339460 308536 364800 308564
rect 339460 308524 339466 308536
rect 364794 308524 364800 308536
rect 364852 308524 364858 308576
rect 268654 308496 268660 308508
rect 253906 308468 268660 308496
rect 268654 308456 268660 308468
rect 268712 308456 268718 308508
rect 304442 308456 304448 308508
rect 304500 308496 304506 308508
rect 347130 308496 347136 308508
rect 304500 308468 347136 308496
rect 304500 308456 304506 308468
rect 347130 308456 347136 308468
rect 347188 308456 347194 308508
rect 350718 308456 350724 308508
rect 350776 308456 350782 308508
rect 352466 308456 352472 308508
rect 352524 308496 352530 308508
rect 367370 308496 367376 308508
rect 352524 308468 367376 308496
rect 352524 308456 352530 308468
rect 367370 308456 367376 308468
rect 367428 308456 367434 308508
rect 170732 308400 219434 308428
rect 170732 308388 170738 308400
rect 231118 308388 231124 308440
rect 231176 308428 231182 308440
rect 239582 308428 239588 308440
rect 231176 308400 239588 308428
rect 231176 308388 231182 308400
rect 239582 308388 239588 308400
rect 239640 308388 239646 308440
rect 269206 308428 269212 308440
rect 253906 308400 269212 308428
rect 173342 308320 173348 308372
rect 173400 308360 173406 308372
rect 241606 308360 241612 308372
rect 173400 308332 241612 308360
rect 173400 308320 173406 308332
rect 241606 308320 241612 308332
rect 241664 308320 241670 308372
rect 243538 308184 243544 308236
rect 243596 308224 243602 308236
rect 251818 308224 251824 308236
rect 243596 308196 251824 308224
rect 243596 308184 243602 308196
rect 251818 308184 251824 308196
rect 251876 308184 251882 308236
rect 232038 308116 232044 308168
rect 232096 308156 232102 308168
rect 243446 308156 243452 308168
rect 232096 308128 243452 308156
rect 232096 308116 232102 308128
rect 243446 308116 243452 308128
rect 243504 308116 243510 308168
rect 246850 308116 246856 308168
rect 246908 308156 246914 308168
rect 252738 308156 252744 308168
rect 246908 308128 252744 308156
rect 246908 308116 246914 308128
rect 252738 308116 252744 308128
rect 252796 308116 252802 308168
rect 231854 308048 231860 308100
rect 231912 308088 231918 308100
rect 246390 308088 246396 308100
rect 231912 308060 246396 308088
rect 231912 308048 231918 308060
rect 246390 308048 246396 308060
rect 246448 308048 246454 308100
rect 250530 308048 250536 308100
rect 250588 308088 250594 308100
rect 253906 308088 253934 308400
rect 269206 308388 269212 308400
rect 269264 308388 269270 308440
rect 295978 308388 295984 308440
rect 296036 308428 296042 308440
rect 349890 308428 349896 308440
rect 296036 308400 349896 308428
rect 296036 308388 296042 308400
rect 349890 308388 349896 308400
rect 349948 308388 349954 308440
rect 350736 308428 350764 308456
rect 367278 308428 367284 308440
rect 350736 308400 367284 308428
rect 367278 308388 367284 308400
rect 367336 308388 367342 308440
rect 312354 308320 312360 308372
rect 312412 308360 312418 308372
rect 313182 308360 313188 308372
rect 312412 308332 313188 308360
rect 312412 308320 312418 308332
rect 313182 308320 313188 308332
rect 313240 308320 313246 308372
rect 313642 308320 313648 308372
rect 313700 308360 313706 308372
rect 314010 308360 314016 308372
rect 313700 308332 314016 308360
rect 313700 308320 313706 308332
rect 314010 308320 314016 308332
rect 314068 308320 314074 308372
rect 314838 308320 314844 308372
rect 314896 308360 314902 308372
rect 315298 308360 315304 308372
rect 314896 308332 315304 308360
rect 314896 308320 314902 308332
rect 315298 308320 315304 308332
rect 315356 308320 315362 308372
rect 316402 308320 316408 308372
rect 316460 308360 316466 308372
rect 317046 308360 317052 308372
rect 316460 308332 317052 308360
rect 316460 308320 316466 308332
rect 317046 308320 317052 308332
rect 317104 308320 317110 308372
rect 317414 308320 317420 308372
rect 317472 308360 317478 308372
rect 317690 308360 317696 308372
rect 317472 308332 317696 308360
rect 317472 308320 317478 308332
rect 317690 308320 317696 308332
rect 317748 308320 317754 308372
rect 317874 308320 317880 308372
rect 317932 308360 317938 308372
rect 318334 308360 318340 308372
rect 317932 308332 318340 308360
rect 317932 308320 317938 308332
rect 318334 308320 318340 308332
rect 318392 308320 318398 308372
rect 318794 308320 318800 308372
rect 318852 308360 318858 308372
rect 319254 308360 319260 308372
rect 318852 308332 319260 308360
rect 318852 308320 318858 308332
rect 319254 308320 319260 308332
rect 319312 308320 319318 308372
rect 319438 308320 319444 308372
rect 319496 308360 319502 308372
rect 319898 308360 319904 308372
rect 319496 308332 319904 308360
rect 319496 308320 319502 308332
rect 319898 308320 319904 308332
rect 319956 308320 319962 308372
rect 320542 308320 320548 308372
rect 320600 308360 320606 308372
rect 321094 308360 321100 308372
rect 320600 308332 321100 308360
rect 320600 308320 320606 308332
rect 321094 308320 321100 308332
rect 321152 308320 321158 308372
rect 340966 308320 340972 308372
rect 341024 308360 341030 308372
rect 343358 308360 343364 308372
rect 341024 308332 343364 308360
rect 341024 308320 341030 308332
rect 343358 308320 343364 308332
rect 343416 308320 343422 308372
rect 344370 308320 344376 308372
rect 344428 308360 344434 308372
rect 360930 308360 360936 308372
rect 344428 308332 360936 308360
rect 344428 308320 344434 308332
rect 360930 308320 360936 308332
rect 360988 308320 360994 308372
rect 273162 308252 273168 308304
rect 273220 308292 273226 308304
rect 273714 308292 273720 308304
rect 273220 308264 273720 308292
rect 273220 308252 273226 308264
rect 273714 308252 273720 308264
rect 273772 308252 273778 308304
rect 311894 308252 311900 308304
rect 311952 308292 311958 308304
rect 312630 308292 312636 308304
rect 311952 308264 312636 308292
rect 311952 308252 311958 308264
rect 312630 308252 312636 308264
rect 312688 308252 312694 308304
rect 313366 308252 313372 308304
rect 313424 308292 313430 308304
rect 313918 308292 313924 308304
rect 313424 308264 313924 308292
rect 313424 308252 313430 308264
rect 313918 308252 313924 308264
rect 313976 308252 313982 308304
rect 314930 308252 314936 308304
rect 314988 308292 314994 308304
rect 315114 308292 315120 308304
rect 314988 308264 315120 308292
rect 314988 308252 314994 308264
rect 315114 308252 315120 308264
rect 315172 308252 315178 308304
rect 316310 308252 316316 308304
rect 316368 308292 316374 308304
rect 317230 308292 317236 308304
rect 316368 308264 317236 308292
rect 316368 308252 316374 308264
rect 317230 308252 317236 308264
rect 317288 308252 317294 308304
rect 319162 308292 319168 308304
rect 318812 308264 319168 308292
rect 318812 308236 318840 308264
rect 319162 308252 319168 308264
rect 319220 308252 319226 308304
rect 320174 308252 320180 308304
rect 320232 308292 320238 308304
rect 321278 308292 321284 308304
rect 320232 308264 321284 308292
rect 320232 308252 320238 308264
rect 321278 308252 321284 308264
rect 321336 308252 321342 308304
rect 350534 308252 350540 308304
rect 350592 308292 350598 308304
rect 350902 308292 350908 308304
rect 350592 308264 350908 308292
rect 350592 308252 350598 308264
rect 350902 308252 350908 308264
rect 350960 308252 350966 308304
rect 363506 308292 363512 308304
rect 351932 308264 363512 308292
rect 312078 308184 312084 308236
rect 312136 308224 312142 308236
rect 312538 308224 312544 308236
rect 312136 308196 312544 308224
rect 312136 308184 312142 308196
rect 312538 308184 312544 308196
rect 312596 308184 312602 308236
rect 313550 308184 313556 308236
rect 313608 308224 313614 308236
rect 314562 308224 314568 308236
rect 313608 308196 314568 308224
rect 313608 308184 313614 308196
rect 314562 308184 314568 308196
rect 314620 308184 314626 308236
rect 314746 308184 314752 308236
rect 314804 308224 314810 308236
rect 315482 308224 315488 308236
rect 314804 308196 315488 308224
rect 314804 308184 314810 308196
rect 315482 308184 315488 308196
rect 315540 308184 315546 308236
rect 316034 308184 316040 308236
rect 316092 308224 316098 308236
rect 316494 308224 316500 308236
rect 316092 308196 316500 308224
rect 316092 308184 316098 308196
rect 316494 308184 316500 308196
rect 316552 308184 316558 308236
rect 317414 308184 317420 308236
rect 317472 308224 317478 308236
rect 318518 308224 318524 308236
rect 317472 308196 318524 308224
rect 317472 308184 317478 308196
rect 318518 308184 318524 308196
rect 318576 308184 318582 308236
rect 318794 308184 318800 308236
rect 318852 308184 318858 308236
rect 350718 308184 350724 308236
rect 350776 308224 350782 308236
rect 351270 308224 351276 308236
rect 350776 308196 351276 308224
rect 350776 308184 350782 308196
rect 351270 308184 351276 308196
rect 351328 308184 351334 308236
rect 312170 308116 312176 308168
rect 312228 308156 312234 308168
rect 312998 308156 313004 308168
rect 312228 308128 313004 308156
rect 312228 308116 312234 308128
rect 312998 308116 313004 308128
rect 313056 308116 313062 308168
rect 313366 308116 313372 308168
rect 313424 308156 313430 308168
rect 314378 308156 314384 308168
rect 313424 308128 314384 308156
rect 313424 308116 313430 308128
rect 314378 308116 314384 308128
rect 314436 308116 314442 308168
rect 314930 308116 314936 308168
rect 314988 308156 314994 308168
rect 315666 308156 315672 308168
rect 314988 308128 315672 308156
rect 314988 308116 314994 308128
rect 315666 308116 315672 308128
rect 315724 308116 315730 308168
rect 319162 308116 319168 308168
rect 319220 308156 319226 308168
rect 319714 308156 319720 308168
rect 319220 308128 319720 308156
rect 319220 308116 319226 308128
rect 319714 308116 319720 308128
rect 319772 308116 319778 308168
rect 350902 308116 350908 308168
rect 350960 308156 350966 308168
rect 351822 308156 351828 308168
rect 350960 308128 351828 308156
rect 350960 308116 350966 308128
rect 351822 308116 351828 308128
rect 351880 308116 351886 308168
rect 250588 308060 253934 308088
rect 250588 308048 250594 308060
rect 318978 308048 318984 308100
rect 319036 308088 319042 308100
rect 319530 308088 319536 308100
rect 319036 308060 319536 308088
rect 319036 308048 319042 308060
rect 319530 308048 319536 308060
rect 319588 308048 319594 308100
rect 347866 308048 347872 308100
rect 347924 308088 347930 308100
rect 351932 308088 351960 308264
rect 363506 308252 363512 308264
rect 363564 308252 363570 308304
rect 347924 308060 351960 308088
rect 347924 308048 347930 308060
rect 250714 307980 250720 308032
rect 250772 308020 250778 308032
rect 254670 308020 254676 308032
rect 250772 307992 254676 308020
rect 250772 307980 250778 307992
rect 254670 307980 254676 307992
rect 254728 307980 254734 308032
rect 275278 307980 275284 308032
rect 275336 308020 275342 308032
rect 280338 308020 280344 308032
rect 275336 307992 280344 308020
rect 275336 307980 275342 307992
rect 280338 307980 280344 307992
rect 280396 307980 280402 308032
rect 311250 307980 311256 308032
rect 311308 308020 311314 308032
rect 312630 308020 312636 308032
rect 311308 307992 312636 308020
rect 311308 307980 311314 307992
rect 312630 307980 312636 307992
rect 312688 307980 312694 308032
rect 316126 307980 316132 308032
rect 316184 308020 316190 308032
rect 316862 308020 316868 308032
rect 316184 307992 316868 308020
rect 316184 307980 316190 307992
rect 316862 307980 316868 307992
rect 316920 307980 316926 308032
rect 319070 307980 319076 308032
rect 319128 308020 319134 308032
rect 320082 308020 320088 308032
rect 319128 307992 320088 308020
rect 319128 307980 319134 307992
rect 320082 307980 320088 307992
rect 320140 307980 320146 308032
rect 249058 307912 249064 307964
rect 249116 307952 249122 307964
rect 255958 307952 255964 307964
rect 249116 307924 255964 307952
rect 249116 307912 249122 307924
rect 255958 307912 255964 307924
rect 256016 307912 256022 307964
rect 270586 307912 270592 307964
rect 270644 307952 270650 307964
rect 271138 307952 271144 307964
rect 270644 307924 271144 307952
rect 270644 307912 270650 307924
rect 271138 307912 271144 307924
rect 271196 307912 271202 307964
rect 278590 307952 278596 307964
rect 273226 307924 278596 307952
rect 242802 307844 242808 307896
rect 242860 307884 242866 307896
rect 250990 307884 250996 307896
rect 242860 307856 250996 307884
rect 242860 307844 242866 307856
rect 250990 307844 250996 307856
rect 251048 307844 251054 307896
rect 257430 307844 257436 307896
rect 257488 307884 257494 307896
rect 263410 307884 263416 307896
rect 257488 307856 263416 307884
rect 257488 307844 257494 307856
rect 263410 307844 263416 307856
rect 263468 307844 263474 307896
rect 272518 307844 272524 307896
rect 272576 307884 272582 307896
rect 273226 307884 273254 307924
rect 278590 307912 278596 307924
rect 278648 307912 278654 307964
rect 318610 307912 318616 307964
rect 318668 307952 318674 307964
rect 319530 307952 319536 307964
rect 318668 307924 319536 307952
rect 318668 307912 318674 307924
rect 319530 307912 319536 307924
rect 319588 307912 319594 307964
rect 330018 307912 330024 307964
rect 330076 307952 330082 307964
rect 331858 307952 331864 307964
rect 330076 307924 331864 307952
rect 330076 307912 330082 307924
rect 331858 307912 331864 307924
rect 331916 307912 331922 307964
rect 345750 307912 345756 307964
rect 345808 307952 345814 307964
rect 352742 307952 352748 307964
rect 345808 307924 352748 307952
rect 345808 307912 345814 307924
rect 352742 307912 352748 307924
rect 352800 307912 352806 307964
rect 272576 307856 273254 307884
rect 272576 307844 272582 307856
rect 278314 307844 278320 307896
rect 278372 307884 278378 307896
rect 280890 307884 280896 307896
rect 278372 307856 280896 307884
rect 278372 307844 278378 307856
rect 280890 307844 280896 307856
rect 280948 307844 280954 307896
rect 325786 307844 325792 307896
rect 325844 307884 325850 307896
rect 329006 307884 329012 307896
rect 325844 307856 329012 307884
rect 325844 307844 325850 307856
rect 329006 307844 329012 307856
rect 329064 307844 329070 307896
rect 347498 307844 347504 307896
rect 347556 307884 347562 307896
rect 359642 307884 359648 307896
rect 347556 307856 359648 307884
rect 347556 307844 347562 307856
rect 359642 307844 359648 307856
rect 359700 307844 359706 307896
rect 237374 307776 237380 307828
rect 237432 307816 237438 307828
rect 240686 307816 240692 307828
rect 237432 307788 240692 307816
rect 237432 307776 237438 307788
rect 240686 307776 240692 307788
rect 240744 307776 240750 307828
rect 247034 307776 247040 307828
rect 247092 307816 247098 307828
rect 250438 307816 250444 307828
rect 247092 307788 250444 307816
rect 247092 307776 247098 307788
rect 250438 307776 250444 307788
rect 250496 307776 250502 307828
rect 251818 307776 251824 307828
rect 251876 307816 251882 307828
rect 259086 307816 259092 307828
rect 251876 307788 259092 307816
rect 251876 307776 251882 307788
rect 259086 307776 259092 307788
rect 259144 307776 259150 307828
rect 270034 307776 270040 307828
rect 270092 307816 270098 307828
rect 270494 307816 270500 307828
rect 270092 307788 270500 307816
rect 270092 307776 270098 307788
rect 270494 307776 270500 307788
rect 270552 307776 270558 307828
rect 275370 307776 275376 307828
rect 275428 307816 275434 307828
rect 277394 307816 277400 307828
rect 275428 307788 277400 307816
rect 275428 307776 275434 307788
rect 277394 307776 277400 307788
rect 277452 307776 277458 307828
rect 278130 307776 278136 307828
rect 278188 307816 278194 307828
rect 278774 307816 278780 307828
rect 278188 307788 278780 307816
rect 278188 307776 278194 307788
rect 278774 307776 278780 307788
rect 278832 307776 278838 307828
rect 306926 307776 306932 307828
rect 306984 307816 306990 307828
rect 308674 307816 308680 307828
rect 306984 307788 308680 307816
rect 306984 307776 306990 307788
rect 308674 307776 308680 307788
rect 308732 307776 308738 307828
rect 309042 307776 309048 307828
rect 309100 307816 309106 307828
rect 310054 307816 310060 307828
rect 309100 307788 310060 307816
rect 309100 307776 309106 307788
rect 310054 307776 310060 307788
rect 310112 307776 310118 307828
rect 321830 307776 321836 307828
rect 321888 307816 321894 307828
rect 323670 307816 323676 307828
rect 321888 307788 323676 307816
rect 321888 307776 321894 307788
rect 323670 307776 323676 307788
rect 323728 307776 323734 307828
rect 324130 307776 324136 307828
rect 324188 307816 324194 307828
rect 325142 307816 325148 307828
rect 324188 307788 325148 307816
rect 324188 307776 324194 307788
rect 325142 307776 325148 307788
rect 325200 307776 325206 307828
rect 325234 307776 325240 307828
rect 325292 307816 325298 307828
rect 327810 307816 327816 307828
rect 325292 307788 327816 307816
rect 325292 307776 325298 307788
rect 327810 307776 327816 307788
rect 327868 307776 327874 307828
rect 328362 307776 328368 307828
rect 328420 307816 328426 307828
rect 329374 307816 329380 307828
rect 328420 307788 329380 307816
rect 328420 307776 328426 307788
rect 329374 307776 329380 307788
rect 329432 307776 329438 307828
rect 331214 307776 331220 307828
rect 331272 307816 331278 307828
rect 333422 307816 333428 307828
rect 331272 307788 333428 307816
rect 331272 307776 331278 307788
rect 333422 307776 333428 307788
rect 333480 307776 333486 307828
rect 341610 307776 341616 307828
rect 341668 307816 341674 307828
rect 342438 307816 342444 307828
rect 341668 307788 342444 307816
rect 341668 307776 341674 307788
rect 342438 307776 342444 307788
rect 342496 307776 342502 307828
rect 229738 307708 229744 307760
rect 229796 307748 229802 307760
rect 243906 307748 243912 307760
rect 229796 307720 243912 307748
rect 229796 307708 229802 307720
rect 243906 307708 243912 307720
rect 243964 307708 243970 307760
rect 227070 307640 227076 307692
rect 227128 307680 227134 307692
rect 241238 307680 241244 307692
rect 227128 307652 241244 307680
rect 227128 307640 227134 307652
rect 241238 307640 241244 307652
rect 241296 307640 241302 307692
rect 172422 307572 172428 307624
rect 172480 307612 172486 307624
rect 245838 307612 245844 307624
rect 172480 307584 245844 307612
rect 172480 307572 172486 307584
rect 245838 307572 245844 307584
rect 245896 307572 245902 307624
rect 220078 307504 220084 307556
rect 220136 307544 220142 307556
rect 242710 307544 242716 307556
rect 220136 307516 242716 307544
rect 220136 307504 220142 307516
rect 242710 307504 242716 307516
rect 242768 307504 242774 307556
rect 228358 307436 228364 307488
rect 228416 307476 228422 307488
rect 248690 307476 248696 307488
rect 228416 307448 248696 307476
rect 228416 307436 228422 307448
rect 248690 307436 248696 307448
rect 248748 307436 248754 307488
rect 224218 307368 224224 307420
rect 224276 307408 224282 307420
rect 241790 307408 241796 307420
rect 224276 307380 241796 307408
rect 224276 307368 224282 307380
rect 241790 307368 241796 307380
rect 241848 307368 241854 307420
rect 170398 307300 170404 307352
rect 170456 307340 170462 307352
rect 249150 307340 249156 307352
rect 170456 307312 249156 307340
rect 170456 307300 170462 307312
rect 249150 307300 249156 307312
rect 249208 307300 249214 307352
rect 170490 307232 170496 307284
rect 170548 307272 170554 307284
rect 236822 307272 236828 307284
rect 170548 307244 236828 307272
rect 170548 307232 170554 307244
rect 236822 307232 236828 307244
rect 236880 307232 236886 307284
rect 323302 307232 323308 307284
rect 323360 307272 323366 307284
rect 323486 307272 323492 307284
rect 323360 307244 323492 307272
rect 323360 307232 323366 307244
rect 323486 307232 323492 307244
rect 323544 307232 323550 307284
rect 215202 307164 215208 307216
rect 215260 307204 215266 307216
rect 290458 307204 290464 307216
rect 215260 307176 290464 307204
rect 215260 307164 215266 307176
rect 290458 307164 290464 307176
rect 290516 307164 290522 307216
rect 316678 307164 316684 307216
rect 316736 307204 316742 307216
rect 437474 307204 437480 307216
rect 316736 307176 437480 307204
rect 316736 307164 316742 307176
rect 437474 307164 437480 307176
rect 437532 307164 437538 307216
rect 210970 307096 210976 307148
rect 211028 307136 211034 307148
rect 339954 307136 339960 307148
rect 211028 307108 339960 307136
rect 211028 307096 211034 307108
rect 339954 307096 339960 307108
rect 340012 307096 340018 307148
rect 350626 307096 350632 307148
rect 350684 307136 350690 307148
rect 351638 307136 351644 307148
rect 350684 307108 351644 307136
rect 350684 307096 350690 307108
rect 351638 307096 351644 307108
rect 351696 307096 351702 307148
rect 195974 307028 195980 307080
rect 196032 307068 196038 307080
rect 280522 307068 280528 307080
rect 196032 307040 280528 307068
rect 196032 307028 196038 307040
rect 280522 307028 280528 307040
rect 280580 307028 280586 307080
rect 326246 307028 326252 307080
rect 326304 307068 326310 307080
rect 500954 307068 500960 307080
rect 326304 307040 500960 307068
rect 326304 307028 326310 307040
rect 500954 307028 500960 307040
rect 501012 307028 501018 307080
rect 171870 306960 171876 307012
rect 171928 307000 171934 307012
rect 171928 306972 234614 307000
rect 171928 306960 171934 306972
rect 234586 306932 234614 306972
rect 251542 306960 251548 307012
rect 251600 306960 251606 307012
rect 269390 306960 269396 307012
rect 269448 307000 269454 307012
rect 269666 307000 269672 307012
rect 269448 306972 269672 307000
rect 269448 306960 269454 306972
rect 269666 306960 269672 306972
rect 269724 306960 269730 307012
rect 325878 306960 325884 307012
rect 325936 307000 325942 307012
rect 326154 307000 326160 307012
rect 325936 306972 326160 307000
rect 325936 306960 325942 306972
rect 326154 306960 326160 306972
rect 326212 306960 326218 307012
rect 337102 306960 337108 307012
rect 337160 306960 337166 307012
rect 246022 306932 246028 306944
rect 234586 306904 246028 306932
rect 246022 306892 246028 306904
rect 246080 306892 246086 306944
rect 251450 306756 251456 306808
rect 251508 306796 251514 306808
rect 251560 306796 251588 306960
rect 261386 306824 261392 306876
rect 261444 306824 261450 306876
rect 283190 306824 283196 306876
rect 283248 306864 283254 306876
rect 283650 306864 283656 306876
rect 283248 306836 283656 306864
rect 283248 306824 283254 306836
rect 283650 306824 283656 306836
rect 283708 306824 283714 306876
rect 294046 306824 294052 306876
rect 294104 306824 294110 306876
rect 251508 306768 251588 306796
rect 251508 306756 251514 306768
rect 261404 306672 261432 306824
rect 263870 306688 263876 306740
rect 263928 306728 263934 306740
rect 264146 306728 264152 306740
rect 263928 306700 264152 306728
rect 263928 306688 263934 306700
rect 264146 306688 264152 306700
rect 264204 306688 264210 306740
rect 294064 306672 294092 306824
rect 337120 306796 337148 306960
rect 337194 306796 337200 306808
rect 337120 306768 337200 306796
rect 337194 306756 337200 306768
rect 337252 306756 337258 306808
rect 332686 306688 332692 306740
rect 332744 306728 332750 306740
rect 333054 306728 333060 306740
rect 332744 306700 333060 306728
rect 332744 306688 332750 306700
rect 333054 306688 333060 306700
rect 333112 306688 333118 306740
rect 261386 306620 261392 306672
rect 261444 306620 261450 306672
rect 294046 306620 294052 306672
rect 294104 306620 294110 306672
rect 263870 306552 263876 306604
rect 263928 306592 263934 306604
rect 264054 306592 264060 306604
rect 263928 306564 264060 306592
rect 263928 306552 263934 306564
rect 264054 306552 264060 306564
rect 264112 306552 264118 306604
rect 300854 306552 300860 306604
rect 300912 306592 300918 306604
rect 301314 306592 301320 306604
rect 300912 306564 301320 306592
rect 300912 306552 300918 306564
rect 301314 306552 301320 306564
rect 301372 306552 301378 306604
rect 252738 306484 252744 306536
rect 252796 306524 252802 306536
rect 253658 306524 253664 306536
rect 252796 306496 253664 306524
rect 252796 306484 252802 306496
rect 253658 306484 253664 306496
rect 253716 306484 253722 306536
rect 263594 306484 263600 306536
rect 263652 306524 263658 306536
rect 264606 306524 264612 306536
rect 263652 306496 264612 306524
rect 263652 306484 263658 306496
rect 264606 306484 264612 306496
rect 264664 306484 264670 306536
rect 282730 306484 282736 306536
rect 282788 306524 282794 306536
rect 289078 306524 289084 306536
rect 282788 306496 289084 306524
rect 282788 306484 282794 306496
rect 289078 306484 289084 306496
rect 289136 306484 289142 306536
rect 309134 306484 309140 306536
rect 309192 306524 309198 306536
rect 309594 306524 309600 306536
rect 309192 306496 309600 306524
rect 309192 306484 309198 306496
rect 309594 306484 309600 306496
rect 309652 306484 309658 306536
rect 329926 306484 329932 306536
rect 329984 306524 329990 306536
rect 330570 306524 330576 306536
rect 329984 306496 330576 306524
rect 329984 306484 329990 306496
rect 330570 306484 330576 306496
rect 330628 306484 330634 306536
rect 248598 306416 248604 306468
rect 248656 306456 248662 306468
rect 249518 306456 249524 306468
rect 248656 306428 249524 306456
rect 248656 306416 248662 306428
rect 249518 306416 249524 306428
rect 249576 306416 249582 306468
rect 252646 306416 252652 306468
rect 252704 306456 252710 306468
rect 253290 306456 253296 306468
rect 252704 306428 253296 306456
rect 252704 306416 252710 306428
rect 253290 306416 253296 306428
rect 253348 306416 253354 306468
rect 255590 306416 255596 306468
rect 255648 306456 255654 306468
rect 255866 306456 255872 306468
rect 255648 306428 255872 306456
rect 255648 306416 255654 306428
rect 255866 306416 255872 306428
rect 255924 306416 255930 306468
rect 258166 306416 258172 306468
rect 258224 306456 258230 306468
rect 258718 306456 258724 306468
rect 258224 306428 258724 306456
rect 258224 306416 258230 306428
rect 258718 306416 258724 306428
rect 258776 306416 258782 306468
rect 262214 306416 262220 306468
rect 262272 306456 262278 306468
rect 262858 306456 262864 306468
rect 262272 306428 262864 306456
rect 262272 306416 262278 306428
rect 262858 306416 262864 306428
rect 262916 306416 262922 306468
rect 263778 306416 263784 306468
rect 263836 306456 263842 306468
rect 264790 306456 264796 306468
rect 263836 306428 264796 306456
rect 263836 306416 263842 306428
rect 264790 306416 264796 306428
rect 264848 306416 264854 306468
rect 264974 306416 264980 306468
rect 265032 306456 265038 306468
rect 265434 306456 265440 306468
rect 265032 306428 265440 306456
rect 265032 306416 265038 306428
rect 265434 306416 265440 306428
rect 265492 306416 265498 306468
rect 266630 306416 266636 306468
rect 266688 306456 266694 306468
rect 266906 306456 266912 306468
rect 266688 306428 266912 306456
rect 266688 306416 266694 306428
rect 266906 306416 266912 306428
rect 266964 306416 266970 306468
rect 269758 306456 269764 306468
rect 269316 306428 269764 306456
rect 269316 306400 269344 306428
rect 269758 306416 269764 306428
rect 269816 306416 269822 306468
rect 271598 306416 271604 306468
rect 271656 306456 271662 306468
rect 272058 306456 272064 306468
rect 271656 306428 272064 306456
rect 271656 306416 271662 306428
rect 272058 306416 272064 306428
rect 272116 306416 272122 306468
rect 272150 306416 272156 306468
rect 272208 306456 272214 306468
rect 272794 306456 272800 306468
rect 272208 306428 272800 306456
rect 272208 306416 272214 306428
rect 272794 306416 272800 306428
rect 272852 306416 272858 306468
rect 273254 306416 273260 306468
rect 273312 306456 273318 306468
rect 273622 306456 273628 306468
rect 273312 306428 273628 306456
rect 273312 306416 273318 306428
rect 273622 306416 273628 306428
rect 273680 306416 273686 306468
rect 276198 306416 276204 306468
rect 276256 306456 276262 306468
rect 276474 306456 276480 306468
rect 276256 306428 276480 306456
rect 276256 306416 276262 306428
rect 276474 306416 276480 306428
rect 276532 306416 276538 306468
rect 277486 306416 277492 306468
rect 277544 306456 277550 306468
rect 278406 306456 278412 306468
rect 277544 306428 278412 306456
rect 277544 306416 277550 306428
rect 278406 306416 278412 306428
rect 278464 306416 278470 306468
rect 280522 306416 280528 306468
rect 280580 306456 280586 306468
rect 281442 306456 281448 306468
rect 280580 306428 281448 306456
rect 280580 306416 280586 306428
rect 281442 306416 281448 306428
rect 281500 306416 281506 306468
rect 281718 306416 281724 306468
rect 281776 306456 281782 306468
rect 282178 306456 282184 306468
rect 281776 306428 282184 306456
rect 281776 306416 281782 306428
rect 282178 306416 282184 306428
rect 282236 306416 282242 306468
rect 287422 306456 287428 306468
rect 282840 306428 287428 306456
rect 233326 306348 233332 306400
rect 233384 306388 233390 306400
rect 234154 306388 234160 306400
rect 233384 306360 234160 306388
rect 233384 306348 233390 306360
rect 234154 306348 234160 306360
rect 234212 306348 234218 306400
rect 241698 306348 241704 306400
rect 241756 306388 241762 306400
rect 242618 306388 242624 306400
rect 241756 306360 242624 306388
rect 241756 306348 241762 306360
rect 242618 306348 242624 306360
rect 242676 306348 242682 306400
rect 247126 306348 247132 306400
rect 247184 306388 247190 306400
rect 247954 306388 247960 306400
rect 247184 306360 247960 306388
rect 247184 306348 247190 306360
rect 247954 306348 247960 306360
rect 248012 306348 248018 306400
rect 248690 306348 248696 306400
rect 248748 306388 248754 306400
rect 249334 306388 249340 306400
rect 248748 306360 249340 306388
rect 248748 306348 248754 306360
rect 249334 306348 249340 306360
rect 249392 306348 249398 306400
rect 251266 306348 251272 306400
rect 251324 306388 251330 306400
rect 252370 306388 252376 306400
rect 251324 306360 252376 306388
rect 251324 306348 251330 306360
rect 252370 306348 252376 306360
rect 252428 306348 252434 306400
rect 252554 306348 252560 306400
rect 252612 306388 252618 306400
rect 253198 306388 253204 306400
rect 252612 306360 253204 306388
rect 252612 306348 252618 306360
rect 253198 306348 253204 306360
rect 253256 306348 253262 306400
rect 256694 306348 256700 306400
rect 256752 306388 256758 306400
rect 257338 306388 257344 306400
rect 256752 306360 257344 306388
rect 256752 306348 256758 306360
rect 257338 306348 257344 306360
rect 257396 306348 257402 306400
rect 258350 306348 258356 306400
rect 258408 306388 258414 306400
rect 258902 306388 258908 306400
rect 258408 306360 258908 306388
rect 258408 306348 258414 306360
rect 258902 306348 258908 306360
rect 258960 306348 258966 306400
rect 259546 306348 259552 306400
rect 259604 306388 259610 306400
rect 259822 306388 259828 306400
rect 259604 306360 259828 306388
rect 259604 306348 259610 306360
rect 259822 306348 259828 306360
rect 259880 306348 259886 306400
rect 259914 306348 259920 306400
rect 259972 306388 259978 306400
rect 260558 306388 260564 306400
rect 259972 306360 260564 306388
rect 259972 306348 259978 306360
rect 260558 306348 260564 306360
rect 260616 306348 260622 306400
rect 262398 306348 262404 306400
rect 262456 306388 262462 306400
rect 263042 306388 263048 306400
rect 262456 306360 263048 306388
rect 262456 306348 262462 306360
rect 263042 306348 263048 306360
rect 263100 306348 263106 306400
rect 263686 306348 263692 306400
rect 263744 306388 263750 306400
rect 264146 306388 264152 306400
rect 263744 306360 264152 306388
rect 263744 306348 263750 306360
rect 264146 306348 264152 306360
rect 264204 306348 264210 306400
rect 269298 306348 269304 306400
rect 269356 306348 269362 306400
rect 270862 306348 270868 306400
rect 270920 306388 270926 306400
rect 271322 306388 271328 306400
rect 270920 306360 271328 306388
rect 270920 306348 270926 306360
rect 271322 306348 271328 306360
rect 271380 306348 271386 306400
rect 272334 306348 272340 306400
rect 272392 306388 272398 306400
rect 273070 306388 273076 306400
rect 272392 306360 273076 306388
rect 272392 306348 272398 306360
rect 273070 306348 273076 306360
rect 273128 306348 273134 306400
rect 273530 306348 273536 306400
rect 273588 306388 273594 306400
rect 273806 306388 273812 306400
rect 273588 306360 273812 306388
rect 273588 306348 273594 306360
rect 273806 306348 273812 306360
rect 273864 306348 273870 306400
rect 275002 306348 275008 306400
rect 275060 306388 275066 306400
rect 275462 306388 275468 306400
rect 275060 306360 275468 306388
rect 275060 306348 275066 306360
rect 275462 306348 275468 306360
rect 275520 306348 275526 306400
rect 276014 306348 276020 306400
rect 276072 306388 276078 306400
rect 277210 306388 277216 306400
rect 276072 306360 277216 306388
rect 276072 306348 276078 306360
rect 277210 306348 277216 306360
rect 277268 306348 277274 306400
rect 277670 306348 277676 306400
rect 277728 306388 277734 306400
rect 278038 306388 278044 306400
rect 277728 306360 278044 306388
rect 277728 306348 277734 306360
rect 278038 306348 278044 306360
rect 278096 306348 278102 306400
rect 278866 306348 278872 306400
rect 278924 306388 278930 306400
rect 279510 306388 279516 306400
rect 278924 306360 279516 306388
rect 278924 306348 278930 306360
rect 279510 306348 279516 306360
rect 279568 306348 279574 306400
rect 280430 306348 280436 306400
rect 280488 306388 280494 306400
rect 281258 306388 281264 306400
rect 280488 306360 281264 306388
rect 280488 306348 280494 306360
rect 281258 306348 281264 306360
rect 281316 306348 281322 306400
rect 3326 306280 3332 306332
rect 3384 306320 3390 306332
rect 94498 306320 94504 306332
rect 3384 306292 94504 306320
rect 3384 306280 3390 306292
rect 94498 306280 94504 306292
rect 94556 306280 94562 306332
rect 218974 306280 218980 306332
rect 219032 306320 219038 306332
rect 282840 306320 282868 306428
rect 287422 306416 287428 306428
rect 287480 306416 287486 306468
rect 307846 306416 307852 306468
rect 307904 306456 307910 306468
rect 308490 306456 308496 306468
rect 307904 306428 308496 306456
rect 307904 306416 307910 306428
rect 308490 306416 308496 306428
rect 308548 306416 308554 306468
rect 309318 306416 309324 306468
rect 309376 306456 309382 306468
rect 309778 306456 309784 306468
rect 309376 306428 309784 306456
rect 309376 306416 309382 306428
rect 309778 306416 309784 306428
rect 309836 306416 309842 306468
rect 310514 306416 310520 306468
rect 310572 306456 310578 306468
rect 310882 306456 310888 306468
rect 310572 306428 310888 306456
rect 310572 306416 310578 306428
rect 310882 306416 310888 306428
rect 310940 306416 310946 306468
rect 322934 306416 322940 306468
rect 322992 306416 322998 306468
rect 327166 306416 327172 306468
rect 327224 306456 327230 306468
rect 327442 306456 327448 306468
rect 327224 306428 327448 306456
rect 327224 306416 327230 306428
rect 327442 306416 327448 306428
rect 327500 306416 327506 306468
rect 330110 306416 330116 306468
rect 330168 306456 330174 306468
rect 330386 306456 330392 306468
rect 330168 306428 330392 306456
rect 330168 306416 330174 306428
rect 330386 306416 330392 306428
rect 330444 306416 330450 306468
rect 333514 306456 333520 306468
rect 332796 306428 333520 306456
rect 291378 306348 291384 306400
rect 291436 306388 291442 306400
rect 291746 306388 291752 306400
rect 291436 306360 291752 306388
rect 291436 306348 291442 306360
rect 291746 306348 291752 306360
rect 291804 306348 291810 306400
rect 295334 306348 295340 306400
rect 295392 306388 295398 306400
rect 296346 306388 296352 306400
rect 295392 306360 296352 306388
rect 295392 306348 295398 306360
rect 296346 306348 296352 306360
rect 296404 306348 296410 306400
rect 296714 306348 296720 306400
rect 296772 306388 296778 306400
rect 297174 306388 297180 306400
rect 296772 306360 297180 306388
rect 296772 306348 296778 306360
rect 297174 306348 297180 306360
rect 297232 306348 297238 306400
rect 301130 306348 301136 306400
rect 301188 306388 301194 306400
rect 301314 306388 301320 306400
rect 301188 306360 301320 306388
rect 301188 306348 301194 306360
rect 301314 306348 301320 306360
rect 301372 306348 301378 306400
rect 303982 306348 303988 306400
rect 304040 306388 304046 306400
rect 304810 306388 304816 306400
rect 304040 306360 304816 306388
rect 304040 306348 304046 306360
rect 304810 306348 304816 306360
rect 304868 306348 304874 306400
rect 304994 306348 305000 306400
rect 305052 306388 305058 306400
rect 305546 306388 305552 306400
rect 305052 306360 305552 306388
rect 305052 306348 305058 306360
rect 305546 306348 305552 306360
rect 305604 306348 305610 306400
rect 321830 306348 321836 306400
rect 321888 306388 321894 306400
rect 322566 306388 322572 306400
rect 321888 306360 322572 306388
rect 321888 306348 321894 306360
rect 322566 306348 322572 306360
rect 322624 306348 322630 306400
rect 219032 306292 282868 306320
rect 219032 306280 219038 306292
rect 286042 306280 286048 306332
rect 286100 306320 286106 306332
rect 286778 306320 286784 306332
rect 286100 306292 286784 306320
rect 286100 306280 286106 306292
rect 286778 306280 286784 306292
rect 286836 306280 286842 306332
rect 289906 306280 289912 306332
rect 289964 306320 289970 306332
rect 290366 306320 290372 306332
rect 289964 306292 290372 306320
rect 289964 306280 289970 306292
rect 290366 306280 290372 306292
rect 290424 306280 290430 306332
rect 291470 306280 291476 306332
rect 291528 306320 291534 306332
rect 292390 306320 292396 306332
rect 291528 306292 292396 306320
rect 291528 306280 291534 306292
rect 292390 306280 292396 306292
rect 292448 306280 292454 306332
rect 292850 306280 292856 306332
rect 292908 306320 292914 306332
rect 293310 306320 293316 306332
rect 292908 306292 293316 306320
rect 292908 306280 292914 306292
rect 293310 306280 293316 306292
rect 293368 306280 293374 306332
rect 293954 306280 293960 306332
rect 294012 306320 294018 306332
rect 294230 306320 294236 306332
rect 294012 306292 294236 306320
rect 294012 306280 294018 306292
rect 294230 306280 294236 306292
rect 294288 306280 294294 306332
rect 295518 306280 295524 306332
rect 295576 306320 295582 306332
rect 296162 306320 296168 306332
rect 295576 306292 296168 306320
rect 295576 306280 295582 306292
rect 296162 306280 296168 306292
rect 296220 306280 296226 306332
rect 299474 306280 299480 306332
rect 299532 306320 299538 306332
rect 299750 306320 299756 306332
rect 299532 306292 299756 306320
rect 299532 306280 299538 306292
rect 299750 306280 299756 306292
rect 299808 306280 299814 306332
rect 303890 306280 303896 306332
rect 303948 306320 303954 306332
rect 304258 306320 304264 306332
rect 303948 306292 304264 306320
rect 303948 306280 303954 306292
rect 304258 306280 304264 306292
rect 304316 306280 304322 306332
rect 305086 306280 305092 306332
rect 305144 306320 305150 306332
rect 305730 306320 305736 306332
rect 305144 306292 305736 306320
rect 305144 306280 305150 306292
rect 305730 306280 305736 306292
rect 305788 306280 305794 306332
rect 306374 306280 306380 306332
rect 306432 306320 306438 306332
rect 307110 306320 307116 306332
rect 306432 306292 307116 306320
rect 306432 306280 306438 306292
rect 307110 306280 307116 306292
rect 307168 306280 307174 306332
rect 321646 306280 321652 306332
rect 321704 306320 321710 306332
rect 322106 306320 322112 306332
rect 321704 306292 322112 306320
rect 321704 306280 321710 306292
rect 322106 306280 322112 306292
rect 322164 306280 322170 306332
rect 218882 306212 218888 306264
rect 218940 306252 218946 306264
rect 282730 306252 282736 306264
rect 218940 306224 282736 306252
rect 218940 306212 218946 306224
rect 282730 306212 282736 306224
rect 282788 306212 282794 306264
rect 283006 306212 283012 306264
rect 283064 306252 283070 306264
rect 283926 306252 283932 306264
rect 283064 306224 283932 306252
rect 283064 306212 283070 306224
rect 283926 306212 283932 306224
rect 283984 306212 283990 306264
rect 288894 306212 288900 306264
rect 288952 306252 288958 306264
rect 289446 306252 289452 306264
rect 288952 306224 289452 306252
rect 288952 306212 288958 306224
rect 289446 306212 289452 306224
rect 289504 306212 289510 306264
rect 290182 306212 290188 306264
rect 290240 306252 290246 306264
rect 290826 306252 290832 306264
rect 290240 306224 290832 306252
rect 290240 306212 290246 306224
rect 290826 306212 290832 306224
rect 290884 306212 290890 306264
rect 291562 306212 291568 306264
rect 291620 306252 291626 306264
rect 292114 306252 292120 306264
rect 291620 306224 292120 306252
rect 291620 306212 291626 306224
rect 292114 306212 292120 306224
rect 292172 306212 292178 306264
rect 296714 306212 296720 306264
rect 296772 306252 296778 306264
rect 297082 306252 297088 306264
rect 296772 306224 297088 306252
rect 296772 306212 296778 306224
rect 297082 306212 297088 306224
rect 297140 306212 297146 306264
rect 302510 306212 302516 306264
rect 302568 306252 302574 306264
rect 303062 306252 303068 306264
rect 302568 306224 303068 306252
rect 302568 306212 302574 306224
rect 303062 306212 303068 306224
rect 303120 306212 303126 306264
rect 303706 306212 303712 306264
rect 303764 306252 303770 306264
rect 304166 306252 304172 306264
rect 303764 306224 304172 306252
rect 303764 306212 303770 306224
rect 304166 306212 304172 306224
rect 304224 306212 304230 306264
rect 305270 306212 305276 306264
rect 305328 306252 305334 306264
rect 305914 306252 305920 306264
rect 305328 306224 305920 306252
rect 305328 306212 305334 306224
rect 305914 306212 305920 306224
rect 305972 306212 305978 306264
rect 309502 306212 309508 306264
rect 309560 306252 309566 306264
rect 310146 306252 310152 306264
rect 309560 306224 310152 306252
rect 309560 306212 309566 306224
rect 310146 306212 310152 306224
rect 310204 306212 310210 306264
rect 310698 306212 310704 306264
rect 310756 306252 310762 306264
rect 310974 306252 310980 306264
rect 310756 306224 310980 306252
rect 310756 306212 310762 306224
rect 310974 306212 310980 306224
rect 311032 306212 311038 306264
rect 321554 306212 321560 306264
rect 321612 306252 321618 306264
rect 322750 306252 322756 306264
rect 321612 306224 322756 306252
rect 321612 306212 321618 306224
rect 322750 306212 322756 306224
rect 322808 306212 322814 306264
rect 169938 306144 169944 306196
rect 169996 306184 170002 306196
rect 238386 306184 238392 306196
rect 169996 306156 238392 306184
rect 169996 306144 170002 306156
rect 238386 306144 238392 306156
rect 238444 306144 238450 306196
rect 239030 306144 239036 306196
rect 239088 306184 239094 306196
rect 239490 306184 239496 306196
rect 239088 306156 239496 306184
rect 239088 306144 239094 306156
rect 239490 306144 239496 306156
rect 239548 306144 239554 306196
rect 242986 306144 242992 306196
rect 243044 306184 243050 306196
rect 244090 306184 244096 306196
rect 243044 306156 244096 306184
rect 243044 306144 243050 306156
rect 244090 306144 244096 306156
rect 244148 306144 244154 306196
rect 244550 306144 244556 306196
rect 244608 306184 244614 306196
rect 245102 306184 245108 306196
rect 244608 306156 245108 306184
rect 244608 306144 244614 306156
rect 245102 306144 245108 306156
rect 245160 306144 245166 306196
rect 250070 306144 250076 306196
rect 250128 306184 250134 306196
rect 250622 306184 250628 306196
rect 250128 306156 250628 306184
rect 250128 306144 250134 306156
rect 250622 306144 250628 306156
rect 250680 306144 250686 306196
rect 251542 306144 251548 306196
rect 251600 306184 251606 306196
rect 252186 306184 252192 306196
rect 251600 306156 252192 306184
rect 251600 306144 251606 306156
rect 252186 306144 252192 306156
rect 252244 306144 252250 306196
rect 252830 306144 252836 306196
rect 252888 306184 252894 306196
rect 253842 306184 253848 306196
rect 252888 306156 253848 306184
rect 252888 306144 252894 306156
rect 253842 306144 253848 306156
rect 253900 306144 253906 306196
rect 254026 306144 254032 306196
rect 254084 306184 254090 306196
rect 255038 306184 255044 306196
rect 254084 306156 255044 306184
rect 254084 306144 254090 306156
rect 255038 306144 255044 306156
rect 255096 306144 255102 306196
rect 255682 306144 255688 306196
rect 255740 306184 255746 306196
rect 256418 306184 256424 306196
rect 255740 306156 256424 306184
rect 255740 306144 255746 306156
rect 256418 306144 256424 306156
rect 256476 306144 256482 306196
rect 256970 306144 256976 306196
rect 257028 306184 257034 306196
rect 257706 306184 257712 306196
rect 257028 306156 257712 306184
rect 257028 306144 257034 306156
rect 257706 306144 257712 306156
rect 257764 306144 257770 306196
rect 258258 306144 258264 306196
rect 258316 306184 258322 306196
rect 258626 306184 258632 306196
rect 258316 306156 258632 306184
rect 258316 306144 258322 306156
rect 258626 306144 258632 306156
rect 258684 306144 258690 306196
rect 259454 306144 259460 306196
rect 259512 306184 259518 306196
rect 259822 306184 259828 306196
rect 259512 306156 259828 306184
rect 259512 306144 259518 306156
rect 259822 306144 259828 306156
rect 259880 306144 259886 306196
rect 261294 306144 261300 306196
rect 261352 306184 261358 306196
rect 261938 306184 261944 306196
rect 261352 306156 261944 306184
rect 261352 306144 261358 306156
rect 261938 306144 261944 306156
rect 261996 306144 262002 306196
rect 263686 306144 263692 306196
rect 263744 306184 263750 306196
rect 264238 306184 264244 306196
rect 263744 306156 264244 306184
rect 263744 306144 263750 306156
rect 264238 306144 264244 306156
rect 264296 306144 264302 306196
rect 265066 306144 265072 306196
rect 265124 306184 265130 306196
rect 265710 306184 265716 306196
rect 265124 306156 265716 306184
rect 265124 306144 265130 306156
rect 265710 306144 265716 306156
rect 265768 306144 265774 306196
rect 266722 306144 266728 306196
rect 266780 306184 266786 306196
rect 267090 306184 267096 306196
rect 266780 306156 267096 306184
rect 266780 306144 266786 306156
rect 267090 306144 267096 306156
rect 267148 306144 267154 306196
rect 269482 306144 269488 306196
rect 269540 306184 269546 306196
rect 270126 306184 270132 306196
rect 269540 306156 270132 306184
rect 269540 306144 269546 306156
rect 270126 306144 270132 306156
rect 270184 306144 270190 306196
rect 271966 306144 271972 306196
rect 272024 306184 272030 306196
rect 272978 306184 272984 306196
rect 272024 306156 272984 306184
rect 272024 306144 272030 306156
rect 272978 306144 272984 306156
rect 273036 306144 273042 306196
rect 273806 306144 273812 306196
rect 273864 306184 273870 306196
rect 274542 306184 274548 306196
rect 273864 306156 274548 306184
rect 273864 306144 273870 306156
rect 274542 306144 274548 306156
rect 274600 306144 274606 306196
rect 274634 306144 274640 306196
rect 274692 306184 274698 306196
rect 275094 306184 275100 306196
rect 274692 306156 275100 306184
rect 274692 306144 274698 306156
rect 275094 306144 275100 306156
rect 275152 306144 275158 306196
rect 278038 306144 278044 306196
rect 278096 306184 278102 306196
rect 278314 306184 278320 306196
rect 278096 306156 278320 306184
rect 278096 306144 278102 306156
rect 278314 306144 278320 306156
rect 278372 306144 278378 306196
rect 280246 306144 280252 306196
rect 280304 306184 280310 306196
rect 280706 306184 280712 306196
rect 280304 306156 280712 306184
rect 280304 306144 280310 306156
rect 280706 306144 280712 306156
rect 280764 306144 280770 306196
rect 282086 306144 282092 306196
rect 282144 306184 282150 306196
rect 282546 306184 282552 306196
rect 282144 306156 282552 306184
rect 282144 306144 282150 306156
rect 282546 306144 282552 306156
rect 282604 306144 282610 306196
rect 288526 306184 288532 306196
rect 283116 306156 288532 306184
rect 216398 306076 216404 306128
rect 216456 306116 216462 306128
rect 283116 306116 283144 306156
rect 288526 306144 288532 306156
rect 288584 306144 288590 306196
rect 290274 306144 290280 306196
rect 290332 306184 290338 306196
rect 291010 306184 291016 306196
rect 290332 306156 291016 306184
rect 290332 306144 290338 306156
rect 291010 306144 291016 306156
rect 291068 306144 291074 306196
rect 293126 306144 293132 306196
rect 293184 306184 293190 306196
rect 293678 306184 293684 306196
rect 293184 306156 293684 306184
rect 293184 306144 293190 306156
rect 293678 306144 293684 306156
rect 293736 306144 293742 306196
rect 294230 306144 294236 306196
rect 294288 306184 294294 306196
rect 294874 306184 294880 306196
rect 294288 306156 294880 306184
rect 294288 306144 294294 306156
rect 294874 306144 294880 306156
rect 294932 306144 294938 306196
rect 298094 306144 298100 306196
rect 298152 306184 298158 306196
rect 299382 306184 299388 306196
rect 298152 306156 299388 306184
rect 298152 306144 298158 306156
rect 299382 306144 299388 306156
rect 299440 306144 299446 306196
rect 299566 306144 299572 306196
rect 299624 306184 299630 306196
rect 300210 306184 300216 306196
rect 299624 306156 300216 306184
rect 299624 306144 299630 306156
rect 300210 306144 300216 306156
rect 300268 306144 300274 306196
rect 302326 306144 302332 306196
rect 302384 306184 302390 306196
rect 303430 306184 303436 306196
rect 302384 306156 303436 306184
rect 302384 306144 302390 306156
rect 303430 306144 303436 306156
rect 303488 306144 303494 306196
rect 303614 306144 303620 306196
rect 303672 306184 303678 306196
rect 304626 306184 304632 306196
rect 303672 306156 304632 306184
rect 303672 306144 303678 306156
rect 304626 306144 304632 306156
rect 304684 306144 304690 306196
rect 305362 306144 305368 306196
rect 305420 306184 305426 306196
rect 306098 306184 306104 306196
rect 305420 306156 306104 306184
rect 305420 306144 305426 306156
rect 306098 306144 306104 306156
rect 306156 306144 306162 306196
rect 309410 306144 309416 306196
rect 309468 306184 309474 306196
rect 310330 306184 310336 306196
rect 309468 306156 310336 306184
rect 309468 306144 309474 306156
rect 310330 306144 310336 306156
rect 310388 306144 310394 306196
rect 321738 306144 321744 306196
rect 321796 306184 321802 306196
rect 322198 306184 322204 306196
rect 321796 306156 322204 306184
rect 321796 306144 321802 306156
rect 322198 306144 322204 306156
rect 322256 306144 322262 306196
rect 322952 306184 322980 306416
rect 332796 306400 332824 306428
rect 333514 306416 333520 306428
rect 333572 306416 333578 306468
rect 337010 306416 337016 306468
rect 337068 306456 337074 306468
rect 337286 306456 337292 306468
rect 337068 306428 337292 306456
rect 337068 306416 337074 306428
rect 337286 306416 337292 306428
rect 337344 306416 337350 306468
rect 349706 306416 349712 306468
rect 349764 306416 349770 306468
rect 332778 306348 332784 306400
rect 332836 306348 332842 306400
rect 336826 306348 336832 306400
rect 336884 306388 336890 306400
rect 337654 306388 337660 306400
rect 336884 306360 337660 306388
rect 336884 306348 336890 306360
rect 337654 306348 337660 306360
rect 337712 306348 337718 306400
rect 324498 306280 324504 306332
rect 324556 306280 324562 306332
rect 327074 306280 327080 306332
rect 327132 306320 327138 306332
rect 327718 306320 327724 306332
rect 327132 306292 327724 306320
rect 327132 306280 327138 306292
rect 327718 306280 327724 306292
rect 327776 306280 327782 306332
rect 328454 306280 328460 306332
rect 328512 306320 328518 306332
rect 329098 306320 329104 306332
rect 328512 306292 329104 306320
rect 328512 306280 328518 306292
rect 329098 306280 329104 306292
rect 329156 306280 329162 306332
rect 330018 306280 330024 306332
rect 330076 306320 330082 306332
rect 330846 306320 330852 306332
rect 330076 306292 330852 306320
rect 330076 306280 330082 306292
rect 330846 306280 330852 306292
rect 330904 306280 330910 306332
rect 333238 306280 333244 306332
rect 333296 306320 333302 306332
rect 333698 306320 333704 306332
rect 333296 306292 333704 306320
rect 333296 306280 333302 306292
rect 333698 306280 333704 306292
rect 333756 306280 333762 306332
rect 334342 306280 334348 306332
rect 334400 306320 334406 306332
rect 334618 306320 334624 306332
rect 334400 306292 334624 306320
rect 334400 306280 334406 306292
rect 334618 306280 334624 306292
rect 334676 306280 334682 306332
rect 336734 306280 336740 306332
rect 336792 306320 336798 306332
rect 337286 306320 337292 306332
rect 336792 306292 337292 306320
rect 336792 306280 336798 306292
rect 337286 306280 337292 306292
rect 337344 306280 337350 306332
rect 341150 306280 341156 306332
rect 341208 306320 341214 306332
rect 341702 306320 341708 306332
rect 341208 306292 341708 306320
rect 341208 306280 341214 306292
rect 341702 306280 341708 306292
rect 341760 306280 341766 306332
rect 343634 306280 343640 306332
rect 343692 306320 343698 306332
rect 344186 306320 344192 306332
rect 343692 306292 344192 306320
rect 343692 306280 343698 306292
rect 344186 306280 344192 306292
rect 344244 306280 344250 306332
rect 349724 306320 349752 306416
rect 366266 306320 366272 306332
rect 349724 306292 366272 306320
rect 366266 306280 366272 306292
rect 366324 306280 366330 306332
rect 323302 306212 323308 306264
rect 323360 306252 323366 306264
rect 323762 306252 323768 306264
rect 323360 306224 323768 306252
rect 323360 306212 323366 306224
rect 323762 306212 323768 306224
rect 323820 306212 323826 306264
rect 323394 306184 323400 306196
rect 322952 306156 323400 306184
rect 323394 306144 323400 306156
rect 323452 306144 323458 306196
rect 216456 306088 283144 306116
rect 216456 306076 216462 306088
rect 283190 306076 283196 306128
rect 283248 306116 283254 306128
rect 283742 306116 283748 306128
rect 283248 306088 283748 306116
rect 283248 306076 283254 306088
rect 283742 306076 283748 306088
rect 283800 306076 283806 306128
rect 292942 306076 292948 306128
rect 293000 306116 293006 306128
rect 293862 306116 293868 306128
rect 293000 306088 293868 306116
rect 293000 306076 293006 306088
rect 293862 306076 293868 306088
rect 293920 306076 293926 306128
rect 294138 306076 294144 306128
rect 294196 306116 294202 306128
rect 295242 306116 295248 306128
rect 294196 306088 295248 306116
rect 294196 306076 294202 306088
rect 295242 306076 295248 306088
rect 295300 306076 295306 306128
rect 299474 306076 299480 306128
rect 299532 306116 299538 306128
rect 300762 306116 300768 306128
rect 299532 306088 300768 306116
rect 299532 306076 299538 306088
rect 300762 306076 300768 306088
rect 300820 306076 300826 306128
rect 301222 306076 301228 306128
rect 301280 306116 301286 306128
rect 301958 306116 301964 306128
rect 301280 306088 301964 306116
rect 301280 306076 301286 306088
rect 301958 306076 301964 306088
rect 302016 306076 302022 306128
rect 304994 306076 305000 306128
rect 305052 306116 305058 306128
rect 306282 306116 306288 306128
rect 305052 306088 306288 306116
rect 305052 306076 305058 306088
rect 306282 306076 306288 306088
rect 306340 306076 306346 306128
rect 306558 306076 306564 306128
rect 306616 306116 306622 306128
rect 307662 306116 307668 306128
rect 306616 306088 307668 306116
rect 306616 306076 306622 306088
rect 307662 306076 307668 306088
rect 307720 306076 307726 306128
rect 310698 306076 310704 306128
rect 310756 306116 310762 306128
rect 311526 306116 311532 306128
rect 310756 306088 311532 306116
rect 310756 306076 310762 306088
rect 311526 306076 311532 306088
rect 311584 306076 311590 306128
rect 321646 306076 321652 306128
rect 321704 306116 321710 306128
rect 322382 306116 322388 306128
rect 321704 306088 322388 306116
rect 321704 306076 321710 306088
rect 322382 306076 322388 306088
rect 322440 306076 322446 306128
rect 323026 306076 323032 306128
rect 323084 306116 323090 306128
rect 323578 306116 323584 306128
rect 323084 306088 323584 306116
rect 323084 306076 323090 306088
rect 323578 306076 323584 306088
rect 323636 306076 323642 306128
rect 324516 306116 324544 306280
rect 325970 306212 325976 306264
rect 326028 306252 326034 306264
rect 326614 306252 326620 306264
rect 326028 306224 326620 306252
rect 326028 306212 326034 306224
rect 326614 306212 326620 306224
rect 326672 306212 326678 306264
rect 327534 306212 327540 306264
rect 327592 306252 327598 306264
rect 328086 306252 328092 306264
rect 327592 306224 328092 306252
rect 327592 306212 327598 306224
rect 328086 306212 328092 306224
rect 328144 306212 328150 306264
rect 329834 306212 329840 306264
rect 329892 306252 329898 306264
rect 330386 306252 330392 306264
rect 329892 306224 330392 306252
rect 329892 306212 329898 306224
rect 330386 306212 330392 306224
rect 330444 306212 330450 306264
rect 336918 306212 336924 306264
rect 336976 306252 336982 306264
rect 337746 306252 337752 306264
rect 336976 306224 337752 306252
rect 336976 306212 336982 306224
rect 337746 306212 337752 306224
rect 337804 306212 337810 306264
rect 340966 306212 340972 306264
rect 341024 306252 341030 306264
rect 341886 306252 341892 306264
rect 341024 306224 341892 306252
rect 341024 306212 341030 306224
rect 341886 306212 341892 306224
rect 341944 306212 341950 306264
rect 342346 306212 342352 306264
rect 342404 306252 342410 306264
rect 342898 306252 342904 306264
rect 342404 306224 342904 306252
rect 342404 306212 342410 306224
rect 342898 306212 342904 306224
rect 342956 306212 342962 306264
rect 349154 306212 349160 306264
rect 349212 306252 349218 306264
rect 350166 306252 350172 306264
rect 349212 306224 350172 306252
rect 349212 306212 349218 306224
rect 350166 306212 350172 306224
rect 350224 306212 350230 306264
rect 350350 306212 350356 306264
rect 350408 306252 350414 306264
rect 366358 306252 366364 306264
rect 350408 306224 366364 306252
rect 350408 306212 350414 306224
rect 366358 306212 366364 306224
rect 366416 306212 366422 306264
rect 325878 306144 325884 306196
rect 325936 306184 325942 306196
rect 326430 306184 326436 306196
rect 325936 306156 326436 306184
rect 325936 306144 325942 306156
rect 326430 306144 326436 306156
rect 326488 306144 326494 306196
rect 327258 306144 327264 306196
rect 327316 306184 327322 306196
rect 327902 306184 327908 306196
rect 327316 306156 327908 306184
rect 327316 306144 327322 306156
rect 327902 306144 327908 306156
rect 327960 306144 327966 306196
rect 331674 306144 331680 306196
rect 331732 306184 331738 306196
rect 332502 306184 332508 306196
rect 331732 306156 332508 306184
rect 331732 306144 331738 306156
rect 332502 306144 332508 306156
rect 332560 306144 332566 306196
rect 332962 306144 332968 306196
rect 333020 306184 333026 306196
rect 333330 306184 333336 306196
rect 333020 306156 333336 306184
rect 333020 306144 333026 306156
rect 333330 306144 333336 306156
rect 333388 306144 333394 306196
rect 335262 306144 335268 306196
rect 335320 306184 335326 306196
rect 335630 306184 335636 306196
rect 335320 306156 335636 306184
rect 335320 306144 335326 306156
rect 335630 306144 335636 306156
rect 335688 306144 335694 306196
rect 335814 306144 335820 306196
rect 335872 306184 335878 306196
rect 336366 306184 336372 306196
rect 335872 306156 336372 306184
rect 335872 306144 335878 306156
rect 336366 306144 336372 306156
rect 336424 306144 336430 306196
rect 336734 306144 336740 306196
rect 336792 306184 336798 306196
rect 337930 306184 337936 306196
rect 336792 306156 337936 306184
rect 336792 306144 336798 306156
rect 337930 306144 337936 306156
rect 337988 306144 337994 306196
rect 338114 306144 338120 306196
rect 338172 306184 338178 306196
rect 338172 306156 338252 306184
rect 338172 306144 338178 306156
rect 324424 306088 324544 306116
rect 214926 306008 214932 306060
rect 214984 306048 214990 306060
rect 214984 306020 273254 306048
rect 214984 306008 214990 306020
rect 172238 305940 172244 305992
rect 172296 305980 172302 305992
rect 244918 305980 244924 305992
rect 172296 305952 244924 305980
rect 172296 305940 172302 305952
rect 244918 305940 244924 305952
rect 244976 305940 244982 305992
rect 254302 305940 254308 305992
rect 254360 305980 254366 305992
rect 255222 305980 255228 305992
rect 254360 305952 255228 305980
rect 254360 305940 254366 305952
rect 255222 305940 255228 305952
rect 255280 305940 255286 305992
rect 255406 305940 255412 305992
rect 255464 305980 255470 305992
rect 256326 305980 256332 305992
rect 255464 305952 256332 305980
rect 255464 305940 255470 305952
rect 256326 305940 256332 305952
rect 256384 305940 256390 305992
rect 257154 305940 257160 305992
rect 257212 305980 257218 305992
rect 257890 305980 257896 305992
rect 257212 305952 257896 305980
rect 257212 305940 257218 305952
rect 257890 305940 257896 305952
rect 257948 305940 257954 305992
rect 258258 305940 258264 305992
rect 258316 305980 258322 305992
rect 259270 305980 259276 305992
rect 258316 305952 259276 305980
rect 258316 305940 258322 305952
rect 259270 305940 259276 305952
rect 259328 305940 259334 305992
rect 259638 305940 259644 305992
rect 259696 305980 259702 305992
rect 260374 305980 260380 305992
rect 259696 305952 260380 305980
rect 259696 305940 259702 305952
rect 260374 305940 260380 305952
rect 260432 305940 260438 305992
rect 261110 305940 261116 305992
rect 261168 305980 261174 305992
rect 261754 305980 261760 305992
rect 261168 305952 261760 305980
rect 261168 305940 261174 305952
rect 261754 305940 261760 305952
rect 261812 305940 261818 305992
rect 263962 305940 263968 305992
rect 264020 305980 264026 305992
rect 264422 305980 264428 305992
rect 264020 305952 264428 305980
rect 264020 305940 264026 305952
rect 264422 305940 264428 305952
rect 264480 305940 264486 305992
rect 265250 305940 265256 305992
rect 265308 305980 265314 305992
rect 265894 305980 265900 305992
rect 265308 305952 265900 305980
rect 265308 305940 265314 305952
rect 265894 305940 265900 305952
rect 265952 305940 265958 305992
rect 266354 305940 266360 305992
rect 266412 305980 266418 305992
rect 266814 305980 266820 305992
rect 266412 305952 266820 305980
rect 266412 305940 266418 305952
rect 266814 305940 266820 305952
rect 266872 305940 266878 305992
rect 269390 305940 269396 305992
rect 269448 305980 269454 305992
rect 270310 305980 270316 305992
rect 269448 305952 270316 305980
rect 269448 305940 269454 305952
rect 270310 305940 270316 305952
rect 270368 305940 270374 305992
rect 270954 305940 270960 305992
rect 271012 305980 271018 305992
rect 271506 305980 271512 305992
rect 271012 305952 271512 305980
rect 271012 305940 271018 305952
rect 271506 305940 271512 305952
rect 271564 305940 271570 305992
rect 273226 305980 273254 306020
rect 273438 306008 273444 306060
rect 273496 306048 273502 306060
rect 273990 306048 273996 306060
rect 273496 306020 273996 306048
rect 273496 306008 273502 306020
rect 273990 306008 273996 306020
rect 274048 306008 274054 306060
rect 274818 306008 274824 306060
rect 274876 306048 274882 306060
rect 275554 306048 275560 306060
rect 274876 306020 275560 306048
rect 274876 306008 274882 306020
rect 275554 306008 275560 306020
rect 275612 306008 275618 306060
rect 276382 306008 276388 306060
rect 276440 306048 276446 306060
rect 277026 306048 277032 306060
rect 276440 306020 277032 306048
rect 276440 306008 276446 306020
rect 277026 306008 277032 306020
rect 277084 306008 277090 306060
rect 277762 306008 277768 306060
rect 277820 306048 277826 306060
rect 278222 306048 278228 306060
rect 277820 306020 278228 306048
rect 277820 306008 277826 306020
rect 278222 306008 278228 306020
rect 278280 306008 278286 306060
rect 279142 306008 279148 306060
rect 279200 306048 279206 306060
rect 279694 306048 279700 306060
rect 279200 306020 279700 306048
rect 279200 306008 279206 306020
rect 279694 306008 279700 306020
rect 279752 306008 279758 306060
rect 281810 306008 281816 306060
rect 281868 306048 281874 306060
rect 282362 306048 282368 306060
rect 281868 306020 282368 306048
rect 281868 306008 281874 306020
rect 282362 306008 282368 306020
rect 282420 306008 282426 306060
rect 287974 306048 287980 306060
rect 283116 306020 287980 306048
rect 283116 305980 283144 306020
rect 287974 306008 287980 306020
rect 288032 306008 288038 306060
rect 292758 306008 292764 306060
rect 292816 306048 292822 306060
rect 293494 306048 293500 306060
rect 292816 306020 293500 306048
rect 292816 306008 292822 306020
rect 293494 306008 293500 306020
rect 293552 306008 293558 306060
rect 296806 306008 296812 306060
rect 296864 306048 296870 306060
rect 297726 306048 297732 306060
rect 296864 306020 297732 306048
rect 296864 306008 296870 306020
rect 297726 306008 297732 306020
rect 297784 306008 297790 306060
rect 300854 306008 300860 306060
rect 300912 306048 300918 306060
rect 301866 306048 301872 306060
rect 300912 306020 301872 306048
rect 300912 306008 300918 306020
rect 301866 306008 301872 306020
rect 301924 306008 301930 306060
rect 323210 306008 323216 306060
rect 323268 306048 323274 306060
rect 323946 306048 323952 306060
rect 323268 306020 323952 306048
rect 323268 306008 323274 306020
rect 323946 306008 323952 306020
rect 324004 306008 324010 306060
rect 324424 305992 324452 306088
rect 324590 306076 324596 306128
rect 324648 306116 324654 306128
rect 325418 306116 325424 306128
rect 324648 306088 325424 306116
rect 324648 306076 324654 306088
rect 325418 306076 325424 306088
rect 325476 306076 325482 306128
rect 327350 306076 327356 306128
rect 327408 306116 327414 306128
rect 328178 306116 328184 306128
rect 327408 306088 328184 306116
rect 327408 306076 327414 306088
rect 328178 306076 328184 306088
rect 328236 306076 328242 306128
rect 328822 306076 328828 306128
rect 328880 306116 328886 306128
rect 329466 306116 329472 306128
rect 328880 306088 329472 306116
rect 328880 306076 328886 306088
rect 329466 306076 329472 306088
rect 329524 306076 329530 306128
rect 331490 306076 331496 306128
rect 331548 306116 331554 306128
rect 331950 306116 331956 306128
rect 331548 306088 331956 306116
rect 331548 306076 331554 306088
rect 331950 306076 331956 306088
rect 332008 306076 332014 306128
rect 334434 306076 334440 306128
rect 334492 306116 334498 306128
rect 334986 306116 334992 306128
rect 334492 306088 334992 306116
rect 334492 306076 334498 306088
rect 334986 306076 334992 306088
rect 335044 306076 335050 306128
rect 335446 306076 335452 306128
rect 335504 306116 335510 306128
rect 336182 306116 336188 306128
rect 335504 306088 336188 306116
rect 335504 306076 335510 306088
rect 336182 306076 336188 306088
rect 336240 306076 336246 306128
rect 328914 306008 328920 306060
rect 328972 306048 328978 306060
rect 329282 306048 329288 306060
rect 328972 306020 329288 306048
rect 328972 306008 328978 306020
rect 329282 306008 329288 306020
rect 329340 306008 329346 306060
rect 331398 306008 331404 306060
rect 331456 306048 331462 306060
rect 332134 306048 332140 306060
rect 331456 306020 332140 306048
rect 331456 306008 331462 306020
rect 332134 306008 332140 306020
rect 332192 306008 332198 306060
rect 334158 306008 334164 306060
rect 334216 306048 334222 306060
rect 334802 306048 334808 306060
rect 334216 306020 334808 306048
rect 334216 306008 334222 306020
rect 334802 306008 334808 306020
rect 334860 306008 334866 306060
rect 338224 305992 338252 306156
rect 349982 306144 349988 306196
rect 350040 306184 350046 306196
rect 367554 306184 367560 306196
rect 350040 306156 367560 306184
rect 350040 306144 350046 306156
rect 367554 306144 367560 306156
rect 367612 306144 367618 306196
rect 348970 306076 348976 306128
rect 349028 306116 349034 306128
rect 365898 306116 365904 306128
rect 349028 306088 365904 306116
rect 349028 306076 349034 306088
rect 365898 306076 365904 306088
rect 365956 306076 365962 306128
rect 349338 306008 349344 306060
rect 349396 306048 349402 306060
rect 367738 306048 367744 306060
rect 349396 306020 367744 306048
rect 349396 306008 349402 306020
rect 367738 306008 367744 306020
rect 367796 306008 367802 306060
rect 273226 305952 283144 305980
rect 296898 305940 296904 305992
rect 296956 305980 296962 305992
rect 297542 305980 297548 305992
rect 296956 305952 297548 305980
rect 296956 305940 296962 305952
rect 297542 305940 297548 305952
rect 297600 305940 297606 305992
rect 324406 305940 324412 305992
rect 324464 305940 324470 305992
rect 324498 305940 324504 305992
rect 324556 305980 324562 305992
rect 325602 305980 325608 305992
rect 324556 305952 325608 305980
rect 324556 305940 324562 305952
rect 325602 305940 325608 305952
rect 325660 305940 325666 305992
rect 328546 305940 328552 305992
rect 328604 305980 328610 305992
rect 329006 305980 329012 305992
rect 328604 305952 329012 305980
rect 328604 305940 328610 305952
rect 329006 305940 329012 305952
rect 329064 305940 329070 305992
rect 329926 305940 329932 305992
rect 329984 305980 329990 305992
rect 331030 305980 331036 305992
rect 329984 305952 331036 305980
rect 329984 305940 329990 305952
rect 331030 305940 331036 305952
rect 331088 305940 331094 305992
rect 334250 305940 334256 305992
rect 334308 305980 334314 305992
rect 335170 305980 335176 305992
rect 334308 305952 335176 305980
rect 334308 305940 334314 305952
rect 335170 305940 335176 305952
rect 335228 305940 335234 305992
rect 338206 305940 338212 305992
rect 338264 305940 338270 305992
rect 348602 305940 348608 305992
rect 348660 305980 348666 305992
rect 367646 305980 367652 305992
rect 348660 305952 367652 305980
rect 348660 305940 348666 305952
rect 367646 305940 367652 305952
rect 367704 305940 367710 305992
rect 216306 305872 216312 305924
rect 216364 305912 216370 305924
rect 290642 305912 290648 305924
rect 216364 305884 290648 305912
rect 216364 305872 216370 305884
rect 290642 305872 290648 305884
rect 290700 305872 290706 305924
rect 324222 305872 324228 305924
rect 324280 305912 324286 305924
rect 324866 305912 324872 305924
rect 324280 305884 324872 305912
rect 324280 305872 324286 305884
rect 324866 305872 324872 305884
rect 324924 305872 324930 305924
rect 331766 305872 331772 305924
rect 331824 305912 331830 305924
rect 332318 305912 332324 305924
rect 331824 305884 332324 305912
rect 331824 305872 331830 305884
rect 332318 305872 332324 305884
rect 332376 305872 332382 305924
rect 344002 305872 344008 305924
rect 344060 305912 344066 305924
rect 367462 305912 367468 305924
rect 344060 305884 367468 305912
rect 344060 305872 344066 305884
rect 367462 305872 367468 305884
rect 367520 305872 367526 305924
rect 216582 305804 216588 305856
rect 216640 305844 216646 305856
rect 291194 305844 291200 305856
rect 216640 305816 291200 305844
rect 216640 305804 216646 305816
rect 291194 305804 291200 305816
rect 291252 305804 291258 305856
rect 328546 305804 328552 305856
rect 328604 305844 328610 305856
rect 329650 305844 329656 305856
rect 328604 305816 329656 305844
rect 328604 305804 328610 305816
rect 329650 305804 329656 305816
rect 329708 305804 329714 305856
rect 332778 305804 332784 305856
rect 332836 305844 332842 305856
rect 333882 305844 333888 305856
rect 332836 305816 333888 305844
rect 332836 305804 332842 305816
rect 333882 305804 333888 305816
rect 333940 305804 333946 305856
rect 344554 305804 344560 305856
rect 344612 305844 344618 305856
rect 367830 305844 367836 305856
rect 344612 305816 367836 305844
rect 344612 305804 344618 305816
rect 367830 305804 367836 305816
rect 367888 305804 367894 305856
rect 213822 305736 213828 305788
rect 213880 305776 213886 305788
rect 290090 305776 290096 305788
rect 213880 305748 290096 305776
rect 213880 305736 213886 305748
rect 290090 305736 290096 305748
rect 290148 305736 290154 305788
rect 342622 305736 342628 305788
rect 342680 305776 342686 305788
rect 368566 305776 368572 305788
rect 342680 305748 368572 305776
rect 342680 305736 342686 305748
rect 368566 305736 368572 305748
rect 368624 305736 368630 305788
rect 212074 305668 212080 305720
rect 212132 305708 212138 305720
rect 289630 305708 289636 305720
rect 212132 305680 289636 305708
rect 212132 305668 212138 305680
rect 289630 305668 289636 305680
rect 289688 305668 289694 305720
rect 343082 305668 343088 305720
rect 343140 305708 343146 305720
rect 368842 305708 368848 305720
rect 343140 305680 368848 305708
rect 343140 305668 343146 305680
rect 368842 305668 368848 305680
rect 368900 305668 368906 305720
rect 175918 305600 175924 305652
rect 175976 305640 175982 305652
rect 274634 305640 274640 305652
rect 175976 305612 274640 305640
rect 175976 305600 175982 305612
rect 274634 305600 274640 305612
rect 274692 305600 274698 305652
rect 274910 305600 274916 305652
rect 274968 305640 274974 305652
rect 275922 305640 275928 305652
rect 274968 305612 275928 305640
rect 274968 305600 274974 305612
rect 275922 305600 275928 305612
rect 275980 305600 275986 305652
rect 278958 305600 278964 305652
rect 279016 305640 279022 305652
rect 279418 305640 279424 305652
rect 279016 305612 279424 305640
rect 279016 305600 279022 305612
rect 279418 305600 279424 305612
rect 279476 305600 279482 305652
rect 281994 305600 282000 305652
rect 282052 305640 282058 305652
rect 282822 305640 282828 305652
rect 282052 305612 282828 305640
rect 282052 305600 282058 305612
rect 282822 305600 282828 305612
rect 282880 305600 282886 305652
rect 298186 305600 298192 305652
rect 298244 305640 298250 305652
rect 299014 305640 299020 305652
rect 298244 305612 299020 305640
rect 298244 305600 298250 305612
rect 299014 305600 299020 305612
rect 299072 305600 299078 305652
rect 342070 305600 342076 305652
rect 342128 305640 342134 305652
rect 368934 305640 368940 305652
rect 342128 305612 368940 305640
rect 342128 305600 342134 305612
rect 368934 305600 368940 305612
rect 368992 305600 368998 305652
rect 219066 305532 219072 305584
rect 219124 305572 219130 305584
rect 286410 305572 286416 305584
rect 219124 305544 286416 305572
rect 219124 305532 219130 305544
rect 286410 305532 286416 305544
rect 286468 305532 286474 305584
rect 350902 305532 350908 305584
rect 350960 305572 350966 305584
rect 366174 305572 366180 305584
rect 350960 305544 366180 305572
rect 350960 305532 350966 305544
rect 366174 305532 366180 305544
rect 366232 305532 366238 305584
rect 219158 305464 219164 305516
rect 219216 305504 219222 305516
rect 285306 305504 285312 305516
rect 219216 305476 285312 305504
rect 219216 305464 219222 305476
rect 285306 305464 285312 305476
rect 285364 305464 285370 305516
rect 350994 305464 351000 305516
rect 351052 305504 351058 305516
rect 366082 305504 366088 305516
rect 351052 305476 366088 305504
rect 351052 305464 351058 305476
rect 366082 305464 366088 305476
rect 366140 305464 366146 305516
rect 172606 305396 172612 305448
rect 172664 305436 172670 305448
rect 236270 305436 236276 305448
rect 172664 305408 236276 305436
rect 172664 305396 172670 305408
rect 236270 305396 236276 305408
rect 236328 305396 236334 305448
rect 238938 305396 238944 305448
rect 238996 305436 239002 305448
rect 239950 305436 239956 305448
rect 238996 305408 239956 305436
rect 238996 305396 239002 305408
rect 239950 305396 239956 305408
rect 240008 305396 240014 305448
rect 254210 305396 254216 305448
rect 254268 305436 254274 305448
rect 254578 305436 254584 305448
rect 254268 305408 254584 305436
rect 254268 305396 254274 305408
rect 254578 305396 254584 305408
rect 254636 305396 254642 305448
rect 256786 305396 256792 305448
rect 256844 305436 256850 305448
rect 257246 305436 257252 305448
rect 256844 305408 257252 305436
rect 256844 305396 256850 305408
rect 257246 305396 257252 305408
rect 257304 305396 257310 305448
rect 259454 305396 259460 305448
rect 259512 305436 259518 305448
rect 260006 305436 260012 305448
rect 259512 305408 260012 305436
rect 259512 305396 259518 305408
rect 260006 305396 260012 305408
rect 260064 305396 260070 305448
rect 260926 305396 260932 305448
rect 260984 305436 260990 305448
rect 261570 305436 261576 305448
rect 260984 305408 261576 305436
rect 260984 305396 260990 305408
rect 261570 305396 261576 305408
rect 261628 305396 261634 305448
rect 265342 305396 265348 305448
rect 265400 305436 265406 305448
rect 266170 305436 266176 305448
rect 265400 305408 266176 305436
rect 265400 305396 265406 305408
rect 266170 305396 266176 305408
rect 266228 305396 266234 305448
rect 266630 305396 266636 305448
rect 266688 305436 266694 305448
rect 267274 305436 267280 305448
rect 266688 305408 267280 305436
rect 266688 305396 266694 305408
rect 267274 305396 267280 305408
rect 267332 305396 267338 305448
rect 267826 305396 267832 305448
rect 267884 305436 267890 305448
rect 268286 305436 268292 305448
rect 267884 305408 268292 305436
rect 267884 305396 267890 305408
rect 268286 305396 268292 305408
rect 268344 305396 268350 305448
rect 273714 305396 273720 305448
rect 273772 305436 273778 305448
rect 274174 305436 274180 305448
rect 273772 305408 274180 305436
rect 273772 305396 273778 305408
rect 274174 305396 274180 305408
rect 274232 305396 274238 305448
rect 274634 305396 274640 305448
rect 274692 305436 274698 305448
rect 276842 305436 276848 305448
rect 274692 305408 276848 305436
rect 274692 305396 274698 305408
rect 276842 305396 276848 305408
rect 276900 305396 276906 305448
rect 278958 305396 278964 305448
rect 279016 305436 279022 305448
rect 280062 305436 280068 305448
rect 279016 305408 280068 305436
rect 279016 305396 279022 305408
rect 280062 305396 280068 305408
rect 280120 305396 280126 305448
rect 281718 305396 281724 305448
rect 281776 305436 281782 305448
rect 282638 305436 282644 305448
rect 281776 305408 282644 305436
rect 281776 305396 281782 305408
rect 282638 305396 282644 305408
rect 282696 305396 282702 305448
rect 351454 305396 351460 305448
rect 351512 305436 351518 305448
rect 361022 305436 361028 305448
rect 351512 305408 361028 305436
rect 351512 305396 351518 305408
rect 361022 305396 361028 305408
rect 361080 305396 361086 305448
rect 238662 305328 238668 305380
rect 238720 305368 238726 305380
rect 239766 305368 239772 305380
rect 238720 305340 239772 305368
rect 238720 305328 238726 305340
rect 239766 305328 239772 305340
rect 239824 305328 239830 305380
rect 267734 305328 267740 305380
rect 267792 305368 267798 305380
rect 268194 305368 268200 305380
rect 267792 305340 268200 305368
rect 267792 305328 267798 305340
rect 268194 305328 268200 305340
rect 268252 305328 268258 305380
rect 238386 305260 238392 305312
rect 238444 305300 238450 305312
rect 242250 305300 242256 305312
rect 238444 305272 242256 305300
rect 238444 305260 238450 305272
rect 242250 305260 242256 305272
rect 242308 305260 242314 305312
rect 256786 305260 256792 305312
rect 256844 305300 256850 305312
rect 257522 305300 257528 305312
rect 256844 305272 257528 305300
rect 256844 305260 256850 305272
rect 257522 305260 257528 305272
rect 257580 305260 257586 305312
rect 267826 305260 267832 305312
rect 267884 305300 267890 305312
rect 268838 305300 268844 305312
rect 267884 305272 268844 305300
rect 267884 305260 267890 305272
rect 268838 305260 268844 305272
rect 268896 305260 268902 305312
rect 97166 305192 97172 305244
rect 97224 305232 97230 305244
rect 97534 305232 97540 305244
rect 97224 305204 97540 305232
rect 97224 305192 97230 305204
rect 97534 305192 97540 305204
rect 97592 305192 97598 305244
rect 307938 305192 307944 305244
rect 307996 305232 308002 305244
rect 308766 305232 308772 305244
rect 307996 305204 308772 305232
rect 307996 305192 308002 305204
rect 308766 305192 308772 305204
rect 308824 305192 308830 305244
rect 97534 305056 97540 305108
rect 97592 305096 97598 305108
rect 97810 305096 97816 305108
rect 97592 305068 97816 305096
rect 97592 305056 97598 305068
rect 97810 305056 97816 305068
rect 97868 305056 97874 305108
rect 262490 304988 262496 305040
rect 262548 305028 262554 305040
rect 262858 305028 262864 305040
rect 262548 305000 262864 305028
rect 262548 304988 262554 305000
rect 262858 304988 262864 305000
rect 262916 304988 262922 305040
rect 172330 304920 172336 304972
rect 172388 304960 172394 304972
rect 244274 304960 244280 304972
rect 172388 304932 244280 304960
rect 172388 304920 172394 304932
rect 244274 304920 244280 304932
rect 244332 304920 244338 304972
rect 247218 304920 247224 304972
rect 247276 304960 247282 304972
rect 249702 304960 249708 304972
rect 247276 304932 249708 304960
rect 247276 304920 247282 304932
rect 249702 304920 249708 304932
rect 249760 304920 249766 304972
rect 262306 304920 262312 304972
rect 262364 304960 262370 304972
rect 262766 304960 262772 304972
rect 262364 304932 262772 304960
rect 262364 304920 262370 304932
rect 262766 304920 262772 304932
rect 262824 304920 262830 304972
rect 262490 304852 262496 304904
rect 262548 304892 262554 304904
rect 263502 304892 263508 304904
rect 262548 304864 263508 304892
rect 262548 304852 262554 304864
rect 263502 304852 263508 304864
rect 263560 304852 263566 304904
rect 325694 304852 325700 304904
rect 325752 304892 325758 304904
rect 326798 304892 326804 304904
rect 325752 304864 326804 304892
rect 325752 304852 325758 304864
rect 326798 304852 326804 304864
rect 326856 304852 326862 304904
rect 301406 304648 301412 304700
rect 301464 304688 301470 304700
rect 302142 304688 302148 304700
rect 301464 304660 302148 304688
rect 301464 304648 301470 304660
rect 302142 304648 302148 304660
rect 302200 304648 302206 304700
rect 169846 304444 169852 304496
rect 169904 304484 169910 304496
rect 237834 304484 237840 304496
rect 169904 304456 237840 304484
rect 169904 304444 169910 304456
rect 237834 304444 237840 304456
rect 237892 304444 237898 304496
rect 342438 304444 342444 304496
rect 342496 304484 342502 304496
rect 342714 304484 342720 304496
rect 342496 304456 342720 304484
rect 342496 304444 342502 304456
rect 342714 304444 342720 304456
rect 342772 304444 342778 304496
rect 171686 304376 171692 304428
rect 171744 304416 171750 304428
rect 244366 304416 244372 304428
rect 171744 304388 244372 304416
rect 171744 304376 171750 304388
rect 244366 304376 244372 304388
rect 244424 304376 244430 304428
rect 308122 304376 308128 304428
rect 308180 304416 308186 304428
rect 308950 304416 308956 304428
rect 308180 304388 308956 304416
rect 308180 304376 308186 304388
rect 308950 304376 308956 304388
rect 309008 304376 309014 304428
rect 170030 304308 170036 304360
rect 170088 304348 170094 304360
rect 247586 304348 247592 304360
rect 170088 304320 247592 304348
rect 170088 304308 170094 304320
rect 247586 304308 247592 304320
rect 247644 304308 247650 304360
rect 171870 304240 171876 304292
rect 171928 304280 171934 304292
rect 254854 304280 254860 304292
rect 171928 304252 254860 304280
rect 171928 304240 171934 304252
rect 254854 304240 254860 304252
rect 254912 304240 254918 304292
rect 271046 304240 271052 304292
rect 271104 304280 271110 304292
rect 271690 304280 271696 304292
rect 271104 304252 271696 304280
rect 271104 304240 271110 304252
rect 271690 304240 271696 304252
rect 271748 304240 271754 304292
rect 236086 304172 236092 304224
rect 236144 304212 236150 304224
rect 236270 304212 236276 304224
rect 236144 304184 236276 304212
rect 236144 304172 236150 304184
rect 236270 304172 236276 304184
rect 236328 304172 236334 304224
rect 255774 304104 255780 304156
rect 255832 304144 255838 304156
rect 256142 304144 256148 304156
rect 255832 304116 256148 304144
rect 255832 304104 255838 304116
rect 256142 304104 256148 304116
rect 256200 304104 256206 304156
rect 310606 304104 310612 304156
rect 310664 304144 310670 304156
rect 310882 304144 310888 304156
rect 310664 304116 310888 304144
rect 310664 304104 310670 304116
rect 310882 304104 310888 304116
rect 310940 304104 310946 304156
rect 337102 304104 337108 304156
rect 337160 304144 337166 304156
rect 337470 304144 337476 304156
rect 337160 304116 337476 304144
rect 337160 304104 337166 304116
rect 337470 304104 337476 304116
rect 337528 304104 337534 304156
rect 310606 303968 310612 304020
rect 310664 304008 310670 304020
rect 311434 304008 311440 304020
rect 310664 303980 311440 304008
rect 310664 303968 310670 303980
rect 311434 303968 311440 303980
rect 311492 303968 311498 304020
rect 302418 303696 302424 303748
rect 302476 303736 302482 303748
rect 302878 303736 302884 303748
rect 302476 303708 302884 303736
rect 302476 303696 302482 303708
rect 302878 303696 302884 303708
rect 302936 303696 302942 303748
rect 216122 303560 216128 303612
rect 216180 303600 216186 303612
rect 285950 303600 285956 303612
rect 216180 303572 285956 303600
rect 216180 303560 216186 303572
rect 285950 303560 285956 303572
rect 286008 303560 286014 303612
rect 349246 303560 349252 303612
rect 349304 303600 349310 303612
rect 371326 303600 371332 303612
rect 349304 303572 371332 303600
rect 349304 303560 349310 303572
rect 371326 303560 371332 303572
rect 371384 303560 371390 303612
rect 214742 303492 214748 303544
rect 214800 303532 214806 303544
rect 285490 303532 285496 303544
rect 214800 303504 285496 303532
rect 214800 303492 214806 303504
rect 285490 303492 285496 303504
rect 285548 303492 285554 303544
rect 349798 303492 349804 303544
rect 349856 303532 349862 303544
rect 371602 303532 371608 303544
rect 349856 303504 371608 303532
rect 349856 303492 349862 303504
rect 371602 303492 371608 303504
rect 371660 303492 371666 303544
rect 216490 303424 216496 303476
rect 216548 303464 216554 303476
rect 287146 303464 287152 303476
rect 216548 303436 287152 303464
rect 216548 303424 216554 303436
rect 287146 303424 287152 303436
rect 287204 303424 287210 303476
rect 348418 303424 348424 303476
rect 348476 303464 348482 303476
rect 370498 303464 370504 303476
rect 348476 303436 370504 303464
rect 348476 303424 348482 303436
rect 370498 303424 370504 303436
rect 370556 303424 370562 303476
rect 216214 303356 216220 303408
rect 216272 303396 216278 303408
rect 288158 303396 288164 303408
rect 216272 303368 288164 303396
rect 216272 303356 216278 303368
rect 288158 303356 288164 303368
rect 288216 303356 288222 303408
rect 347682 303356 347688 303408
rect 347740 303396 347746 303408
rect 369118 303396 369124 303408
rect 347740 303368 369124 303396
rect 347740 303356 347746 303368
rect 369118 303356 369124 303368
rect 369176 303356 369182 303408
rect 214834 303288 214840 303340
rect 214892 303328 214898 303340
rect 286594 303328 286600 303340
rect 214892 303300 286600 303328
rect 214892 303288 214898 303300
rect 286594 303288 286600 303300
rect 286652 303288 286658 303340
rect 346670 303288 346676 303340
rect 346728 303328 346734 303340
rect 369946 303328 369952 303340
rect 346728 303300 369952 303328
rect 346728 303288 346734 303300
rect 369946 303288 369952 303300
rect 370004 303288 370010 303340
rect 214650 303220 214656 303272
rect 214708 303260 214714 303272
rect 287606 303260 287612 303272
rect 214708 303232 287612 303260
rect 214708 303220 214714 303232
rect 287606 303220 287612 303232
rect 287664 303220 287670 303272
rect 349522 303220 349528 303272
rect 349580 303260 349586 303272
rect 372982 303260 372988 303272
rect 349580 303232 372988 303260
rect 349580 303220 349586 303232
rect 372982 303220 372988 303232
rect 373040 303220 373046 303272
rect 215018 303152 215024 303204
rect 215076 303192 215082 303204
rect 292298 303192 292304 303204
rect 215076 303164 292304 303192
rect 215076 303152 215082 303164
rect 292298 303152 292304 303164
rect 292356 303152 292362 303204
rect 347314 303152 347320 303204
rect 347372 303192 347378 303204
rect 370682 303192 370688 303204
rect 347372 303164 370688 303192
rect 347372 303152 347378 303164
rect 370682 303152 370688 303164
rect 370740 303152 370746 303204
rect 213454 303084 213460 303136
rect 213512 303124 213518 303136
rect 290458 303124 290464 303136
rect 213512 303096 290464 303124
rect 213512 303084 213518 303096
rect 290458 303084 290464 303096
rect 290516 303084 290522 303136
rect 347038 303084 347044 303136
rect 347096 303124 347102 303136
rect 370590 303124 370596 303136
rect 347096 303096 370596 303124
rect 347096 303084 347102 303096
rect 370590 303084 370596 303096
rect 370648 303084 370654 303136
rect 212442 303016 212448 303068
rect 212500 303056 212506 303068
rect 291838 303056 291844 303068
rect 212500 303028 291844 303056
rect 212500 303016 212506 303028
rect 291838 303016 291844 303028
rect 291896 303016 291902 303068
rect 346302 303016 346308 303068
rect 346360 303056 346366 303068
rect 370130 303056 370136 303068
rect 346360 303028 370136 303056
rect 346360 303016 346366 303028
rect 370130 303016 370136 303028
rect 370188 303016 370194 303068
rect 171962 302948 171968 303000
rect 172020 302988 172026 303000
rect 252002 302988 252008 303000
rect 172020 302960 252008 302988
rect 172020 302948 172026 302960
rect 252002 302948 252008 302960
rect 252060 302948 252066 303000
rect 345934 302948 345940 303000
rect 345992 302988 345998 303000
rect 370038 302988 370044 303000
rect 345992 302960 370044 302988
rect 345992 302948 345998 302960
rect 370038 302948 370044 302960
rect 370096 302948 370102 303000
rect 175274 302880 175280 302932
rect 175332 302920 175338 302932
rect 275370 302920 275376 302932
rect 175332 302892 275376 302920
rect 175332 302880 175338 302892
rect 275370 302880 275376 302892
rect 275428 302880 275434 302932
rect 345566 302880 345572 302932
rect 345624 302920 345630 302932
rect 370222 302920 370228 302932
rect 345624 302892 370228 302920
rect 345624 302880 345630 302892
rect 370222 302880 370228 302892
rect 370280 302880 370286 302932
rect 216030 302812 216036 302864
rect 216088 302852 216094 302864
rect 285674 302852 285680 302864
rect 216088 302824 285680 302852
rect 216088 302812 216094 302824
rect 285674 302812 285680 302824
rect 285732 302812 285738 302864
rect 348786 302812 348792 302864
rect 348844 302852 348850 302864
rect 369210 302852 369216 302864
rect 348844 302824 369216 302852
rect 348844 302812 348850 302824
rect 369210 302812 369216 302824
rect 369268 302812 369274 302864
rect 215110 302744 215116 302796
rect 215168 302784 215174 302796
rect 285122 302784 285128 302796
rect 215168 302756 285128 302784
rect 215168 302744 215174 302756
rect 285122 302744 285128 302756
rect 285180 302744 285186 302796
rect 352006 302744 352012 302796
rect 352064 302784 352070 302796
rect 373074 302784 373080 302796
rect 352064 302756 373080 302784
rect 352064 302744 352070 302756
rect 373074 302744 373080 302756
rect 373132 302744 373138 302796
rect 172330 302676 172336 302728
rect 172388 302716 172394 302728
rect 234798 302716 234804 302728
rect 172388 302688 234804 302716
rect 172388 302676 172394 302688
rect 234798 302676 234804 302688
rect 234856 302676 234862 302728
rect 236454 302676 236460 302728
rect 236512 302716 236518 302728
rect 237282 302716 237288 302728
rect 236512 302688 237288 302716
rect 236512 302676 236518 302688
rect 237282 302676 237288 302688
rect 237340 302676 237346 302728
rect 348050 302676 348056 302728
rect 348108 302716 348114 302728
rect 358170 302716 358176 302728
rect 348108 302688 358176 302716
rect 348108 302676 348114 302688
rect 358170 302676 358176 302688
rect 358228 302676 358234 302728
rect 261018 302472 261024 302524
rect 261076 302512 261082 302524
rect 262122 302512 262128 302524
rect 261076 302484 262128 302512
rect 261076 302472 261082 302484
rect 262122 302472 262128 302484
rect 262180 302472 262186 302524
rect 339954 302268 339960 302320
rect 340012 302308 340018 302320
rect 340598 302308 340604 302320
rect 340012 302280 340604 302308
rect 340012 302268 340018 302280
rect 340598 302268 340604 302280
rect 340656 302268 340662 302320
rect 172422 302132 172428 302184
rect 172480 302172 172486 302184
rect 238662 302172 238668 302184
rect 172480 302144 238668 302172
rect 172480 302132 172486 302144
rect 238662 302132 238668 302144
rect 238720 302132 238726 302184
rect 219342 301588 219348 301640
rect 219400 301628 219406 301640
rect 290274 301628 290280 301640
rect 219400 301600 290280 301628
rect 219400 301588 219406 301600
rect 290274 301588 290280 301600
rect 290332 301588 290338 301640
rect 211982 301520 211988 301572
rect 212040 301560 212046 301572
rect 340414 301560 340420 301572
rect 212040 301532 340420 301560
rect 212040 301520 212046 301532
rect 340414 301520 340420 301532
rect 340472 301520 340478 301572
rect 213362 301452 213368 301504
rect 213420 301492 213426 301504
rect 341058 301492 341064 301504
rect 213420 301464 341064 301492
rect 213420 301452 213426 301464
rect 341058 301452 341064 301464
rect 341116 301452 341122 301504
rect 251358 301316 251364 301368
rect 251416 301356 251422 301368
rect 251634 301356 251640 301368
rect 251416 301328 251640 301356
rect 251416 301316 251422 301328
rect 251634 301316 251640 301328
rect 251692 301316 251698 301368
rect 97442 300772 97448 300824
rect 97500 300812 97506 300824
rect 248874 300812 248880 300824
rect 97500 300784 248880 300812
rect 97500 300772 97506 300784
rect 248874 300772 248880 300784
rect 248932 300772 248938 300824
rect 343726 300772 343732 300824
rect 343784 300812 343790 300824
rect 365070 300812 365076 300824
rect 343784 300784 365076 300812
rect 343784 300772 343790 300784
rect 365070 300772 365076 300784
rect 365128 300772 365134 300824
rect 97258 300704 97264 300756
rect 97316 300744 97322 300756
rect 247034 300744 247040 300756
rect 97316 300716 247040 300744
rect 97316 300704 97322 300716
rect 247034 300704 247040 300716
rect 247092 300704 247098 300756
rect 350534 300704 350540 300756
rect 350592 300744 350598 300756
rect 372706 300744 372712 300756
rect 350592 300716 372712 300744
rect 350592 300704 350598 300716
rect 372706 300704 372712 300716
rect 372764 300704 372770 300756
rect 99374 300636 99380 300688
rect 99432 300676 99438 300688
rect 248598 300676 248604 300688
rect 99432 300648 248604 300676
rect 99432 300636 99438 300648
rect 248598 300636 248604 300648
rect 248656 300636 248662 300688
rect 349154 300636 349160 300688
rect 349212 300676 349218 300688
rect 373258 300676 373264 300688
rect 349212 300648 373264 300676
rect 349212 300636 349218 300648
rect 373258 300636 373264 300648
rect 373316 300636 373322 300688
rect 97718 300568 97724 300620
rect 97776 300608 97782 300620
rect 244550 300608 244556 300620
rect 97776 300580 244556 300608
rect 97776 300568 97782 300580
rect 244550 300568 244556 300580
rect 244608 300568 244614 300620
rect 342622 300568 342628 300620
rect 342680 300608 342686 300620
rect 369302 300608 369308 300620
rect 342680 300580 369308 300608
rect 342680 300568 342686 300580
rect 369302 300568 369308 300580
rect 369360 300568 369366 300620
rect 97810 300500 97816 300552
rect 97868 300540 97874 300552
rect 242802 300540 242808 300552
rect 97868 300512 242808 300540
rect 97868 300500 97874 300512
rect 242802 300500 242808 300512
rect 242860 300500 242866 300552
rect 342438 300500 342444 300552
rect 342496 300540 342502 300552
rect 371418 300540 371424 300552
rect 342496 300512 371424 300540
rect 342496 300500 342502 300512
rect 371418 300500 371424 300512
rect 371476 300500 371482 300552
rect 99006 300432 99012 300484
rect 99064 300472 99070 300484
rect 243078 300472 243084 300484
rect 99064 300444 243084 300472
rect 99064 300432 99070 300444
rect 243078 300432 243084 300444
rect 243136 300432 243142 300484
rect 341150 300432 341156 300484
rect 341208 300472 341214 300484
rect 370314 300472 370320 300484
rect 341208 300444 370320 300472
rect 341208 300432 341214 300444
rect 370314 300432 370320 300444
rect 370372 300432 370378 300484
rect 97626 300364 97632 300416
rect 97684 300404 97690 300416
rect 241974 300404 241980 300416
rect 97684 300376 241980 300404
rect 97684 300364 97690 300376
rect 241974 300364 241980 300376
rect 242032 300364 242038 300416
rect 343634 300364 343640 300416
rect 343692 300404 343698 300416
rect 372798 300404 372804 300416
rect 343692 300376 372804 300404
rect 343692 300364 343698 300376
rect 372798 300364 372804 300376
rect 372856 300364 372862 300416
rect 99466 300296 99472 300348
rect 99524 300336 99530 300348
rect 240594 300336 240600 300348
rect 99524 300308 240600 300336
rect 99524 300296 99530 300308
rect 240594 300296 240600 300308
rect 240652 300296 240658 300348
rect 342530 300296 342536 300348
rect 342588 300336 342594 300348
rect 373166 300336 373172 300348
rect 342588 300308 373172 300336
rect 342588 300296 342594 300308
rect 373166 300296 373172 300308
rect 373224 300296 373230 300348
rect 97350 300228 97356 300280
rect 97408 300268 97414 300280
rect 237374 300268 237380 300280
rect 97408 300240 237380 300268
rect 97408 300228 97414 300240
rect 237374 300228 237380 300240
rect 237432 300228 237438 300280
rect 343358 300228 343364 300280
rect 343416 300268 343422 300280
rect 371786 300268 371792 300280
rect 343416 300240 371792 300268
rect 343416 300228 343422 300240
rect 371786 300228 371792 300240
rect 371844 300228 371850 300280
rect 99834 300160 99840 300212
rect 99892 300200 99898 300212
rect 238938 300200 238944 300212
rect 99892 300172 238944 300200
rect 99892 300160 99898 300172
rect 238938 300160 238944 300172
rect 238996 300160 239002 300212
rect 339678 300160 339684 300212
rect 339736 300200 339742 300212
rect 372890 300200 372896 300212
rect 339736 300172 372896 300200
rect 339736 300160 339742 300172
rect 372890 300160 372896 300172
rect 372948 300160 372954 300212
rect 99190 300092 99196 300144
rect 99248 300132 99254 300144
rect 237190 300132 237196 300144
rect 99248 300104 237196 300132
rect 99248 300092 99254 300104
rect 237190 300092 237196 300104
rect 237248 300092 237254 300144
rect 294138 300092 294144 300144
rect 294196 300132 294202 300144
rect 369026 300132 369032 300144
rect 294196 300104 369032 300132
rect 294196 300092 294202 300104
rect 369026 300092 369032 300104
rect 369084 300092 369090 300144
rect 98914 300024 98920 300076
rect 98972 300064 98978 300076
rect 233418 300064 233424 300076
rect 98972 300036 233424 300064
rect 98972 300024 98978 300036
rect 233418 300024 233424 300036
rect 233476 300024 233482 300076
rect 350626 300024 350632 300076
rect 350684 300064 350690 300076
rect 371878 300064 371884 300076
rect 350684 300036 371884 300064
rect 350684 300024 350690 300036
rect 371878 300024 371884 300036
rect 371936 300024 371942 300076
rect 217962 299956 217968 300008
rect 218020 299996 218026 300008
rect 292666 299996 292672 300008
rect 218020 299968 292672 299996
rect 218020 299956 218026 299968
rect 292666 299956 292672 299968
rect 292724 299956 292730 300008
rect 350718 299956 350724 300008
rect 350776 299996 350782 300008
rect 371694 299996 371700 300008
rect 350776 299968 371700 299996
rect 350776 299956 350782 299968
rect 371694 299956 371700 299968
rect 371752 299956 371758 300008
rect 213546 299888 213552 299940
rect 213604 299928 213610 299940
rect 286042 299928 286048 299940
rect 213604 299900 286048 299928
rect 213604 299888 213610 299900
rect 286042 299888 286048 299900
rect 286100 299888 286106 299940
rect 350810 299888 350816 299940
rect 350868 299928 350874 299940
rect 371510 299928 371516 299940
rect 350868 299900 371516 299928
rect 350868 299888 350874 299900
rect 371510 299888 371516 299900
rect 371568 299888 371574 299940
rect 271138 299752 271144 299804
rect 271196 299792 271202 299804
rect 271598 299792 271604 299804
rect 271196 299764 271604 299792
rect 271196 299752 271202 299764
rect 271598 299752 271604 299764
rect 271656 299752 271662 299804
rect 97902 299412 97908 299464
rect 97960 299452 97966 299464
rect 241698 299452 241704 299464
rect 97960 299424 241704 299452
rect 97960 299412 97966 299424
rect 241698 299412 241704 299424
rect 241756 299412 241762 299464
rect 352650 299412 352656 299464
rect 352708 299452 352714 299464
rect 580166 299452 580172 299464
rect 352708 299424 580172 299452
rect 352708 299412 352714 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 98638 299344 98644 299396
rect 98696 299384 98702 299396
rect 239306 299384 239312 299396
rect 98696 299356 239312 299384
rect 98696 299344 98702 299356
rect 239306 299344 239312 299356
rect 239364 299344 239370 299396
rect 98822 299276 98828 299328
rect 98880 299316 98886 299328
rect 237466 299316 237472 299328
rect 98880 299288 237472 299316
rect 98880 299276 98886 299288
rect 237466 299276 237472 299288
rect 237524 299276 237530 299328
rect 98546 299208 98552 299260
rect 98604 299248 98610 299260
rect 236178 299248 236184 299260
rect 98604 299220 236184 299248
rect 98604 299208 98610 299220
rect 236178 299208 236184 299220
rect 236236 299208 236242 299260
rect 104526 299140 104532 299192
rect 104584 299180 104590 299192
rect 234706 299180 234712 299192
rect 104584 299152 234712 299180
rect 104584 299140 104590 299152
rect 234706 299140 234712 299152
rect 234764 299140 234770 299192
rect 114830 299072 114836 299124
rect 114888 299112 114894 299124
rect 242986 299112 242992 299124
rect 114888 299084 242992 299112
rect 114888 299072 114894 299084
rect 242986 299072 242992 299084
rect 243044 299072 243050 299124
rect 119982 299004 119988 299056
rect 120040 299044 120046 299056
rect 246114 299044 246120 299056
rect 120040 299016 246120 299044
rect 120040 299004 120046 299016
rect 246114 299004 246120 299016
rect 246172 299004 246178 299056
rect 125134 298936 125140 298988
rect 125192 298976 125198 298988
rect 239122 298976 239128 298988
rect 125192 298948 239128 298976
rect 125192 298936 125198 298948
rect 239122 298936 239128 298948
rect 239180 298936 239186 298988
rect 140590 298868 140596 298920
rect 140648 298908 140654 298920
rect 249886 298908 249892 298920
rect 140648 298880 249892 298908
rect 140648 298868 140654 298880
rect 249886 298868 249892 298880
rect 249944 298868 249950 298920
rect 156046 298800 156052 298852
rect 156104 298840 156110 298852
rect 250070 298840 250076 298852
rect 156104 298812 250076 298840
rect 156104 298800 156110 298812
rect 250070 298800 250076 298812
rect 250128 298800 250134 298852
rect 146938 298732 146944 298784
rect 146996 298772 147002 298784
rect 248690 298772 248696 298784
rect 146996 298744 248696 298772
rect 146996 298732 147002 298744
rect 248690 298732 248696 298744
rect 248748 298732 248754 298784
rect 333238 298732 333244 298784
rect 333296 298772 333302 298784
rect 538858 298772 538864 298784
rect 333296 298744 538864 298772
rect 333296 298732 333302 298744
rect 538858 298732 538864 298744
rect 538916 298732 538922 298784
rect 145742 298664 145748 298716
rect 145800 298704 145806 298716
rect 236270 298704 236276 298716
rect 145800 298676 236276 298704
rect 145800 298664 145806 298676
rect 236270 298664 236276 298676
rect 236328 298664 236334 298716
rect 161198 298596 161204 298648
rect 161256 298636 161262 298648
rect 247310 298636 247316 298648
rect 161256 298608 247316 298636
rect 161256 298596 161262 298608
rect 247310 298596 247316 298608
rect 247368 298596 247374 298648
rect 163774 298528 163780 298580
rect 163832 298568 163838 298580
rect 234522 298568 234528 298580
rect 163832 298540 234528 298568
rect 163832 298528 163838 298540
rect 234522 298528 234528 298540
rect 234580 298528 234586 298580
rect 158622 298052 158628 298104
rect 158680 298092 158686 298104
rect 169938 298092 169944 298104
rect 158680 298064 169944 298092
rect 158680 298052 158686 298064
rect 169938 298052 169944 298064
rect 169996 298052 170002 298104
rect 132862 297916 132868 297968
rect 132920 297956 132926 297968
rect 247218 297956 247224 297968
rect 132920 297928 247224 297956
rect 132920 297916 132926 297928
rect 247218 297916 247224 297928
rect 247276 297916 247282 297968
rect 122558 297848 122564 297900
rect 122616 297888 122622 297900
rect 236362 297888 236368 297900
rect 122616 297860 236368 297888
rect 122616 297848 122622 297860
rect 236362 297848 236368 297860
rect 236420 297848 236426 297900
rect 138014 297780 138020 297832
rect 138072 297820 138078 297832
rect 237558 297820 237564 297832
rect 138072 297792 237564 297820
rect 138072 297780 138078 297792
rect 237558 297780 237564 297792
rect 237616 297780 237622 297832
rect 130286 297712 130292 297764
rect 130344 297752 130350 297764
rect 146938 297752 146944 297764
rect 130344 297724 146944 297752
rect 130344 297712 130350 297724
rect 146938 297712 146944 297724
rect 146996 297712 147002 297764
rect 148318 297712 148324 297764
rect 148376 297752 148382 297764
rect 234798 297752 234804 297764
rect 148376 297724 234804 297752
rect 148376 297712 148382 297724
rect 234798 297712 234804 297724
rect 234856 297712 234862 297764
rect 100018 297644 100024 297696
rect 100076 297684 100082 297696
rect 172238 297684 172244 297696
rect 100076 297656 172244 297684
rect 100076 297644 100082 297656
rect 172238 297644 172244 297656
rect 172296 297644 172302 297696
rect 213730 297644 213736 297696
rect 213788 297684 213794 297696
rect 291746 297684 291752 297696
rect 213788 297656 291752 297684
rect 213788 297644 213794 297656
rect 291746 297644 291752 297656
rect 291804 297644 291810 297696
rect 107102 297576 107108 297628
rect 107160 297616 107166 297628
rect 170490 297616 170496 297628
rect 107160 297588 170496 297616
rect 107160 297576 107166 297588
rect 170490 297576 170496 297588
rect 170548 297576 170554 297628
rect 211706 297576 211712 297628
rect 211764 297616 211770 297628
rect 290366 297616 290372 297628
rect 211764 297588 290372 297616
rect 211764 297576 211770 297588
rect 290366 297576 290372 297588
rect 290424 297576 290430 297628
rect 109678 297508 109684 297560
rect 109736 297548 109742 297560
rect 170030 297548 170036 297560
rect 109736 297520 170036 297548
rect 109736 297508 109742 297520
rect 170030 297508 170036 297520
rect 170088 297508 170094 297560
rect 213270 297508 213276 297560
rect 213328 297548 213334 297560
rect 338390 297548 338396 297560
rect 213328 297520 338396 297548
rect 213328 297508 213334 297520
rect 338390 297508 338396 297520
rect 338448 297508 338454 297560
rect 112254 297440 112260 297492
rect 112312 297480 112318 297492
rect 172606 297480 172612 297492
rect 112312 297452 172612 297480
rect 112312 297440 112318 297452
rect 172606 297440 172612 297452
rect 172664 297440 172670 297492
rect 213178 297440 213184 297492
rect 213236 297480 213242 297492
rect 339586 297480 339592 297492
rect 213236 297452 339592 297480
rect 213236 297440 213242 297452
rect 339586 297440 339592 297452
rect 339644 297440 339650 297492
rect 135438 297372 135444 297424
rect 135496 297412 135502 297424
rect 171686 297412 171692 297424
rect 135496 297384 171692 297412
rect 135496 297372 135502 297384
rect 171686 297372 171692 297384
rect 171744 297372 171750 297424
rect 212258 297372 212264 297424
rect 212316 297412 212322 297424
rect 291930 297412 291936 297424
rect 212316 297384 291936 297412
rect 212316 297372 212322 297384
rect 291930 297372 291936 297384
rect 291988 297372 291994 297424
rect 337286 297372 337292 297424
rect 337344 297412 337350 297424
rect 567838 297412 567844 297424
rect 337344 297384 567844 297412
rect 337344 297372 337350 297384
rect 567838 297372 567844 297384
rect 567896 297372 567902 297424
rect 143166 297304 143172 297356
rect 143224 297344 143230 297356
rect 172330 297344 172336 297356
rect 143224 297316 172336 297344
rect 143224 297304 143230 297316
rect 172330 297304 172336 297316
rect 172388 297304 172394 297356
rect 213638 297304 213644 297356
rect 213696 297344 213702 297356
rect 289998 297344 290004 297356
rect 213696 297316 290004 297344
rect 213696 297304 213702 297316
rect 289998 297304 290004 297316
rect 290056 297304 290062 297356
rect 215938 297236 215944 297288
rect 215996 297276 216002 297288
rect 291470 297276 291476 297288
rect 215996 297248 291476 297276
rect 215996 297236 216002 297248
rect 291470 297236 291476 297248
rect 291528 297236 291534 297288
rect 218790 297168 218796 297220
rect 218848 297208 218854 297220
rect 290182 297208 290188 297220
rect 218848 297180 290188 297208
rect 218848 297168 218854 297180
rect 290182 297168 290188 297180
rect 290240 297168 290246 297220
rect 98730 297100 98736 297152
rect 98788 297140 98794 297152
rect 245838 297140 245844 297152
rect 98788 297112 245844 297140
rect 98788 297100 98794 297112
rect 245838 297100 245844 297112
rect 245896 297100 245902 297152
rect 101950 297032 101956 297084
rect 102008 297072 102014 297084
rect 247494 297072 247500 297084
rect 102008 297044 247500 297072
rect 102008 297032 102014 297044
rect 247494 297032 247500 297044
rect 247552 297032 247558 297084
rect 99098 296624 99104 296676
rect 99156 296664 99162 296676
rect 240318 296664 240324 296676
rect 99156 296636 240324 296664
rect 99156 296624 99162 296636
rect 240318 296624 240324 296636
rect 240376 296624 240382 296676
rect 117314 296556 117320 296608
rect 117372 296596 117378 296608
rect 243170 296596 243176 296608
rect 117372 296568 243176 296596
rect 117372 296556 117378 296568
rect 243170 296556 243176 296568
rect 243228 296556 243234 296608
rect 126974 296488 126980 296540
rect 127032 296528 127038 296540
rect 247126 296528 247132 296540
rect 127032 296500 247132 296528
rect 127032 296488 127038 296500
rect 247126 296488 247132 296500
rect 247184 296488 247190 296540
rect 153194 296420 153200 296472
rect 153252 296460 153258 296472
rect 247402 296460 247408 296472
rect 153252 296432 247408 296460
rect 153252 296420 153258 296432
rect 247402 296420 247408 296432
rect 247460 296420 247466 296472
rect 149054 296080 149060 296132
rect 149112 296120 149118 296132
rect 273346 296120 273352 296132
rect 149112 296092 273352 296120
rect 149112 296080 149118 296092
rect 273346 296080 273352 296092
rect 273404 296080 273410 296132
rect 143534 296012 143540 296064
rect 143592 296052 143598 296064
rect 272610 296052 272616 296064
rect 143592 296024 272616 296052
rect 143592 296012 143598 296024
rect 272610 296012 272616 296024
rect 272668 296012 272674 296064
rect 125594 295944 125600 295996
rect 125652 295984 125658 295996
rect 269666 295984 269672 295996
rect 125652 295956 269672 295984
rect 125652 295944 125658 295956
rect 269666 295944 269672 295956
rect 269724 295944 269730 295996
rect 210878 295196 210884 295248
rect 210936 295236 210942 295248
rect 283282 295236 283288 295248
rect 210936 295208 283288 295236
rect 210936 295196 210942 295208
rect 283282 295196 283288 295208
rect 283340 295196 283346 295248
rect 217870 295128 217876 295180
rect 217928 295168 217934 295180
rect 293034 295168 293040 295180
rect 217928 295140 293040 295168
rect 217928 295128 217934 295140
rect 293034 295128 293040 295140
rect 293092 295128 293098 295180
rect 215846 295060 215852 295112
rect 215904 295100 215910 295112
rect 292942 295100 292948 295112
rect 215904 295072 292948 295100
rect 215904 295060 215910 295072
rect 292942 295060 292948 295072
rect 293000 295060 293006 295112
rect 214374 294992 214380 295044
rect 214432 295032 214438 295044
rect 292574 295032 292580 295044
rect 214432 295004 292580 295032
rect 214432 294992 214438 295004
rect 292574 294992 292580 295004
rect 292632 294992 292638 295044
rect 213086 294924 213092 294976
rect 213144 294964 213150 294976
rect 291654 294964 291660 294976
rect 213144 294936 291660 294964
rect 213144 294924 213150 294936
rect 291654 294924 291660 294936
rect 291712 294924 291718 294976
rect 214466 294856 214472 294908
rect 214524 294896 214530 294908
rect 292758 294896 292764 294908
rect 214524 294868 292764 294896
rect 214524 294856 214530 294868
rect 292758 294856 292764 294868
rect 292816 294856 292822 294908
rect 211614 294788 211620 294840
rect 211672 294828 211678 294840
rect 291562 294828 291568 294840
rect 211672 294800 291568 294828
rect 211672 294788 211678 294800
rect 291562 294788 291568 294800
rect 291620 294788 291626 294840
rect 212994 294720 213000 294772
rect 213052 294760 213058 294772
rect 292850 294760 292856 294772
rect 213052 294732 292856 294760
rect 213052 294720 213058 294732
rect 292850 294720 292856 294732
rect 292908 294720 292914 294772
rect 164234 294652 164240 294704
rect 164292 294692 164298 294704
rect 275462 294692 275468 294704
rect 164292 294664 275468 294692
rect 164292 294652 164298 294664
rect 275462 294652 275468 294664
rect 275520 294652 275526 294704
rect 139394 294584 139400 294636
rect 139452 294624 139458 294636
rect 271138 294624 271144 294636
rect 139452 294596 271144 294624
rect 139452 294584 139458 294596
rect 271138 294584 271144 294596
rect 271196 294584 271202 294636
rect 321922 294584 321928 294636
rect 321980 294624 321986 294636
rect 471238 294624 471244 294636
rect 321980 294596 471244 294624
rect 321980 294584 321986 294596
rect 471238 294584 471244 294596
rect 471296 294584 471302 294636
rect 217686 293360 217692 293412
rect 217744 293400 217750 293412
rect 341518 293400 341524 293412
rect 217744 293372 341524 293400
rect 217744 293360 217750 293372
rect 341518 293360 341524 293372
rect 341576 293360 341582 293412
rect 150434 293292 150440 293344
rect 150492 293332 150498 293344
rect 273254 293332 273260 293344
rect 150492 293304 273260 293332
rect 150492 293292 150498 293304
rect 273254 293292 273260 293304
rect 273312 293292 273318 293344
rect 333146 293292 333152 293344
rect 333204 293332 333210 293344
rect 543734 293332 543740 293344
rect 333204 293304 543740 293332
rect 333204 293292 333210 293304
rect 543734 293292 543740 293304
rect 543792 293292 543798 293344
rect 64874 293224 64880 293276
rect 64932 293264 64938 293276
rect 260834 293264 260840 293276
rect 64932 293236 260840 293264
rect 64932 293224 64938 293236
rect 260834 293224 260840 293236
rect 260892 293224 260898 293276
rect 337194 293224 337200 293276
rect 337252 293264 337258 293276
rect 571978 293264 571984 293276
rect 337252 293236 571984 293264
rect 337252 293224 337258 293236
rect 571978 293224 571984 293236
rect 572036 293224 572042 293276
rect 184198 291864 184204 291916
rect 184256 291904 184262 291916
rect 276382 291904 276388 291916
rect 184256 291876 276388 291904
rect 184256 291864 184262 291876
rect 276382 291864 276388 291876
rect 276440 291864 276446 291916
rect 315206 291864 315212 291916
rect 315264 291904 315270 291916
rect 422938 291904 422944 291916
rect 315264 291876 422944 291904
rect 315264 291864 315270 291876
rect 422938 291864 422944 291876
rect 422996 291864 423002 291916
rect 128354 291796 128360 291848
rect 128412 291836 128418 291848
rect 269758 291836 269764 291848
rect 128412 291808 269764 291836
rect 128412 291796 128418 291808
rect 269758 291796 269764 291808
rect 269816 291796 269822 291848
rect 333054 291796 333060 291848
rect 333112 291836 333118 291848
rect 547874 291836 547880 291848
rect 333112 291808 547880 291836
rect 333112 291796 333118 291808
rect 547874 291796 547880 291808
rect 547932 291796 547938 291848
rect 132494 290504 132500 290556
rect 132552 290544 132558 290556
rect 271230 290544 271236 290556
rect 132552 290516 271236 290544
rect 132552 290504 132558 290516
rect 271230 290504 271236 290516
rect 271288 290504 271294 290556
rect 22738 290436 22744 290488
rect 22796 290476 22802 290488
rect 254394 290476 254400 290488
rect 22796 290448 254400 290476
rect 22796 290436 22802 290448
rect 254394 290436 254400 290448
rect 254452 290436 254458 290488
rect 316494 290436 316500 290488
rect 316552 290476 316558 290488
rect 431954 290476 431960 290488
rect 316552 290448 431960 290476
rect 316552 290436 316558 290448
rect 431954 290436 431960 290448
rect 432012 290436 432018 290488
rect 312446 289416 312452 289468
rect 312504 289456 312510 289468
rect 407114 289456 407120 289468
rect 312504 289428 407120 289456
rect 312504 289416 312510 289428
rect 407114 289416 407120 289428
rect 407172 289416 407178 289468
rect 315114 289348 315120 289400
rect 315172 289388 315178 289400
rect 413278 289388 413284 289400
rect 315172 289360 413284 289388
rect 315172 289348 315178 289360
rect 413278 289348 413284 289360
rect 413336 289348 413342 289400
rect 312538 289280 312544 289332
rect 312596 289320 312602 289332
rect 411254 289320 411260 289332
rect 312596 289292 411260 289320
rect 312596 289280 312602 289292
rect 411254 289280 411260 289292
rect 411312 289280 411318 289332
rect 313918 289212 313924 289264
rect 313976 289252 313982 289264
rect 415394 289252 415400 289264
rect 313976 289224 415400 289252
rect 313976 289212 313982 289224
rect 415394 289212 415400 289224
rect 415452 289212 415458 289264
rect 313826 289144 313832 289196
rect 313884 289184 313890 289196
rect 418154 289184 418160 289196
rect 313884 289156 418160 289184
rect 313884 289144 313890 289156
rect 418154 289144 418160 289156
rect 418212 289144 418218 289196
rect 135254 289076 135260 289128
rect 135312 289116 135318 289128
rect 270954 289116 270960 289128
rect 135312 289088 270960 289116
rect 135312 289076 135318 289088
rect 270954 289076 270960 289088
rect 271012 289076 271018 289128
rect 337102 289076 337108 289128
rect 337160 289116 337166 289128
rect 575474 289116 575480 289128
rect 337160 289088 575480 289116
rect 337160 289076 337166 289088
rect 575474 289076 575480 289088
rect 575532 289076 575538 289128
rect 308306 287988 308312 288040
rect 308364 288028 308370 288040
rect 382274 288028 382280 288040
rect 308364 288000 382280 288028
rect 308364 287988 308370 288000
rect 382274 287988 382280 288000
rect 382332 287988 382338 288040
rect 309778 287920 309784 287972
rect 309836 287960 309842 287972
rect 386414 287960 386420 287972
rect 309836 287932 386420 287960
rect 309836 287920 309842 287932
rect 386414 287920 386420 287932
rect 386472 287920 386478 287972
rect 312630 287852 312636 287904
rect 312688 287892 312694 287904
rect 400214 287892 400220 287904
rect 312688 287864 400220 287892
rect 312688 287852 312694 287864
rect 400214 287852 400220 287864
rect 400272 287852 400278 287904
rect 146294 287784 146300 287836
rect 146352 287824 146358 287836
rect 272334 287824 272340 287836
rect 146352 287796 272340 287824
rect 146352 287784 146358 287796
rect 272334 287784 272340 287796
rect 272392 287784 272398 287836
rect 311066 287784 311072 287836
rect 311124 287824 311130 287836
rect 404354 287824 404360 287836
rect 311124 287796 404360 287824
rect 311124 287784 311130 287796
rect 404354 287784 404360 287796
rect 404412 287784 404418 287836
rect 71038 287716 71044 287768
rect 71096 287756 71102 287768
rect 261386 287756 261392 287768
rect 71096 287728 261392 287756
rect 71096 287716 71102 287728
rect 261386 287716 261392 287728
rect 261444 287716 261450 287768
rect 323670 287716 323676 287768
rect 323728 287756 323734 287768
rect 471974 287756 471980 287768
rect 323728 287728 471980 287756
rect 323728 287716 323734 287728
rect 471974 287716 471980 287728
rect 472032 287716 472038 287768
rect 39298 287648 39304 287700
rect 39356 287688 39362 287700
rect 257246 287688 257252 287700
rect 39356 287660 257252 287688
rect 39356 287648 39362 287660
rect 257246 287648 257252 287660
rect 257304 287648 257310 287700
rect 324866 287648 324872 287700
rect 324924 287688 324930 287700
rect 488534 287688 488540 287700
rect 324924 287660 488540 287688
rect 324924 287648 324930 287660
rect 488534 287648 488540 287660
rect 488592 287648 488598 287700
rect 306926 286628 306932 286680
rect 306984 286668 306990 286680
rect 375374 286668 375380 286680
rect 306984 286640 375380 286668
rect 306984 286628 306990 286640
rect 375374 286628 375380 286640
rect 375432 286628 375438 286680
rect 310974 286560 310980 286612
rect 311032 286600 311038 286612
rect 397454 286600 397460 286612
rect 311032 286572 397460 286600
rect 311032 286560 311038 286572
rect 397454 286560 397460 286572
rect 397512 286560 397518 286612
rect 313734 286492 313740 286544
rect 313792 286532 313798 286544
rect 416774 286532 416780 286544
rect 313792 286504 416780 286532
rect 313792 286492 313798 286504
rect 416774 286492 416780 286504
rect 416832 286492 416838 286544
rect 217778 286424 217784 286476
rect 217836 286464 217842 286476
rect 338206 286464 338212 286476
rect 217836 286436 338212 286464
rect 217836 286424 217842 286436
rect 338206 286424 338212 286436
rect 338264 286424 338270 286476
rect 153194 286356 153200 286408
rect 153252 286396 153258 286408
rect 273714 286396 273720 286408
rect 153252 286368 273720 286396
rect 153252 286356 153258 286368
rect 273714 286356 273720 286368
rect 273772 286356 273778 286408
rect 324774 286356 324780 286408
rect 324832 286396 324838 286408
rect 492674 286396 492680 286408
rect 324832 286368 492680 286396
rect 324832 286356 324838 286368
rect 492674 286356 492680 286368
rect 492732 286356 492738 286408
rect 12434 286288 12440 286340
rect 12492 286328 12498 286340
rect 253014 286328 253020 286340
rect 12492 286300 253020 286328
rect 12492 286288 12498 286300
rect 253014 286288 253020 286300
rect 253072 286288 253078 286340
rect 327626 286288 327632 286340
rect 327684 286328 327690 286340
rect 509234 286328 509240 286340
rect 327684 286300 509240 286328
rect 327684 286288 327690 286300
rect 509234 286288 509240 286300
rect 509292 286288 509298 286340
rect 308490 285200 308496 285252
rect 308548 285240 308554 285252
rect 372614 285240 372620 285252
rect 308548 285212 372620 285240
rect 308548 285200 308554 285212
rect 372614 285200 372620 285212
rect 372672 285200 372678 285252
rect 309686 285132 309692 285184
rect 309744 285172 309750 285184
rect 391934 285172 391940 285184
rect 309744 285144 391940 285172
rect 309744 285132 309750 285144
rect 391934 285132 391940 285144
rect 391992 285132 391998 285184
rect 157334 285064 157340 285116
rect 157392 285104 157398 285116
rect 275094 285104 275100 285116
rect 157392 285076 275100 285104
rect 157392 285064 157398 285076
rect 275094 285064 275100 285076
rect 275152 285064 275158 285116
rect 310882 285064 310888 285116
rect 310940 285104 310946 285116
rect 396074 285104 396080 285116
rect 310940 285076 396080 285104
rect 310940 285064 310946 285076
rect 396074 285064 396080 285076
rect 396132 285064 396138 285116
rect 135346 284996 135352 285048
rect 135404 285036 135410 285048
rect 270862 285036 270868 285048
rect 135404 285008 270868 285036
rect 135404 284996 135410 285008
rect 270862 284996 270868 285008
rect 270920 284996 270926 285048
rect 310790 284996 310796 285048
rect 310848 285036 310854 285048
rect 398834 285036 398840 285048
rect 310848 285008 398840 285036
rect 310848 284996 310854 285008
rect 398834 284996 398840 285008
rect 398892 284996 398898 285048
rect 103514 284928 103520 284980
rect 103572 284968 103578 284980
rect 266906 284968 266912 284980
rect 103572 284940 266912 284968
rect 103572 284928 103578 284940
rect 266906 284928 266912 284940
rect 266964 284928 266970 284980
rect 312354 284928 312360 284980
rect 312412 284968 312418 284980
rect 414014 284968 414020 284980
rect 312412 284940 414020 284968
rect 312412 284928 312418 284940
rect 414014 284928 414020 284940
rect 414072 284928 414078 284980
rect 218422 283772 218428 283824
rect 218480 283812 218486 283824
rect 283006 283812 283012 283824
rect 218480 283784 283012 283812
rect 218480 283772 218486 283784
rect 283006 283772 283012 283784
rect 283064 283772 283070 283824
rect 126974 283704 126980 283756
rect 127032 283744 127038 283756
rect 269482 283744 269488 283756
rect 127032 283716 269488 283744
rect 127032 283704 127038 283716
rect 269482 283704 269488 283716
rect 269540 283704 269546 283756
rect 308214 283704 308220 283756
rect 308272 283744 308278 283756
rect 378134 283744 378140 283756
rect 308272 283716 378140 283744
rect 308272 283704 308278 283716
rect 378134 283704 378140 283716
rect 378192 283704 378198 283756
rect 111794 283636 111800 283688
rect 111852 283676 111858 283688
rect 268286 283676 268292 283688
rect 111852 283648 268292 283676
rect 111852 283636 111858 283648
rect 268286 283636 268292 283648
rect 268344 283636 268350 283688
rect 308122 283636 308128 283688
rect 308180 283676 308186 283688
rect 385034 283676 385040 283688
rect 308180 283648 385040 283676
rect 308180 283636 308186 283648
rect 385034 283636 385040 283648
rect 385092 283636 385098 283688
rect 31754 283568 31760 283620
rect 31812 283608 31818 283620
rect 249058 283608 249064 283620
rect 31812 283580 249064 283608
rect 31812 283568 31818 283580
rect 249058 283568 249064 283580
rect 249116 283568 249122 283620
rect 309594 283568 309600 283620
rect 309652 283608 309658 283620
rect 389174 283608 389180 283620
rect 309652 283580 389180 283608
rect 309652 283568 309658 283580
rect 389174 283568 389180 283580
rect 389232 283568 389238 283620
rect 306742 282548 306748 282600
rect 306800 282588 306806 282600
rect 371234 282588 371240 282600
rect 306800 282560 371240 282588
rect 306800 282548 306806 282560
rect 371234 282548 371240 282560
rect 371292 282548 371298 282600
rect 306834 282480 306840 282532
rect 306892 282520 306898 282532
rect 373994 282520 374000 282532
rect 306892 282492 374000 282520
rect 306892 282480 306898 282492
rect 373994 282480 374000 282492
rect 374052 282480 374058 282532
rect 310698 282412 310704 282464
rect 310756 282452 310762 282464
rect 402974 282452 402980 282464
rect 310756 282424 402980 282452
rect 310756 282412 310762 282424
rect 402974 282412 402980 282424
rect 403032 282412 403038 282464
rect 217410 282344 217416 282396
rect 217468 282384 217474 282396
rect 342346 282384 342352 282396
rect 217468 282356 342352 282384
rect 217468 282344 217474 282356
rect 342346 282344 342352 282356
rect 342404 282344 342410 282396
rect 161474 282276 161480 282328
rect 161532 282316 161538 282328
rect 275002 282316 275008 282328
rect 161532 282288 275008 282316
rect 161532 282276 161538 282288
rect 275002 282276 275008 282288
rect 275060 282276 275066 282328
rect 321830 282276 321836 282328
rect 321888 282316 321894 282328
rect 475378 282316 475384 282328
rect 321888 282288 475384 282316
rect 321888 282276 321894 282288
rect 475378 282276 475384 282288
rect 475436 282276 475442 282328
rect 131114 282208 131120 282260
rect 131172 282248 131178 282260
rect 270770 282248 270776 282260
rect 131172 282220 270776 282248
rect 131172 282208 131178 282220
rect 270770 282208 270776 282220
rect 270828 282208 270834 282260
rect 330386 282208 330392 282260
rect 330444 282248 330450 282260
rect 524414 282248 524420 282260
rect 330444 282220 524420 282248
rect 330444 282208 330450 282220
rect 524414 282208 524420 282220
rect 524472 282208 524478 282260
rect 44174 282140 44180 282192
rect 44232 282180 44238 282192
rect 257154 282180 257160 282192
rect 44232 282152 257160 282180
rect 44232 282140 44238 282152
rect 257154 282140 257160 282152
rect 257212 282140 257218 282192
rect 337010 282140 337016 282192
rect 337068 282180 337074 282192
rect 574094 282180 574100 282192
rect 337068 282152 574100 282180
rect 337068 282140 337074 282152
rect 574094 282140 574100 282152
rect 574152 282140 574158 282192
rect 165614 280984 165620 281036
rect 165672 281024 165678 281036
rect 274910 281024 274916 281036
rect 165672 280996 274916 281024
rect 165672 280984 165678 280996
rect 274910 280984 274916 280996
rect 274968 280984 274974 281036
rect 315022 280984 315028 281036
rect 315080 281024 315086 281036
rect 426434 281024 426440 281036
rect 315080 280996 426440 281024
rect 315080 280984 315086 280996
rect 426434 280984 426440 280996
rect 426492 280984 426498 281036
rect 218698 280916 218704 280968
rect 218756 280956 218762 280968
rect 339954 280956 339960 280968
rect 218756 280928 339960 280956
rect 218756 280916 218762 280928
rect 339954 280916 339960 280928
rect 340012 280916 340018 280968
rect 140774 280848 140780 280900
rect 140832 280888 140838 280900
rect 272242 280888 272248 280900
rect 140832 280860 272248 280888
rect 140832 280848 140838 280860
rect 272242 280848 272248 280860
rect 272300 280848 272306 280900
rect 316402 280848 316408 280900
rect 316460 280888 316466 280900
rect 440234 280888 440240 280900
rect 316460 280860 440240 280888
rect 316460 280848 316466 280860
rect 440234 280848 440240 280860
rect 440292 280848 440298 280900
rect 110414 280780 110420 280832
rect 110472 280820 110478 280832
rect 268194 280820 268200 280832
rect 110472 280792 268200 280820
rect 110472 280780 110478 280792
rect 268194 280780 268200 280792
rect 268252 280780 268258 280832
rect 323486 280780 323492 280832
rect 323544 280820 323550 280832
rect 481634 280820 481640 280832
rect 323544 280792 481640 280820
rect 323544 280780 323550 280792
rect 481634 280780 481640 280792
rect 481692 280780 481698 280832
rect 181438 279692 181444 279744
rect 181496 279732 181502 279744
rect 277854 279732 277860 279744
rect 181496 279704 277860 279732
rect 181496 279692 181502 279704
rect 277854 279692 277860 279704
rect 277912 279692 277918 279744
rect 303982 279692 303988 279744
rect 304040 279732 304046 279744
rect 357434 279732 357440 279744
rect 304040 279704 357440 279732
rect 304040 279692 304046 279704
rect 357434 279692 357440 279704
rect 357492 279692 357498 279744
rect 168466 279624 168472 279676
rect 168524 279664 168530 279676
rect 276290 279664 276296 279676
rect 168524 279636 276296 279664
rect 168524 279624 168530 279636
rect 276290 279624 276296 279636
rect 276348 279624 276354 279676
rect 314930 279624 314936 279676
rect 314988 279664 314994 279676
rect 430574 279664 430580 279676
rect 314988 279636 430580 279664
rect 314988 279624 314994 279636
rect 430574 279624 430580 279636
rect 430632 279624 430638 279676
rect 102134 279556 102140 279608
rect 102192 279596 102198 279608
rect 266814 279596 266820 279608
rect 102192 279568 266820 279596
rect 102192 279556 102198 279568
rect 266814 279556 266820 279568
rect 266872 279556 266878 279608
rect 324682 279556 324688 279608
rect 324740 279596 324746 279608
rect 491294 279596 491300 279608
rect 324740 279568 491300 279596
rect 324740 279556 324746 279568
rect 491294 279556 491300 279568
rect 491352 279556 491358 279608
rect 45554 279488 45560 279540
rect 45612 279528 45618 279540
rect 246390 279528 246396 279540
rect 45612 279500 246396 279528
rect 45612 279488 45618 279500
rect 246390 279488 246396 279500
rect 246448 279488 246454 279540
rect 332962 279488 332968 279540
rect 333020 279528 333026 279540
rect 547966 279528 547972 279540
rect 333020 279500 547972 279528
rect 333020 279488 333026 279500
rect 547966 279488 547972 279500
rect 548024 279488 548030 279540
rect 13078 279420 13084 279472
rect 13136 279460 13142 279472
rect 252922 279460 252928 279472
rect 13136 279432 252928 279460
rect 13136 279420 13142 279432
rect 252922 279420 252928 279432
rect 252980 279420 252986 279472
rect 334526 279420 334532 279472
rect 334584 279460 334590 279472
rect 556154 279460 556160 279472
rect 334584 279432 556160 279460
rect 334584 279420 334590 279432
rect 556154 279420 556160 279432
rect 556212 279420 556218 279472
rect 308030 278196 308036 278248
rect 308088 278236 308094 278248
rect 382366 278236 382372 278248
rect 308088 278208 382372 278236
rect 308088 278196 308094 278208
rect 382366 278196 382372 278208
rect 382424 278196 382430 278248
rect 316310 278128 316316 278180
rect 316368 278168 316374 278180
rect 440326 278168 440332 278180
rect 316368 278140 440332 278168
rect 316368 278128 316374 278140
rect 440326 278128 440332 278140
rect 440384 278128 440390 278180
rect 147674 278060 147680 278112
rect 147732 278100 147738 278112
rect 273622 278100 273628 278112
rect 147732 278072 273628 278100
rect 147732 278060 147738 278072
rect 273622 278060 273628 278072
rect 273680 278060 273686 278112
rect 333330 278060 333336 278112
rect 333388 278100 333394 278112
rect 534074 278100 534080 278112
rect 333388 278072 534080 278100
rect 333388 278060 333394 278072
rect 534074 278060 534080 278072
rect 534132 278060 534138 278112
rect 117314 277992 117320 278044
rect 117372 278032 117378 278044
rect 251910 278032 251916 278044
rect 117372 278004 251916 278032
rect 117372 277992 117378 278004
rect 251910 277992 251916 278004
rect 251968 277992 251974 278044
rect 331766 277992 331772 278044
rect 331824 278032 331830 278044
rect 540974 278032 540980 278044
rect 331824 278004 540980 278032
rect 331824 277992 331830 278004
rect 540974 277992 540980 278004
rect 541032 277992 541038 278044
rect 318150 276972 318156 277024
rect 318208 277012 318214 277024
rect 433334 277012 433340 277024
rect 318208 276984 433340 277012
rect 318208 276972 318214 276984
rect 433334 276972 433340 276984
rect 433392 276972 433398 277024
rect 326154 276904 326160 276956
rect 326212 276944 326218 276956
rect 506566 276944 506572 276956
rect 326212 276916 506572 276944
rect 326212 276904 326218 276916
rect 506566 276904 506572 276916
rect 506624 276904 506630 276956
rect 151814 276836 151820 276888
rect 151872 276876 151878 276888
rect 273530 276876 273536 276888
rect 151872 276848 273536 276876
rect 151872 276836 151878 276848
rect 273530 276836 273536 276848
rect 273588 276836 273594 276888
rect 327534 276836 327540 276888
rect 327592 276876 327598 276888
rect 511258 276876 511264 276888
rect 327592 276848 511264 276876
rect 327592 276836 327598 276848
rect 511258 276836 511264 276848
rect 511316 276836 511322 276888
rect 106274 276768 106280 276820
rect 106332 276808 106338 276820
rect 266722 276808 266728 276820
rect 106332 276780 266728 276808
rect 106332 276768 106338 276780
rect 266722 276768 266728 276780
rect 266780 276768 266786 276820
rect 330294 276768 330300 276820
rect 330352 276808 330358 276820
rect 531314 276808 531320 276820
rect 330352 276780 531320 276808
rect 330352 276768 330358 276780
rect 531314 276768 531320 276780
rect 531372 276768 531378 276820
rect 84194 276700 84200 276752
rect 84252 276740 84258 276752
rect 264146 276740 264152 276752
rect 84252 276712 264152 276740
rect 84252 276700 84258 276712
rect 264146 276700 264152 276712
rect 264204 276700 264210 276752
rect 331674 276700 331680 276752
rect 331732 276740 331738 276752
rect 542354 276740 542360 276752
rect 331732 276712 542360 276740
rect 331732 276700 331738 276712
rect 542354 276700 542360 276712
rect 542412 276700 542418 276752
rect 71774 276632 71780 276684
rect 71832 276672 71838 276684
rect 261294 276672 261300 276684
rect 71832 276644 261300 276672
rect 71832 276632 71838 276644
rect 261294 276632 261300 276644
rect 261352 276632 261358 276684
rect 332870 276632 332876 276684
rect 332928 276672 332934 276684
rect 546494 276672 546500 276684
rect 332928 276644 546500 276672
rect 332928 276632 332934 276644
rect 546494 276632 546500 276644
rect 546552 276632 546558 276684
rect 309502 275612 309508 275664
rect 309560 275652 309566 275664
rect 393314 275652 393320 275664
rect 309560 275624 393320 275652
rect 309560 275612 309566 275624
rect 393314 275612 393320 275624
rect 393372 275612 393378 275664
rect 313642 275544 313648 275596
rect 313700 275584 313706 275596
rect 419534 275584 419540 275596
rect 313700 275556 419540 275584
rect 313700 275544 313706 275556
rect 419534 275544 419540 275556
rect 419592 275544 419598 275596
rect 313550 275476 313556 275528
rect 313608 275516 313614 275528
rect 423766 275516 423772 275528
rect 313608 275488 423772 275516
rect 313608 275476 313614 275488
rect 423766 275476 423772 275488
rect 423824 275476 423830 275528
rect 316218 275408 316224 275460
rect 316276 275448 316282 275460
rect 434714 275448 434720 275460
rect 316276 275420 434720 275448
rect 316276 275408 316282 275420
rect 434714 275408 434720 275420
rect 434772 275408 434778 275460
rect 184934 275340 184940 275392
rect 184992 275380 184998 275392
rect 278130 275380 278136 275392
rect 184992 275352 278136 275380
rect 184992 275340 184998 275352
rect 278130 275340 278136 275352
rect 278188 275340 278194 275392
rect 326062 275340 326068 275392
rect 326120 275380 326126 275392
rect 498194 275380 498200 275392
rect 326120 275352 498200 275380
rect 326120 275340 326126 275352
rect 498194 275340 498200 275352
rect 498252 275340 498258 275392
rect 129734 275272 129740 275324
rect 129792 275312 129798 275324
rect 270678 275312 270684 275324
rect 129792 275284 270684 275312
rect 129792 275272 129798 275284
rect 270678 275272 270684 275284
rect 270736 275272 270742 275324
rect 330202 275272 330208 275324
rect 330260 275312 330266 275324
rect 527174 275312 527180 275324
rect 330260 275284 527180 275312
rect 330260 275272 330266 275284
rect 527174 275272 527180 275284
rect 527232 275272 527238 275324
rect 313458 274252 313464 274304
rect 313516 274292 313522 274304
rect 415486 274292 415492 274304
rect 313516 274264 415492 274292
rect 313516 274252 313522 274264
rect 415486 274252 415492 274264
rect 415544 274252 415550 274304
rect 320818 274184 320824 274236
rect 320876 274224 320882 274236
rect 469214 274224 469220 274236
rect 320876 274196 469220 274224
rect 320876 274184 320882 274196
rect 469214 274184 469220 274196
rect 469272 274184 469278 274236
rect 321738 274116 321744 274168
rect 321796 274156 321802 274168
rect 473446 274156 473452 274168
rect 321796 274128 473452 274156
rect 321796 274116 321802 274128
rect 473446 274116 473452 274128
rect 473504 274116 473510 274168
rect 127066 274048 127072 274100
rect 127124 274088 127130 274100
rect 269390 274088 269396 274100
rect 127124 274060 269396 274088
rect 127124 274048 127130 274060
rect 269390 274048 269396 274060
rect 269448 274048 269454 274100
rect 323394 274048 323400 274100
rect 323452 274088 323458 274100
rect 476758 274088 476764 274100
rect 323452 274060 476764 274088
rect 323452 274048 323458 274060
rect 476758 274048 476764 274060
rect 476816 274048 476822 274100
rect 85574 273980 85580 274032
rect 85632 274020 85638 274032
rect 264054 274020 264060 274032
rect 85632 273992 264060 274020
rect 85632 273980 85638 273992
rect 264054 273980 264060 273992
rect 264112 273980 264118 274032
rect 329006 273980 329012 274032
rect 329064 274020 329070 274032
rect 516134 274020 516140 274032
rect 329064 273992 516140 274020
rect 329064 273980 329070 273992
rect 516134 273980 516140 273992
rect 516192 273980 516198 274032
rect 39390 273912 39396 273964
rect 39448 273952 39454 273964
rect 255774 273952 255780 273964
rect 39448 273924 255780 273952
rect 39448 273912 39454 273924
rect 255774 273912 255780 273924
rect 255832 273912 255838 273964
rect 331582 273912 331588 273964
rect 331640 273952 331646 273964
rect 538214 273952 538220 273964
rect 331640 273924 538220 273952
rect 331640 273912 331646 273924
rect 538214 273912 538220 273924
rect 538272 273912 538278 273964
rect 355318 273164 355324 273216
rect 355376 273204 355382 273216
rect 579982 273204 579988 273216
rect 355376 273176 579988 273204
rect 355376 273164 355382 273176
rect 579982 273164 579988 273176
rect 580040 273164 580046 273216
rect 166994 272688 167000 272740
rect 167052 272728 167058 272740
rect 276198 272728 276204 272740
rect 167052 272700 276204 272728
rect 167052 272688 167058 272700
rect 276198 272688 276204 272700
rect 276256 272688 276262 272740
rect 312262 272688 312268 272740
rect 312320 272728 312326 272740
rect 407206 272728 407212 272740
rect 312320 272700 407212 272728
rect 312320 272688 312326 272700
rect 407206 272688 407212 272700
rect 407264 272688 407270 272740
rect 88334 272620 88340 272672
rect 88392 272660 88398 272672
rect 263962 272660 263968 272672
rect 88392 272632 263968 272660
rect 88392 272620 88398 272632
rect 263962 272620 263968 272632
rect 264020 272620 264026 272672
rect 312170 272620 312176 272672
rect 312228 272660 312234 272672
rect 412634 272660 412640 272672
rect 312228 272632 412640 272660
rect 312228 272620 312234 272632
rect 412634 272620 412640 272632
rect 412692 272620 412698 272672
rect 66254 272552 66260 272604
rect 66312 272592 66318 272604
rect 261202 272592 261208 272604
rect 66312 272564 261208 272592
rect 66312 272552 66318 272564
rect 261202 272552 261208 272564
rect 261260 272552 261266 272604
rect 319530 272552 319536 272604
rect 319588 272592 319594 272604
rect 449894 272592 449900 272604
rect 319588 272564 449900 272592
rect 319588 272552 319594 272564
rect 449894 272552 449900 272564
rect 449952 272552 449958 272604
rect 2774 272484 2780 272536
rect 2832 272524 2838 272536
rect 251450 272524 251456 272536
rect 2832 272496 251456 272524
rect 2832 272484 2838 272496
rect 251450 272484 251456 272496
rect 251508 272484 251514 272536
rect 335998 272484 336004 272536
rect 336056 272524 336062 272536
rect 569954 272524 569960 272536
rect 336056 272496 569960 272524
rect 336056 272484 336062 272496
rect 569954 272484 569960 272496
rect 570012 272484 570018 272536
rect 209774 271396 209780 271448
rect 209832 271436 209838 271448
rect 282086 271436 282092 271448
rect 209832 271408 282092 271436
rect 209832 271396 209838 271408
rect 282086 271396 282092 271408
rect 282144 271396 282150 271448
rect 312078 271396 312084 271448
rect 312136 271436 312142 271448
rect 408494 271436 408500 271448
rect 312136 271408 408500 271436
rect 312136 271396 312142 271408
rect 408494 271396 408500 271408
rect 408552 271396 408558 271448
rect 205634 271328 205640 271380
rect 205692 271368 205698 271380
rect 282178 271368 282184 271380
rect 205692 271340 282184 271368
rect 205692 271328 205698 271340
rect 282178 271328 282184 271340
rect 282236 271328 282242 271380
rect 320726 271328 320732 271380
rect 320784 271368 320790 271380
rect 465074 271368 465080 271380
rect 320784 271340 465080 271368
rect 320784 271328 320790 271340
rect 465074 271328 465080 271340
rect 465132 271328 465138 271380
rect 151906 271260 151912 271312
rect 151964 271300 151970 271312
rect 273438 271300 273444 271312
rect 151964 271272 273444 271300
rect 151964 271260 151970 271272
rect 273438 271260 273444 271272
rect 273496 271260 273502 271312
rect 323302 271260 323308 271312
rect 323360 271300 323366 271312
rect 484394 271300 484400 271312
rect 323360 271272 484400 271300
rect 323360 271260 323366 271272
rect 484394 271260 484400 271272
rect 484452 271260 484458 271312
rect 143626 271192 143632 271244
rect 143684 271232 143690 271244
rect 272150 271232 272156 271244
rect 143684 271204 272156 271232
rect 143684 271192 143690 271204
rect 272150 271192 272156 271204
rect 272208 271192 272214 271244
rect 330110 271192 330116 271244
rect 330168 271232 330174 271244
rect 528554 271232 528560 271244
rect 330168 271204 528560 271232
rect 330168 271192 330174 271204
rect 528554 271192 528560 271204
rect 528612 271192 528618 271244
rect 81434 271124 81440 271176
rect 81492 271164 81498 271176
rect 257338 271164 257344 271176
rect 81492 271136 257344 271164
rect 81492 271124 81498 271136
rect 257338 271124 257344 271136
rect 257396 271124 257402 271176
rect 332778 271124 332784 271176
rect 332836 271164 332842 271176
rect 552014 271164 552020 271176
rect 332836 271136 552020 271164
rect 332836 271124 332842 271136
rect 552014 271124 552020 271136
rect 552072 271124 552078 271176
rect 198734 270172 198740 270224
rect 198792 270212 198798 270224
rect 278038 270212 278044 270224
rect 198792 270184 278044 270212
rect 198792 270172 198798 270184
rect 278038 270172 278044 270184
rect 278096 270172 278102 270224
rect 194594 270104 194600 270156
rect 194652 270144 194658 270156
rect 275278 270144 275284 270156
rect 194652 270116 275284 270144
rect 194652 270104 194658 270116
rect 275278 270104 275284 270116
rect 275336 270104 275342 270156
rect 310606 270104 310612 270156
rect 310664 270144 310670 270156
rect 401594 270144 401600 270156
rect 310664 270116 401600 270144
rect 310664 270104 310670 270116
rect 401594 270104 401600 270116
rect 401652 270104 401658 270156
rect 133874 270036 133880 270088
rect 133932 270076 133938 270088
rect 270586 270076 270592 270088
rect 133932 270048 270592 270076
rect 133932 270036 133938 270048
rect 270586 270036 270592 270048
rect 270644 270036 270650 270088
rect 319438 270036 319444 270088
rect 319496 270076 319502 270088
rect 458174 270076 458180 270088
rect 319496 270048 458180 270076
rect 319496 270036 319502 270048
rect 458174 270036 458180 270048
rect 458232 270036 458238 270088
rect 124214 269968 124220 270020
rect 124272 270008 124278 270020
rect 269298 270008 269304 270020
rect 124272 269980 269304 270008
rect 124272 269968 124278 269980
rect 269298 269968 269304 269980
rect 269356 269968 269362 270020
rect 320634 269968 320640 270020
rect 320692 270008 320698 270020
rect 465166 270008 465172 270020
rect 320692 269980 465172 270008
rect 320692 269968 320698 269980
rect 465166 269968 465172 269980
rect 465224 269968 465230 270020
rect 107654 269900 107660 269952
rect 107712 269940 107718 269952
rect 266630 269940 266636 269952
rect 107712 269912 266636 269940
rect 107712 269900 107718 269912
rect 266630 269900 266636 269912
rect 266688 269900 266694 269952
rect 324590 269900 324596 269952
rect 324648 269940 324654 269952
rect 495434 269940 495440 269952
rect 324648 269912 495440 269940
rect 324648 269900 324654 269912
rect 495434 269900 495440 269912
rect 495492 269900 495498 269952
rect 99374 269832 99380 269884
rect 99432 269872 99438 269884
rect 265618 269872 265624 269884
rect 99432 269844 265624 269872
rect 99432 269832 99438 269844
rect 265618 269832 265624 269844
rect 265676 269832 265682 269884
rect 327442 269832 327448 269884
rect 327500 269872 327506 269884
rect 504358 269872 504364 269884
rect 327500 269844 504364 269872
rect 327500 269832 327506 269844
rect 504358 269832 504364 269844
rect 504416 269832 504422 269884
rect 17954 269764 17960 269816
rect 18012 269804 18018 269816
rect 252830 269804 252836 269816
rect 18012 269776 252836 269804
rect 18012 269764 18018 269776
rect 252830 269764 252836 269776
rect 252888 269764 252894 269816
rect 334434 269764 334440 269816
rect 334492 269804 334498 269816
rect 558914 269804 558920 269816
rect 334492 269776 558920 269804
rect 334492 269764 334498 269776
rect 558914 269764 558920 269776
rect 558972 269764 558978 269816
rect 201494 268676 201500 268728
rect 201552 268716 201558 268728
rect 280522 268716 280528 268728
rect 201552 268688 280528 268716
rect 201552 268676 201558 268688
rect 280522 268676 280528 268688
rect 280580 268676 280586 268728
rect 310514 268676 310520 268728
rect 310572 268716 310578 268728
rect 398926 268716 398932 268728
rect 310572 268688 398932 268716
rect 310572 268676 310578 268688
rect 398926 268676 398932 268688
rect 398984 268676 398990 268728
rect 191834 268608 191840 268660
rect 191892 268648 191898 268660
rect 279326 268648 279332 268660
rect 191892 268620 279332 268648
rect 191892 268608 191898 268620
rect 279326 268608 279332 268620
rect 279384 268608 279390 268660
rect 317966 268608 317972 268660
rect 318024 268648 318030 268660
rect 447134 268648 447140 268660
rect 318024 268620 447140 268648
rect 318024 268608 318030 268620
rect 447134 268608 447140 268620
rect 447192 268608 447198 268660
rect 136634 268540 136640 268592
rect 136692 268580 136698 268592
rect 271046 268580 271052 268592
rect 136692 268552 271052 268580
rect 136692 268540 136698 268552
rect 271046 268540 271052 268552
rect 271104 268540 271110 268592
rect 319346 268540 319352 268592
rect 319404 268580 319410 268592
rect 455414 268580 455420 268592
rect 319404 268552 455420 268580
rect 319404 268540 319410 268552
rect 455414 268540 455420 268552
rect 455472 268540 455478 268592
rect 115934 268472 115940 268524
rect 115992 268512 115998 268524
rect 268102 268512 268108 268524
rect 115992 268484 268108 268512
rect 115992 268472 115998 268484
rect 268102 268472 268108 268484
rect 268160 268472 268166 268524
rect 325878 268472 325884 268524
rect 325936 268512 325942 268524
rect 502334 268512 502340 268524
rect 325936 268484 502340 268512
rect 325936 268472 325942 268484
rect 502334 268472 502340 268484
rect 502392 268472 502398 268524
rect 95234 268404 95240 268456
rect 95292 268444 95298 268456
rect 265526 268444 265532 268456
rect 95292 268416 265532 268444
rect 95292 268404 95298 268416
rect 265526 268404 265532 268416
rect 265584 268404 265590 268456
rect 325970 268404 325976 268456
rect 326028 268444 326034 268456
rect 503714 268444 503720 268456
rect 326028 268416 503720 268444
rect 326028 268404 326034 268416
rect 503714 268404 503720 268416
rect 503772 268404 503778 268456
rect 92474 268336 92480 268388
rect 92532 268376 92538 268388
rect 265434 268376 265440 268388
rect 92532 268348 265440 268376
rect 92532 268336 92538 268348
rect 265434 268336 265440 268348
rect 265492 268336 265498 268388
rect 335906 268336 335912 268388
rect 335964 268376 335970 268388
rect 565814 268376 565820 268388
rect 335964 268348 565820 268376
rect 335964 268336 335970 268348
rect 565814 268336 565820 268348
rect 565872 268336 565878 268388
rect 3510 267656 3516 267708
rect 3568 267696 3574 267708
rect 225598 267696 225604 267708
rect 3568 267668 225604 267696
rect 3568 267656 3574 267668
rect 225598 267656 225604 267668
rect 225656 267656 225662 267708
rect 309318 267248 309324 267300
rect 309376 267288 309382 267300
rect 390554 267288 390560 267300
rect 309376 267260 390560 267288
rect 309376 267248 309382 267260
rect 390554 267248 390560 267260
rect 390612 267248 390618 267300
rect 187694 267180 187700 267232
rect 187752 267220 187758 267232
rect 279234 267220 279240 267232
rect 187752 267192 279240 267220
rect 187752 267180 187758 267192
rect 279234 267180 279240 267192
rect 279292 267180 279298 267232
rect 309410 267180 309416 267232
rect 309468 267220 309474 267232
rect 394694 267220 394700 267232
rect 309468 267192 394700 267220
rect 309468 267180 309474 267192
rect 394694 267180 394700 267192
rect 394752 267180 394758 267232
rect 122834 267112 122840 267164
rect 122892 267152 122898 267164
rect 269206 267152 269212 267164
rect 122892 267124 269212 267152
rect 122892 267112 122898 267124
rect 269206 267112 269212 267124
rect 269264 267112 269270 267164
rect 314838 267112 314844 267164
rect 314896 267152 314902 267164
rect 427814 267152 427820 267164
rect 314896 267124 427820 267152
rect 314896 267112 314902 267124
rect 427814 267112 427820 267124
rect 427872 267112 427878 267164
rect 114554 267044 114560 267096
rect 114612 267084 114618 267096
rect 268010 267084 268016 267096
rect 114612 267056 268016 267084
rect 114612 267044 114618 267056
rect 268010 267044 268016 267056
rect 268068 267044 268074 267096
rect 319254 267044 319260 267096
rect 319312 267084 319318 267096
rect 451274 267084 451280 267096
rect 319312 267056 451280 267084
rect 319312 267044 319318 267056
rect 451274 267044 451280 267056
rect 451332 267044 451338 267096
rect 63494 266976 63500 267028
rect 63552 267016 63558 267028
rect 260098 267016 260104 267028
rect 63552 266988 260104 267016
rect 63552 266976 63558 266988
rect 260098 266976 260104 266988
rect 260156 266976 260162 267028
rect 327350 266976 327356 267028
rect 327408 267016 327414 267028
rect 514018 267016 514024 267028
rect 327408 266988 514024 267016
rect 327408 266976 327414 266988
rect 514018 266976 514024 266988
rect 514076 266976 514082 267028
rect 162854 265888 162860 265940
rect 162912 265928 162918 265940
rect 274818 265928 274824 265940
rect 162912 265900 274824 265928
rect 162912 265888 162918 265900
rect 274818 265888 274824 265900
rect 274876 265888 274882 265940
rect 307938 265888 307944 265940
rect 307996 265928 308002 265940
rect 383654 265928 383660 265940
rect 307996 265900 383660 265928
rect 307996 265888 308002 265900
rect 383654 265888 383660 265900
rect 383712 265888 383718 265940
rect 138014 265820 138020 265872
rect 138072 265860 138078 265872
rect 272058 265860 272064 265872
rect 138072 265832 272064 265860
rect 138072 265820 138078 265832
rect 272058 265820 272064 265832
rect 272116 265820 272122 265872
rect 309226 265820 309232 265872
rect 309284 265860 309290 265872
rect 387794 265860 387800 265872
rect 309284 265832 387800 265860
rect 309284 265820 309290 265832
rect 387794 265820 387800 265832
rect 387852 265820 387858 265872
rect 70394 265752 70400 265804
rect 70452 265792 70458 265804
rect 261110 265792 261116 265804
rect 70452 265764 261116 265792
rect 70452 265752 70458 265764
rect 261110 265752 261116 265764
rect 261168 265752 261174 265804
rect 311986 265752 311992 265804
rect 312044 265792 312050 265804
rect 405734 265792 405740 265804
rect 312044 265764 405740 265792
rect 312044 265752 312050 265764
rect 405734 265752 405740 265764
rect 405792 265752 405798 265804
rect 60734 265684 60740 265736
rect 60792 265724 60798 265736
rect 260006 265724 260012 265736
rect 60792 265696 260012 265724
rect 60792 265684 60798 265696
rect 260006 265684 260012 265696
rect 260064 265684 260070 265736
rect 316126 265684 316132 265736
rect 316184 265724 316190 265736
rect 438854 265724 438860 265736
rect 316184 265696 438860 265724
rect 316184 265684 316190 265696
rect 438854 265684 438860 265696
rect 438912 265684 438918 265736
rect 40034 265616 40040 265668
rect 40092 265656 40098 265668
rect 257062 265656 257068 265668
rect 40092 265628 257068 265656
rect 40092 265616 40098 265628
rect 257062 265616 257068 265628
rect 257120 265616 257126 265668
rect 330018 265616 330024 265668
rect 330076 265656 330082 265668
rect 531406 265656 531412 265668
rect 330076 265628 531412 265656
rect 330076 265616 330082 265628
rect 531406 265616 531412 265628
rect 531464 265616 531470 265668
rect 208394 264596 208400 264648
rect 208452 264636 208458 264648
rect 281810 264636 281816 264648
rect 208452 264608 281816 264636
rect 208452 264596 208458 264608
rect 281810 264596 281816 264608
rect 281868 264596 281874 264648
rect 204254 264528 204260 264580
rect 204312 264568 204318 264580
rect 281902 264568 281908 264580
rect 204312 264540 281908 264568
rect 204312 264528 204318 264540
rect 281902 264528 281908 264540
rect 281960 264528 281966 264580
rect 306558 264528 306564 264580
rect 306616 264568 306622 264580
rect 376754 264568 376760 264580
rect 306616 264540 376760 264568
rect 306616 264528 306622 264540
rect 376754 264528 376760 264540
rect 376812 264528 376818 264580
rect 174538 264460 174544 264512
rect 174596 264500 174602 264512
rect 276566 264500 276572 264512
rect 174596 264472 276572 264500
rect 174596 264460 174602 264472
rect 276566 264460 276572 264472
rect 276624 264460 276630 264512
rect 307846 264460 307852 264512
rect 307904 264500 307910 264512
rect 380894 264500 380900 264512
rect 307904 264472 380900 264500
rect 307904 264460 307910 264472
rect 380894 264460 380900 264472
rect 380952 264460 380958 264512
rect 144914 264392 144920 264444
rect 144972 264432 144978 264444
rect 271966 264432 271972 264444
rect 144972 264404 271972 264432
rect 144972 264392 144978 264404
rect 271966 264392 271972 264404
rect 272024 264392 272030 264444
rect 317874 264392 317880 264444
rect 317932 264432 317938 264444
rect 448514 264432 448520 264444
rect 317932 264404 448520 264432
rect 317932 264392 317938 264404
rect 448514 264392 448520 264404
rect 448572 264392 448578 264444
rect 100754 264324 100760 264376
rect 100812 264364 100818 264376
rect 265342 264364 265348 264376
rect 100812 264336 265348 264364
rect 100812 264324 100818 264336
rect 265342 264324 265348 264336
rect 265400 264324 265406 264376
rect 325786 264324 325792 264376
rect 325844 264364 325850 264376
rect 499574 264364 499580 264376
rect 325844 264336 499580 264364
rect 325844 264324 325850 264336
rect 499574 264324 499580 264336
rect 499632 264324 499638 264376
rect 74534 264256 74540 264308
rect 74592 264296 74598 264308
rect 262766 264296 262772 264308
rect 74592 264268 262772 264296
rect 74592 264256 74598 264268
rect 262766 264256 262772 264268
rect 262824 264256 262830 264308
rect 328914 264256 328920 264308
rect 328972 264296 328978 264308
rect 521654 264296 521660 264308
rect 328972 264268 521660 264296
rect 328972 264256 328978 264268
rect 521654 264256 521660 264268
rect 521712 264256 521718 264308
rect 46198 264188 46204 264240
rect 46256 264228 46262 264240
rect 256970 264228 256976 264240
rect 46256 264200 256976 264228
rect 46256 264188 46262 264200
rect 256970 264188 256976 264200
rect 257028 264188 257034 264240
rect 331490 264188 331496 264240
rect 331548 264228 331554 264240
rect 539594 264228 539600 264240
rect 331548 264200 539600 264228
rect 331548 264188 331554 264200
rect 539594 264188 539600 264200
rect 539652 264188 539658 264240
rect 201586 263168 201592 263220
rect 201644 263208 201650 263220
rect 280430 263208 280436 263220
rect 201644 263180 280436 263208
rect 201644 263168 201650 263180
rect 280430 263168 280436 263180
rect 280488 263168 280494 263220
rect 154574 263100 154580 263152
rect 154632 263140 154638 263152
rect 273898 263140 273904 263152
rect 154632 263112 273904 263140
rect 154632 263100 154638 263112
rect 273898 263100 273904 263112
rect 273956 263100 273962 263152
rect 306374 263100 306380 263152
rect 306432 263140 306438 263152
rect 374086 263140 374092 263152
rect 306432 263112 374092 263140
rect 306432 263100 306438 263112
rect 374086 263100 374092 263112
rect 374144 263100 374150 263152
rect 113174 263032 113180 263084
rect 113232 263072 113238 263084
rect 267918 263072 267924 263084
rect 113232 263044 267924 263072
rect 113232 263032 113238 263044
rect 267918 263032 267924 263044
rect 267976 263032 267982 263084
rect 317690 263032 317696 263084
rect 317748 263072 317754 263084
rect 441614 263072 441620 263084
rect 317748 263044 441620 263072
rect 317748 263032 317754 263044
rect 441614 263032 441620 263044
rect 441672 263032 441678 263084
rect 104894 262964 104900 263016
rect 104952 263004 104958 263016
rect 266538 263004 266544 263016
rect 104952 262976 266544 263004
rect 104952 262964 104958 262976
rect 266538 262964 266544 262976
rect 266596 262964 266602 263016
rect 317782 262964 317788 263016
rect 317840 263004 317846 263016
rect 444374 263004 444380 263016
rect 317840 262976 444380 263004
rect 317840 262964 317846 262976
rect 444374 262964 444380 262976
rect 444432 262964 444438 263016
rect 52454 262896 52460 262948
rect 52512 262936 52518 262948
rect 251818 262936 251824 262948
rect 52512 262908 251824 262936
rect 52512 262896 52518 262908
rect 251818 262896 251824 262908
rect 251876 262896 251882 262948
rect 320542 262896 320548 262948
rect 320600 262936 320606 262948
rect 466454 262936 466460 262948
rect 320600 262908 466460 262936
rect 320600 262896 320606 262908
rect 466454 262896 466460 262908
rect 466512 262896 466518 262948
rect 16574 262828 16580 262880
rect 16632 262868 16638 262880
rect 252738 262868 252744 262880
rect 16632 262840 252744 262868
rect 16632 262828 16638 262840
rect 252738 262828 252744 262840
rect 252796 262828 252802 262880
rect 336918 262828 336924 262880
rect 336976 262868 336982 262880
rect 578234 262868 578240 262880
rect 336976 262840 578240 262868
rect 336976 262828 336982 262840
rect 578234 262828 578240 262840
rect 578292 262828 578298 262880
rect 197354 261876 197360 261928
rect 197412 261916 197418 261928
rect 280246 261916 280252 261928
rect 197412 261888 280252 261916
rect 197412 261876 197418 261888
rect 280246 261876 280252 261888
rect 280304 261876 280310 261928
rect 193214 261808 193220 261860
rect 193272 261848 193278 261860
rect 280338 261848 280344 261860
rect 193272 261820 280344 261848
rect 193272 261808 193278 261820
rect 280338 261808 280344 261820
rect 280396 261808 280402 261860
rect 180794 261740 180800 261792
rect 180852 261780 180858 261792
rect 277762 261780 277768 261792
rect 180852 261752 277768 261780
rect 180852 261740 180858 261752
rect 277762 261740 277768 261752
rect 277820 261740 277826 261792
rect 97994 261672 98000 261724
rect 98052 261712 98058 261724
rect 265250 261712 265256 261724
rect 98052 261684 265256 261712
rect 98052 261672 98058 261684
rect 265250 261672 265256 261684
rect 265308 261672 265314 261724
rect 320450 261672 320456 261724
rect 320508 261712 320514 261724
rect 462314 261712 462320 261724
rect 320508 261684 462320 261712
rect 320508 261672 320514 261684
rect 462314 261672 462320 261684
rect 462372 261672 462378 261724
rect 85666 261604 85672 261656
rect 85724 261644 85730 261656
rect 263870 261644 263876 261656
rect 85724 261616 263876 261644
rect 85724 261604 85730 261616
rect 263870 261604 263876 261616
rect 263928 261604 263934 261656
rect 320358 261604 320364 261656
rect 320416 261644 320422 261656
rect 463694 261644 463700 261656
rect 320416 261616 463700 261644
rect 320416 261604 320422 261616
rect 463694 261604 463700 261616
rect 463752 261604 463758 261656
rect 49694 261536 49700 261588
rect 49752 261576 49758 261588
rect 258534 261576 258540 261588
rect 49752 261548 258540 261576
rect 49752 261536 49758 261548
rect 258534 261536 258540 261548
rect 258592 261536 258598 261588
rect 321646 261536 321652 261588
rect 321704 261576 321710 261588
rect 474734 261576 474740 261588
rect 321704 261548 474740 261576
rect 321704 261536 321710 261548
rect 474734 261536 474740 261548
rect 474792 261536 474798 261588
rect 25590 261468 25596 261520
rect 25648 261508 25654 261520
rect 252646 261508 252652 261520
rect 25648 261480 252652 261508
rect 25648 261468 25654 261480
rect 252646 261468 252652 261480
rect 252704 261468 252710 261520
rect 324498 261468 324504 261520
rect 324556 261508 324562 261520
rect 496078 261508 496084 261520
rect 324556 261480 496084 261508
rect 324556 261468 324562 261480
rect 496078 261468 496084 261480
rect 496136 261468 496142 261520
rect 190454 260516 190460 260568
rect 190512 260556 190518 260568
rect 279142 260556 279148 260568
rect 190512 260528 279148 260556
rect 190512 260516 190518 260528
rect 279142 260516 279148 260528
rect 279200 260516 279206 260568
rect 186314 260448 186320 260500
rect 186372 260488 186378 260500
rect 279050 260488 279056 260500
rect 186372 260460 279056 260488
rect 186372 260448 186378 260460
rect 279050 260448 279056 260460
rect 279108 260448 279114 260500
rect 217594 260380 217600 260432
rect 217652 260420 217658 260432
rect 338114 260420 338120 260432
rect 217652 260392 338120 260420
rect 217652 260380 217658 260392
rect 338114 260380 338120 260392
rect 338172 260380 338178 260432
rect 110506 260312 110512 260364
rect 110564 260352 110570 260364
rect 250622 260352 250628 260364
rect 110564 260324 250628 260352
rect 110564 260312 110570 260324
rect 250622 260312 250628 260324
rect 250680 260312 250686 260364
rect 329926 260312 329932 260364
rect 329984 260352 329990 260364
rect 532694 260352 532700 260364
rect 329984 260324 532700 260352
rect 329984 260312 329990 260324
rect 532694 260312 532700 260324
rect 532752 260312 532758 260364
rect 27614 260244 27620 260296
rect 27672 260284 27678 260296
rect 254302 260284 254308 260296
rect 27672 260256 254308 260284
rect 27672 260244 27678 260256
rect 254302 260244 254308 260256
rect 254360 260244 254366 260296
rect 331306 260244 331312 260296
rect 331364 260284 331370 260296
rect 536834 260284 536840 260296
rect 331364 260256 536840 260284
rect 331364 260244 331370 260256
rect 536834 260244 536840 260256
rect 536892 260244 536898 260296
rect 9674 260176 9680 260228
rect 9732 260216 9738 260228
rect 253198 260216 253204 260228
rect 9732 260188 253204 260216
rect 9732 260176 9738 260188
rect 253198 260176 253204 260188
rect 253256 260176 253262 260228
rect 331398 260176 331404 260228
rect 331456 260216 331462 260228
rect 539686 260216 539692 260228
rect 331456 260188 539692 260216
rect 331456 260176 331462 260188
rect 539686 260176 539692 260188
rect 539744 260176 539750 260228
rect 7558 260108 7564 260160
rect 7616 260148 7622 260160
rect 251358 260148 251364 260160
rect 7616 260120 251364 260148
rect 7616 260108 7622 260120
rect 251358 260108 251364 260120
rect 251416 260108 251422 260160
rect 335814 260108 335820 260160
rect 335872 260148 335878 260160
rect 568574 260148 568580 260160
rect 335872 260120 568580 260148
rect 335872 260108 335878 260120
rect 568574 260108 568580 260120
rect 568632 260108 568638 260160
rect 353938 259360 353944 259412
rect 353996 259400 354002 259412
rect 579798 259400 579804 259412
rect 353996 259372 579804 259400
rect 353996 259360 354002 259372
rect 579798 259360 579804 259372
rect 579856 259360 579862 259412
rect 183554 258884 183560 258936
rect 183612 258924 183618 258936
rect 272518 258924 272524 258936
rect 183612 258896 272524 258924
rect 183612 258884 183618 258896
rect 272518 258884 272524 258896
rect 272576 258884 272582 258936
rect 179414 258816 179420 258868
rect 179472 258856 179478 258868
rect 277670 258856 277676 258868
rect 179472 258828 277676 258856
rect 179472 258816 179478 258828
rect 277670 258816 277676 258828
rect 277728 258816 277734 258868
rect 176654 258748 176660 258800
rect 176712 258788 176718 258800
rect 277578 258788 277584 258800
rect 176712 258760 277584 258788
rect 176712 258748 176718 258760
rect 277578 258748 277584 258760
rect 277636 258748 277642 258800
rect 331950 258748 331956 258800
rect 332008 258788 332014 258800
rect 525794 258788 525800 258800
rect 332008 258760 525800 258788
rect 332008 258748 332014 258760
rect 525794 258748 525800 258760
rect 525852 258748 525858 258800
rect 93854 258680 93860 258732
rect 93912 258720 93918 258732
rect 265158 258720 265164 258732
rect 93912 258692 265164 258720
rect 93912 258680 93918 258692
rect 265158 258680 265164 258692
rect 265216 258680 265222 258732
rect 329834 258680 329840 258732
rect 329892 258720 329898 258732
rect 529934 258720 529940 258732
rect 329892 258692 529940 258720
rect 329892 258680 329898 258692
rect 529934 258680 529940 258692
rect 529992 258680 529998 258732
rect 209866 257660 209872 257712
rect 209924 257700 209930 257712
rect 281718 257700 281724 257712
rect 209924 257672 281724 257700
rect 209924 257660 209930 257672
rect 281718 257660 281724 257672
rect 281776 257660 281782 257712
rect 96614 257592 96620 257644
rect 96672 257632 96678 257644
rect 265066 257632 265072 257644
rect 96672 257604 265072 257632
rect 96672 257592 96678 257604
rect 265066 257592 265072 257604
rect 265124 257592 265130 257644
rect 42794 257524 42800 257576
rect 42852 257564 42858 257576
rect 256786 257564 256792 257576
rect 42852 257536 256792 257564
rect 42852 257524 42858 257536
rect 256786 257524 256792 257536
rect 256844 257524 256850 257576
rect 38654 257456 38660 257508
rect 38712 257496 38718 257508
rect 256878 257496 256884 257508
rect 38712 257468 256884 257496
rect 38712 257456 38718 257468
rect 256878 257456 256884 257468
rect 256936 257456 256942 257508
rect 329190 257456 329196 257508
rect 329248 257496 329254 257508
rect 514846 257496 514852 257508
rect 329248 257468 514852 257496
rect 329248 257456 329254 257468
rect 514846 257456 514852 257468
rect 514904 257456 514910 257508
rect 35894 257388 35900 257440
rect 35952 257428 35958 257440
rect 255682 257428 255688 257440
rect 35952 257400 255688 257428
rect 35952 257388 35958 257400
rect 255682 257388 255688 257400
rect 255740 257388 255746 257440
rect 328822 257388 328828 257440
rect 328880 257428 328886 257440
rect 523034 257428 523040 257440
rect 328880 257400 523040 257428
rect 328880 257388 328886 257400
rect 523034 257388 523040 257400
rect 523092 257388 523098 257440
rect 22094 257320 22100 257372
rect 22152 257360 22158 257372
rect 254210 257360 254216 257372
rect 22152 257332 254216 257360
rect 22152 257320 22158 257332
rect 254210 257320 254216 257332
rect 254268 257320 254274 257372
rect 335722 257320 335728 257372
rect 335780 257360 335786 257372
rect 564434 257360 564440 257372
rect 335780 257332 564440 257360
rect 335780 257320 335786 257332
rect 564434 257320 564440 257332
rect 564492 257320 564498 257372
rect 207014 256368 207020 256420
rect 207072 256408 207078 256420
rect 281626 256408 281632 256420
rect 207072 256380 281632 256408
rect 207072 256368 207078 256380
rect 281626 256368 281632 256380
rect 281684 256368 281690 256420
rect 313366 256368 313372 256420
rect 313424 256408 313430 256420
rect 422294 256408 422300 256420
rect 313424 256380 422300 256408
rect 313424 256368 313430 256380
rect 422294 256368 422300 256380
rect 422352 256368 422358 256420
rect 217134 256300 217140 256352
rect 217192 256340 217198 256352
rect 342898 256340 342904 256352
rect 217192 256312 342904 256340
rect 217192 256300 217198 256312
rect 342898 256300 342904 256312
rect 342956 256300 342962 256352
rect 80054 256232 80060 256284
rect 80112 256272 80118 256284
rect 262674 256272 262680 256284
rect 80112 256244 262680 256272
rect 80112 256232 80118 256244
rect 262674 256232 262680 256244
rect 262732 256232 262738 256284
rect 314746 256232 314752 256284
rect 314804 256272 314810 256284
rect 428458 256272 428464 256284
rect 314804 256244 428464 256272
rect 314804 256232 314810 256244
rect 428458 256232 428464 256244
rect 428516 256232 428522 256284
rect 41414 256164 41420 256216
rect 41472 256204 41478 256216
rect 256694 256204 256700 256216
rect 41472 256176 256700 256204
rect 41472 256164 41478 256176
rect 256694 256164 256700 256176
rect 256752 256164 256758 256216
rect 316034 256164 316040 256216
rect 316092 256204 316098 256216
rect 436094 256204 436100 256216
rect 316092 256176 436100 256204
rect 316092 256164 316098 256176
rect 436094 256164 436100 256176
rect 436152 256164 436158 256216
rect 34514 256096 34520 256148
rect 34572 256136 34578 256148
rect 255406 256136 255412 256148
rect 34572 256108 255412 256136
rect 34572 256096 34578 256108
rect 255406 256096 255412 256108
rect 255464 256096 255470 256148
rect 317598 256096 317604 256148
rect 317656 256136 317662 256148
rect 442994 256136 443000 256148
rect 317656 256108 443000 256136
rect 317656 256096 317662 256108
rect 442994 256096 443000 256108
rect 443052 256096 443058 256148
rect 30374 256028 30380 256080
rect 30432 256068 30438 256080
rect 255590 256068 255596 256080
rect 30432 256040 255596 256068
rect 30432 256028 30438 256040
rect 255590 256028 255596 256040
rect 255648 256028 255654 256080
rect 325694 256028 325700 256080
rect 325752 256068 325758 256080
rect 505094 256068 505100 256080
rect 325752 256040 505100 256068
rect 325752 256028 325758 256040
rect 505094 256028 505100 256040
rect 505152 256028 505158 256080
rect 27706 255960 27712 256012
rect 27764 256000 27770 256012
rect 255498 256000 255504 256012
rect 27764 255972 255504 256000
rect 27764 255960 27770 255972
rect 255498 255960 255504 255972
rect 255556 255960 255562 256012
rect 327258 255960 327264 256012
rect 327316 256000 327322 256012
rect 511994 256000 512000 256012
rect 327316 255972 512000 256000
rect 327316 255960 327322 255972
rect 511994 255960 512000 255972
rect 512052 255960 512058 256012
rect 3510 255144 3516 255196
rect 3568 255184 3574 255196
rect 8938 255184 8944 255196
rect 3568 255156 8944 255184
rect 3568 255144 3574 255156
rect 8938 255144 8944 255156
rect 8996 255144 9002 255196
rect 202874 254940 202880 254992
rect 202932 254980 202938 254992
rect 281534 254980 281540 254992
rect 202932 254952 281540 254980
rect 202932 254940 202938 254952
rect 281534 254940 281540 254952
rect 281592 254940 281598 254992
rect 200114 254872 200120 254924
rect 200172 254912 200178 254924
rect 280614 254912 280620 254924
rect 200172 254884 280620 254912
rect 200172 254872 200178 254884
rect 280614 254872 280620 254884
rect 280672 254872 280678 254924
rect 307754 254872 307760 254924
rect 307812 254912 307818 254924
rect 379514 254912 379520 254924
rect 307812 254884 379520 254912
rect 307812 254872 307818 254884
rect 379514 254872 379520 254884
rect 379572 254872 379578 254924
rect 102226 254804 102232 254856
rect 102284 254844 102290 254856
rect 266446 254844 266452 254856
rect 102284 254816 266452 254844
rect 102284 254804 102290 254816
rect 266446 254804 266452 254816
rect 266504 254804 266510 254856
rect 309134 254804 309140 254856
rect 309192 254844 309198 254856
rect 390646 254844 390652 254856
rect 309192 254816 390652 254844
rect 309192 254804 309198 254816
rect 390646 254804 390652 254816
rect 390704 254804 390710 254856
rect 93946 254736 93952 254788
rect 94004 254776 94010 254788
rect 264974 254776 264980 254788
rect 94004 254748 264980 254776
rect 94004 254736 94010 254748
rect 264974 254736 264980 254748
rect 265032 254736 265038 254788
rect 320266 254736 320272 254788
rect 320324 254776 320330 254788
rect 460934 254776 460940 254788
rect 320324 254748 460940 254776
rect 320324 254736 320330 254748
rect 460934 254736 460940 254748
rect 460992 254736 460998 254788
rect 91094 254668 91100 254720
rect 91152 254708 91158 254720
rect 263778 254708 263784 254720
rect 91152 254680 263784 254708
rect 91152 254668 91158 254680
rect 263778 254668 263784 254680
rect 263836 254668 263842 254720
rect 329098 254668 329104 254720
rect 329156 254708 329162 254720
rect 498286 254708 498292 254720
rect 329156 254680 498292 254708
rect 329156 254668 329162 254680
rect 498286 254668 498292 254680
rect 498344 254668 498350 254720
rect 77294 254600 77300 254652
rect 77352 254640 77358 254652
rect 262582 254640 262588 254652
rect 77352 254612 262588 254640
rect 77352 254600 77358 254612
rect 262582 254600 262588 254612
rect 262640 254600 262646 254652
rect 334342 254600 334348 254652
rect 334400 254640 334406 254652
rect 556246 254640 556252 254652
rect 334400 254612 556252 254640
rect 334400 254600 334406 254612
rect 556246 254600 556252 254612
rect 556304 254600 556310 254652
rect 73154 254532 73160 254584
rect 73212 254572 73218 254584
rect 261018 254572 261024 254584
rect 73212 254544 261024 254572
rect 73212 254532 73218 254544
rect 261018 254532 261024 254544
rect 261076 254532 261082 254584
rect 334250 254532 334256 254584
rect 334308 254572 334314 254584
rect 560294 254572 560300 254584
rect 334308 254544 560300 254572
rect 334308 254532 334314 254544
rect 560294 254532 560300 254544
rect 560352 254532 560358 254584
rect 193306 253648 193312 253700
rect 193364 253688 193370 253700
rect 278958 253688 278964 253700
rect 193364 253660 278964 253688
rect 193364 253648 193370 253660
rect 278958 253648 278964 253660
rect 279016 253648 279022 253700
rect 217042 253580 217048 253632
rect 217100 253620 217106 253632
rect 340966 253620 340972 253632
rect 217100 253592 340972 253620
rect 217100 253580 217106 253592
rect 340966 253580 340972 253592
rect 341024 253580 341030 253632
rect 121454 253512 121460 253564
rect 121512 253552 121518 253564
rect 269574 253552 269580 253564
rect 121512 253524 269580 253552
rect 121512 253512 121518 253524
rect 269574 253512 269580 253524
rect 269632 253512 269638 253564
rect 319162 253512 319168 253564
rect 319220 253552 319226 253564
rect 456794 253552 456800 253564
rect 319220 253524 456800 253552
rect 319220 253512 319226 253524
rect 456794 253512 456800 253524
rect 456852 253512 456858 253564
rect 118694 253444 118700 253496
rect 118752 253484 118758 253496
rect 267826 253484 267832 253496
rect 118752 253456 267832 253484
rect 118752 253444 118758 253456
rect 267826 253444 267832 253456
rect 267884 253444 267890 253496
rect 323210 253444 323216 253496
rect 323268 253484 323274 253496
rect 485774 253484 485780 253496
rect 323268 253456 485780 253484
rect 323268 253444 323274 253456
rect 485774 253444 485780 253456
rect 485832 253444 485838 253496
rect 82814 253376 82820 253428
rect 82872 253416 82878 253428
rect 262490 253416 262496 253428
rect 82872 253388 262496 253416
rect 82872 253376 82878 253388
rect 262490 253376 262496 253388
rect 262548 253376 262554 253428
rect 324406 253376 324412 253428
rect 324464 253416 324470 253428
rect 489914 253416 489920 253428
rect 324464 253388 489920 253416
rect 324464 253376 324470 253388
rect 489914 253376 489920 253388
rect 489972 253376 489978 253428
rect 69014 253308 69020 253360
rect 69072 253348 69078 253360
rect 260926 253348 260932 253360
rect 69072 253320 260932 253348
rect 69072 253308 69078 253320
rect 260926 253308 260932 253320
rect 260984 253308 260990 253360
rect 327166 253308 327172 253360
rect 327224 253348 327230 253360
rect 507854 253348 507860 253360
rect 327224 253320 507860 253348
rect 327224 253308 327230 253320
rect 507854 253308 507860 253320
rect 507912 253308 507918 253360
rect 62114 253240 62120 253292
rect 62172 253280 62178 253292
rect 259914 253280 259920 253292
rect 62172 253252 259920 253280
rect 62172 253240 62178 253252
rect 259914 253240 259920 253252
rect 259972 253240 259978 253292
rect 331214 253240 331220 253292
rect 331272 253280 331278 253292
rect 535454 253280 535460 253292
rect 331272 253252 535460 253280
rect 331272 253240 331278 253252
rect 535454 253240 535460 253252
rect 535512 253240 535518 253292
rect 23474 253172 23480 253224
rect 23532 253212 23538 253224
rect 250530 253212 250536 253224
rect 23532 253184 250536 253212
rect 23532 253172 23538 253184
rect 250530 253172 250536 253184
rect 250588 253172 250594 253224
rect 335630 253172 335636 253224
rect 335688 253212 335694 253224
rect 561674 253212 561680 253224
rect 335688 253184 561680 253212
rect 335688 253172 335694 253184
rect 561674 253172 561680 253184
rect 561732 253172 561738 253224
rect 218514 252152 218520 252204
rect 218572 252192 218578 252204
rect 341426 252192 341432 252204
rect 218572 252164 341432 252192
rect 218572 252152 218578 252164
rect 341426 252152 341432 252164
rect 341484 252152 341490 252204
rect 86954 252084 86960 252136
rect 87012 252124 87018 252136
rect 263686 252124 263692 252136
rect 87012 252096 263692 252124
rect 87012 252084 87018 252096
rect 263686 252084 263692 252096
rect 263744 252084 263750 252136
rect 313274 252084 313280 252136
rect 313332 252124 313338 252136
rect 420914 252124 420920 252136
rect 313332 252096 420920 252124
rect 313332 252084 313338 252096
rect 420914 252084 420920 252096
rect 420972 252084 420978 252136
rect 78674 252016 78680 252068
rect 78732 252056 78738 252068
rect 262398 252056 262404 252068
rect 78732 252028 262404 252056
rect 78732 252016 78738 252028
rect 262398 252016 262404 252028
rect 262456 252016 262462 252068
rect 319070 252016 319076 252068
rect 319128 252056 319134 252068
rect 459554 252056 459560 252068
rect 319128 252028 459560 252056
rect 319128 252016 319134 252028
rect 459554 252016 459560 252028
rect 459612 252016 459618 252068
rect 26234 251948 26240 252000
rect 26292 251988 26298 252000
rect 254026 251988 254032 252000
rect 26292 251960 254032 251988
rect 26292 251948 26298 251960
rect 254026 251948 254032 251960
rect 254084 251948 254090 252000
rect 328730 251948 328736 252000
rect 328788 251988 328794 252000
rect 518894 251988 518900 252000
rect 328788 251960 518900 251988
rect 328788 251948 328794 251960
rect 518894 251948 518900 251960
rect 518952 251948 518958 252000
rect 19334 251880 19340 251932
rect 19392 251920 19398 251932
rect 254118 251920 254124 251932
rect 19392 251892 254124 251920
rect 19392 251880 19398 251892
rect 254118 251880 254124 251892
rect 254176 251880 254182 251932
rect 332686 251880 332692 251932
rect 332744 251920 332750 251932
rect 549254 251920 549260 251932
rect 332744 251892 549260 251920
rect 332744 251880 332750 251892
rect 549254 251880 549260 251892
rect 549312 251880 549318 251932
rect 8294 251812 8300 251864
rect 8352 251852 8358 251864
rect 251266 251852 251272 251864
rect 8352 251824 251272 251852
rect 8352 251812 8358 251824
rect 251266 251812 251272 251824
rect 251324 251812 251330 251864
rect 335538 251812 335544 251864
rect 335596 251852 335602 251864
rect 564526 251852 564532 251864
rect 335596 251824 564532 251852
rect 335596 251812 335602 251824
rect 564526 251812 564532 251824
rect 564584 251812 564590 251864
rect 301498 251132 301504 251184
rect 301556 251172 301562 251184
rect 363046 251172 363052 251184
rect 301556 251144 363052 251172
rect 301556 251132 301562 251144
rect 363046 251132 363052 251144
rect 363104 251132 363110 251184
rect 301314 251064 301320 251116
rect 301372 251104 301378 251116
rect 362954 251104 362960 251116
rect 301372 251076 362960 251104
rect 301372 251064 301378 251076
rect 362954 251064 362960 251076
rect 363012 251064 363018 251116
rect 301406 250996 301412 251048
rect 301464 251036 301470 251048
rect 363230 251036 363236 251048
rect 301464 251008 363236 251036
rect 301464 250996 301470 251008
rect 363230 250996 363236 251008
rect 363288 250996 363294 251048
rect 298278 250928 298284 250980
rect 298336 250968 298342 250980
rect 360654 250968 360660 250980
rect 298336 250940 360660 250968
rect 298336 250928 298342 250940
rect 360654 250928 360660 250940
rect 360712 250928 360718 250980
rect 300026 250860 300032 250912
rect 300084 250900 300090 250912
rect 363138 250900 363144 250912
rect 300084 250872 363144 250900
rect 300084 250860 300090 250872
rect 363138 250860 363144 250872
rect 363196 250860 363202 250912
rect 311894 250792 311900 250844
rect 311952 250832 311958 250844
rect 409874 250832 409880 250844
rect 311952 250804 409880 250832
rect 311952 250792 311958 250804
rect 409874 250792 409880 250804
rect 409932 250792 409938 250844
rect 142154 250724 142160 250776
rect 142212 250764 142218 250776
rect 272426 250764 272432 250776
rect 142212 250736 272432 250764
rect 142212 250724 142218 250736
rect 272426 250724 272432 250736
rect 272484 250724 272490 250776
rect 317506 250724 317512 250776
rect 317564 250764 317570 250776
rect 445754 250764 445760 250776
rect 317564 250736 445760 250764
rect 317564 250724 317570 250736
rect 445754 250724 445760 250736
rect 445812 250724 445818 250776
rect 77386 250656 77392 250708
rect 77444 250696 77450 250708
rect 262306 250696 262312 250708
rect 77444 250668 262312 250696
rect 77444 250656 77450 250668
rect 262306 250656 262312 250668
rect 262364 250656 262370 250708
rect 325050 250656 325056 250708
rect 325108 250696 325114 250708
rect 487154 250696 487160 250708
rect 325108 250668 487160 250696
rect 325108 250656 325114 250668
rect 487154 250656 487160 250668
rect 487212 250656 487218 250708
rect 75914 250588 75920 250640
rect 75972 250628 75978 250640
rect 262858 250628 262864 250640
rect 75972 250600 262864 250628
rect 75972 250588 75978 250600
rect 262858 250588 262864 250600
rect 262916 250588 262922 250640
rect 327810 250588 327816 250640
rect 327868 250628 327874 250640
rect 494054 250628 494060 250640
rect 327868 250600 494060 250628
rect 327868 250588 327874 250600
rect 494054 250588 494060 250600
rect 494112 250588 494118 250640
rect 55214 250520 55220 250572
rect 55272 250560 55278 250572
rect 259822 250560 259828 250572
rect 55272 250532 259828 250560
rect 55272 250520 55278 250532
rect 259822 250520 259828 250532
rect 259880 250520 259886 250572
rect 328638 250520 328644 250572
rect 328696 250560 328702 250572
rect 517514 250560 517520 250572
rect 328696 250532 517520 250560
rect 328696 250520 328702 250532
rect 517514 250520 517520 250532
rect 517572 250520 517578 250572
rect 11054 250452 11060 250504
rect 11112 250492 11118 250504
rect 246298 250492 246304 250504
rect 11112 250464 246304 250492
rect 11112 250452 11118 250464
rect 246298 250452 246304 250464
rect 246356 250452 246362 250504
rect 336826 250452 336832 250504
rect 336884 250492 336890 250504
rect 576854 250492 576860 250504
rect 336884 250464 576860 250492
rect 336884 250452 336890 250464
rect 576854 250452 576860 250464
rect 576912 250452 576918 250504
rect 189074 249364 189080 249416
rect 189132 249404 189138 249416
rect 278866 249404 278872 249416
rect 189132 249376 278872 249404
rect 189132 249364 189138 249376
rect 278866 249364 278872 249376
rect 278924 249364 278930 249416
rect 89714 249296 89720 249348
rect 89772 249336 89778 249348
rect 263594 249336 263600 249348
rect 89772 249308 263600 249336
rect 89772 249296 89778 249308
rect 263594 249296 263600 249308
rect 263652 249296 263658 249348
rect 318886 249296 318892 249348
rect 318944 249336 318950 249348
rect 452654 249336 452660 249348
rect 318944 249308 452660 249336
rect 318944 249296 318950 249308
rect 452654 249296 452660 249308
rect 452712 249296 452718 249348
rect 60826 249228 60832 249280
rect 60884 249268 60890 249280
rect 259638 249268 259644 249280
rect 60884 249240 259644 249268
rect 60884 249228 60890 249240
rect 259638 249228 259644 249240
rect 259696 249228 259702 249280
rect 318978 249228 318984 249280
rect 319036 249268 319042 249280
rect 456886 249268 456892 249280
rect 319036 249240 456892 249268
rect 319036 249228 319042 249240
rect 456886 249228 456892 249240
rect 456944 249228 456950 249280
rect 56594 249160 56600 249212
rect 56652 249200 56658 249212
rect 259730 249200 259736 249212
rect 56652 249172 259736 249200
rect 56652 249160 56658 249172
rect 259730 249160 259736 249172
rect 259788 249160 259794 249212
rect 324314 249160 324320 249212
rect 324372 249200 324378 249212
rect 490006 249200 490012 249212
rect 324372 249172 490012 249200
rect 324372 249160 324378 249172
rect 490006 249160 490012 249172
rect 490064 249160 490070 249212
rect 48314 249092 48320 249144
rect 48372 249132 48378 249144
rect 258442 249132 258448 249144
rect 48372 249104 258448 249132
rect 48372 249092 48378 249104
rect 258442 249092 258448 249104
rect 258500 249092 258506 249144
rect 328546 249092 328552 249144
rect 328604 249132 328610 249144
rect 523126 249132 523132 249144
rect 328604 249104 523132 249132
rect 328604 249092 328610 249104
rect 523126 249092 523132 249104
rect 523184 249092 523190 249144
rect 4154 249024 4160 249076
rect 4212 249064 4218 249076
rect 243538 249064 243544 249076
rect 4212 249036 243544 249064
rect 4212 249024 4218 249036
rect 243538 249024 243544 249036
rect 243596 249024 243602 249076
rect 335446 249024 335452 249076
rect 335504 249064 335510 249076
rect 567194 249064 567200 249076
rect 335504 249036 567200 249064
rect 335504 249024 335510 249036
rect 567194 249024 567200 249036
rect 567252 249024 567258 249076
rect 303798 248344 303804 248396
rect 303856 248384 303862 248396
rect 361942 248384 361948 248396
rect 303856 248356 361948 248384
rect 303856 248344 303862 248356
rect 361942 248344 361948 248356
rect 362000 248344 362006 248396
rect 302602 248276 302608 248328
rect 302660 248316 302666 248328
rect 361758 248316 361764 248328
rect 302660 248288 361764 248316
rect 302660 248276 302666 248288
rect 361758 248276 361764 248288
rect 361816 248276 361822 248328
rect 301222 248208 301228 248260
rect 301280 248248 301286 248260
rect 360562 248248 360568 248260
rect 301280 248220 360568 248248
rect 301280 248208 301286 248220
rect 360562 248208 360568 248220
rect 360620 248208 360626 248260
rect 204898 248140 204904 248192
rect 204956 248180 204962 248192
rect 258350 248180 258356 248192
rect 204956 248152 258356 248180
rect 204956 248140 204962 248152
rect 258350 248140 258356 248152
rect 258408 248140 258414 248192
rect 301038 248140 301044 248192
rect 301096 248180 301102 248192
rect 360470 248180 360476 248192
rect 301096 248152 360476 248180
rect 301096 248140 301102 248152
rect 360470 248140 360476 248152
rect 360528 248140 360534 248192
rect 185026 248072 185032 248124
rect 185084 248112 185090 248124
rect 279418 248112 279424 248124
rect 185084 248084 279424 248112
rect 185084 248072 185090 248084
rect 279418 248072 279424 248084
rect 279476 248072 279482 248124
rect 301130 248072 301136 248124
rect 301188 248112 301194 248124
rect 361666 248112 361672 248124
rect 301188 248084 361672 248112
rect 301188 248072 301194 248084
rect 361666 248072 361672 248084
rect 361724 248072 361730 248124
rect 182174 248004 182180 248056
rect 182232 248044 182238 248056
rect 277486 248044 277492 248056
rect 182232 248016 277492 248044
rect 182232 248004 182238 248016
rect 277486 248004 277492 248016
rect 277544 248004 277550 248056
rect 299842 248004 299848 248056
rect 299900 248044 299906 248056
rect 360746 248044 360752 248056
rect 299900 248016 360752 248044
rect 299900 248004 299906 248016
rect 360746 248004 360752 248016
rect 360804 248004 360810 248056
rect 173894 247936 173900 247988
rect 173952 247976 173958 247988
rect 276014 247976 276020 247988
rect 173952 247948 276020 247976
rect 173952 247936 173958 247948
rect 276014 247936 276020 247948
rect 276072 247936 276078 247988
rect 299934 247936 299940 247988
rect 299992 247976 299998 247988
rect 361850 247976 361856 247988
rect 299992 247948 361856 247976
rect 299992 247936 299998 247948
rect 361850 247936 361856 247948
rect 361908 247936 361914 247988
rect 155954 247868 155960 247920
rect 156012 247908 156018 247920
rect 273806 247908 273812 247920
rect 156012 247880 273812 247908
rect 156012 247868 156018 247880
rect 273806 247868 273812 247880
rect 273864 247868 273870 247920
rect 297082 247868 297088 247920
rect 297140 247908 297146 247920
rect 365806 247908 365812 247920
rect 297140 247880 365812 247908
rect 297140 247868 297146 247880
rect 365806 247868 365812 247880
rect 365864 247868 365870 247920
rect 67634 247800 67640 247852
rect 67692 247840 67698 247852
rect 261478 247840 261484 247852
rect 67692 247812 261484 247840
rect 67692 247800 67698 247812
rect 261478 247800 261484 247812
rect 261536 247800 261542 247852
rect 317414 247800 317420 247852
rect 317472 247840 317478 247852
rect 448606 247840 448612 247852
rect 317472 247812 448612 247840
rect 317472 247800 317478 247812
rect 448606 247800 448612 247812
rect 448664 247800 448670 247852
rect 57974 247732 57980 247784
rect 58032 247772 58038 247784
rect 259546 247772 259552 247784
rect 58032 247744 259552 247772
rect 58032 247732 58038 247744
rect 259546 247732 259552 247744
rect 259604 247732 259610 247784
rect 318794 247732 318800 247784
rect 318852 247772 318858 247784
rect 454034 247772 454040 247784
rect 318852 247744 454040 247772
rect 318852 247732 318858 247744
rect 454034 247732 454040 247744
rect 454092 247732 454098 247784
rect 20714 247664 20720 247716
rect 20772 247704 20778 247716
rect 254486 247704 254492 247716
rect 20772 247676 254492 247704
rect 20772 247664 20778 247676
rect 254486 247664 254492 247676
rect 254544 247664 254550 247716
rect 321554 247664 321560 247716
rect 321612 247704 321618 247716
rect 477494 247704 477500 247716
rect 321612 247676 477500 247704
rect 321612 247664 321618 247676
rect 477494 247664 477500 247676
rect 477552 247664 477558 247716
rect 299750 247596 299756 247648
rect 299808 247636 299814 247648
rect 357710 247636 357716 247648
rect 299808 247608 357716 247636
rect 299808 247596 299814 247608
rect 357710 247596 357716 247608
rect 357768 247596 357774 247648
rect 302510 247528 302516 247580
rect 302568 247568 302574 247580
rect 360378 247568 360384 247580
rect 302568 247540 360384 247568
rect 302568 247528 302574 247540
rect 360378 247528 360384 247540
rect 360436 247528 360442 247580
rect 347130 247460 347136 247512
rect 347188 247500 347194 247512
rect 369854 247500 369860 247512
rect 347188 247472 369860 247500
rect 347188 247460 347194 247472
rect 369854 247460 369860 247472
rect 369912 247460 369918 247512
rect 178034 246644 178040 246696
rect 178092 246684 178098 246696
rect 277946 246684 277952 246696
rect 178092 246656 277952 246684
rect 178092 246644 178098 246656
rect 277946 246644 277952 246656
rect 278004 246644 278010 246696
rect 118786 246576 118792 246628
rect 118844 246616 118850 246628
rect 268378 246616 268384 246628
rect 118844 246588 268384 246616
rect 118844 246576 118850 246588
rect 268378 246576 268384 246588
rect 268436 246576 268442 246628
rect 327074 246576 327080 246628
rect 327132 246616 327138 246628
rect 510614 246616 510620 246628
rect 327132 246588 510620 246616
rect 327132 246576 327138 246588
rect 510614 246576 510620 246588
rect 510672 246576 510678 246628
rect 59354 246508 59360 246560
rect 59412 246548 59418 246560
rect 259454 246548 259460 246560
rect 59412 246520 259460 246548
rect 59412 246508 59418 246520
rect 259454 246508 259460 246520
rect 259512 246508 259518 246560
rect 333974 246508 333980 246560
rect 334032 246548 334038 246560
rect 553394 246548 553400 246560
rect 334032 246520 553400 246548
rect 334032 246508 334038 246520
rect 553394 246508 553400 246520
rect 553452 246508 553458 246560
rect 53834 246440 53840 246492
rect 53892 246480 53898 246492
rect 258258 246480 258264 246492
rect 53892 246452 258264 246480
rect 53892 246440 53898 246452
rect 258258 246440 258264 246452
rect 258316 246440 258322 246492
rect 334066 246440 334072 246492
rect 334124 246480 334130 246492
rect 554774 246480 554780 246492
rect 334124 246452 554780 246480
rect 334124 246440 334130 246452
rect 554774 246440 554780 246452
rect 554832 246440 554838 246492
rect 51074 246372 51080 246424
rect 51132 246412 51138 246424
rect 258166 246412 258172 246424
rect 51132 246384 258172 246412
rect 51132 246372 51138 246384
rect 258166 246372 258172 246384
rect 258224 246372 258230 246424
rect 335354 246372 335360 246424
rect 335412 246412 335418 246424
rect 563054 246412 563060 246424
rect 335412 246384 563060 246412
rect 335412 246372 335418 246384
rect 563054 246372 563060 246384
rect 563112 246372 563118 246424
rect 6914 246304 6920 246356
rect 6972 246344 6978 246356
rect 251542 246344 251548 246356
rect 6972 246316 251548 246344
rect 6972 246304 6978 246316
rect 251542 246304 251548 246316
rect 251600 246304 251606 246356
rect 352558 246304 352564 246356
rect 352616 246344 352622 246356
rect 580166 246344 580172 246356
rect 352616 246316 580172 246344
rect 352616 246304 352622 246316
rect 580166 246304 580172 246316
rect 580224 246304 580230 246356
rect 300946 245556 300952 245608
rect 301004 245596 301010 245608
rect 359274 245596 359280 245608
rect 301004 245568 359280 245596
rect 301004 245556 301010 245568
rect 359274 245556 359280 245568
rect 359332 245556 359338 245608
rect 362494 245556 362500 245608
rect 362552 245596 362558 245608
rect 365714 245596 365720 245608
rect 362552 245568 365720 245596
rect 362552 245556 362558 245568
rect 365714 245556 365720 245568
rect 365772 245556 365778 245608
rect 299658 245488 299664 245540
rect 299716 245528 299722 245540
rect 358998 245528 359004 245540
rect 299716 245500 359004 245528
rect 299716 245488 299722 245500
rect 358998 245488 359004 245500
rect 359056 245488 359062 245540
rect 299474 245420 299480 245472
rect 299532 245460 299538 245472
rect 358906 245460 358912 245472
rect 299532 245432 358912 245460
rect 299532 245420 299538 245432
rect 358906 245420 358912 245432
rect 358964 245420 358970 245472
rect 299566 245352 299572 245404
rect 299624 245392 299630 245404
rect 359182 245392 359188 245404
rect 299624 245364 359188 245392
rect 299624 245352 299630 245364
rect 359182 245352 359188 245364
rect 359240 245352 359246 245404
rect 160186 245284 160192 245336
rect 160244 245324 160250 245336
rect 275186 245324 275192 245336
rect 160244 245296 275192 245324
rect 160244 245284 160250 245296
rect 275186 245284 275192 245296
rect 275244 245284 275250 245336
rect 296898 245284 296904 245336
rect 296956 245324 296962 245336
rect 357802 245324 357808 245336
rect 296956 245296 357808 245324
rect 296956 245284 296962 245296
rect 357802 245284 357808 245296
rect 357860 245284 357866 245336
rect 158714 245216 158720 245268
rect 158772 245256 158778 245268
rect 274726 245256 274732 245268
rect 158772 245228 274732 245256
rect 158772 245216 158778 245228
rect 274726 245216 274732 245228
rect 274784 245216 274790 245268
rect 296806 245216 296812 245268
rect 296864 245256 296870 245268
rect 359366 245256 359372 245268
rect 296864 245228 359372 245256
rect 296864 245216 296870 245228
rect 359366 245216 359372 245228
rect 359424 245216 359430 245268
rect 217226 245148 217232 245200
rect 217284 245188 217290 245200
rect 336734 245188 336740 245200
rect 217284 245160 336740 245188
rect 217284 245148 217290 245160
rect 336734 245148 336740 245160
rect 336792 245148 336798 245200
rect 349890 245148 349896 245200
rect 349948 245188 349954 245200
rect 362034 245188 362040 245200
rect 349948 245160 362040 245188
rect 349948 245148 349954 245160
rect 362034 245148 362040 245160
rect 362092 245148 362098 245200
rect 120074 245080 120080 245132
rect 120132 245120 120138 245132
rect 250438 245120 250444 245132
rect 120132 245092 250444 245120
rect 120132 245080 120138 245092
rect 250438 245080 250444 245092
rect 250496 245080 250502 245132
rect 295794 245080 295800 245132
rect 295852 245120 295858 245132
rect 363322 245120 363328 245132
rect 295852 245092 363328 245120
rect 295852 245080 295858 245092
rect 363322 245080 363328 245092
rect 363380 245080 363386 245132
rect 109034 245012 109040 245064
rect 109092 245052 109098 245064
rect 266998 245052 267004 245064
rect 109092 245024 267004 245052
rect 109092 245012 109098 245024
rect 266998 245012 267004 245024
rect 267056 245012 267062 245064
rect 298094 245012 298100 245064
rect 298152 245052 298158 245064
rect 368474 245052 368480 245064
rect 298152 245024 368480 245052
rect 298152 245012 298158 245024
rect 368474 245012 368480 245024
rect 368532 245012 368538 245064
rect 46934 244944 46940 244996
rect 46992 244984 46998 244996
rect 258626 244984 258632 244996
rect 46992 244956 258632 244984
rect 46992 244944 46998 244956
rect 258626 244944 258632 244956
rect 258684 244944 258690 244996
rect 296714 244944 296720 244996
rect 296772 244984 296778 244996
rect 367186 244984 367192 244996
rect 296772 244956 367192 244984
rect 296772 244944 296778 244956
rect 367186 244944 367192 244956
rect 367244 244944 367250 244996
rect 35986 244876 35992 244928
rect 36044 244916 36050 244928
rect 255958 244916 255964 244928
rect 36044 244888 255964 244916
rect 36044 244876 36050 244888
rect 255958 244876 255964 244888
rect 256016 244876 256022 244928
rect 314654 244876 314660 244928
rect 314712 244916 314718 244928
rect 432046 244916 432052 244928
rect 314712 244888 432052 244916
rect 314712 244876 314718 244888
rect 432046 244876 432052 244888
rect 432104 244876 432110 244928
rect 300854 244808 300860 244860
rect 300912 244848 300918 244860
rect 359090 244848 359096 244860
rect 300912 244820 359096 244848
rect 300912 244808 300918 244820
rect 359090 244808 359096 244820
rect 359148 244808 359154 244860
rect 302326 244740 302332 244792
rect 302384 244780 302390 244792
rect 357618 244780 357624 244792
rect 302384 244752 357624 244780
rect 302384 244740 302390 244752
rect 357618 244740 357624 244752
rect 357676 244740 357682 244792
rect 355410 244468 355416 244520
rect 355468 244508 355474 244520
rect 363414 244508 363420 244520
rect 355468 244480 363420 244508
rect 355468 244468 355474 244480
rect 363414 244468 363420 244480
rect 363472 244468 363478 244520
rect 218606 243720 218612 243772
rect 218664 243760 218670 243772
rect 293218 243760 293224 243772
rect 218664 243732 293224 243760
rect 218664 243720 218670 243732
rect 293218 243720 293224 243732
rect 293276 243720 293282 243772
rect 295702 243720 295708 243772
rect 295760 243760 295766 243772
rect 357894 243760 357900 243772
rect 295760 243732 357900 243760
rect 295760 243720 295766 243732
rect 357894 243720 357900 243732
rect 357952 243720 357958 243772
rect 219250 243652 219256 243704
rect 219308 243692 219314 243704
rect 293954 243692 293960 243704
rect 219308 243664 293960 243692
rect 219308 243652 219314 243664
rect 293954 243652 293960 243664
rect 294012 243652 294018 243704
rect 295610 243652 295616 243704
rect 295668 243692 295674 243704
rect 359458 243692 359464 243704
rect 295668 243664 359464 243692
rect 295668 243652 295674 243664
rect 359458 243652 359464 243664
rect 359516 243652 359522 243704
rect 217502 243584 217508 243636
rect 217560 243624 217566 243636
rect 294046 243624 294052 243636
rect 217560 243596 294052 243624
rect 217560 243584 217566 243596
rect 294046 243584 294052 243596
rect 294104 243584 294110 243636
rect 295518 243584 295524 243636
rect 295576 243624 295582 243636
rect 360838 243624 360844 243636
rect 295576 243596 360844 243624
rect 295576 243584 295582 243596
rect 360838 243584 360844 243596
rect 360896 243584 360902 243636
rect 215754 243516 215760 243568
rect 215812 243556 215818 243568
rect 293126 243556 293132 243568
rect 215812 243528 293132 243556
rect 215812 243516 215818 243528
rect 293126 243516 293132 243528
rect 293184 243516 293190 243568
rect 295334 243516 295340 243568
rect 295392 243556 295398 243568
rect 362126 243556 362132 243568
rect 295392 243528 362132 243556
rect 295392 243516 295398 243528
rect 362126 243516 362132 243528
rect 362184 243516 362190 243568
rect 3510 241408 3516 241460
rect 3568 241448 3574 241460
rect 14550 241448 14556 241460
rect 3568 241420 14556 241448
rect 3568 241408 3574 241420
rect 14550 241408 14556 241420
rect 14608 241408 14614 241460
rect 577590 219172 577596 219224
rect 577648 219212 577654 219224
rect 579706 219212 579712 219224
rect 577648 219184 579712 219212
rect 577648 219172 577654 219184
rect 579706 219172 579712 219184
rect 579764 219172 579770 219224
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 209038 215268 209044 215280
rect 3384 215240 209044 215268
rect 3384 215228 3390 215240
rect 209038 215228 209044 215240
rect 209096 215228 209102 215280
rect 358078 206932 358084 206984
rect 358136 206972 358142 206984
rect 579614 206972 579620 206984
rect 358136 206944 579620 206972
rect 358136 206932 358142 206944
rect 579614 206932 579620 206944
rect 579672 206932 579678 206984
rect 358354 204824 358360 204876
rect 358412 204864 358418 204876
rect 363782 204864 363788 204876
rect 358412 204836 363788 204864
rect 358412 204824 358418 204836
rect 363782 204824 363788 204836
rect 363840 204824 363846 204876
rect 358262 204688 358268 204740
rect 358320 204728 358326 204740
rect 363782 204728 363788 204740
rect 358320 204700 363788 204728
rect 358320 204688 358326 204700
rect 363782 204688 363788 204700
rect 363840 204688 363846 204740
rect 3050 202784 3056 202836
rect 3108 202824 3114 202836
rect 199378 202824 199384 202836
rect 3108 202796 199384 202824
rect 3108 202784 3114 202796
rect 199378 202784 199384 202796
rect 199436 202784 199442 202836
rect 214374 195508 214380 195560
rect 214432 195548 214438 195560
rect 217134 195548 217140 195560
rect 214432 195520 217140 195548
rect 214432 195508 214438 195520
rect 217134 195508 217140 195520
rect 217192 195508 217198 195560
rect 212994 195236 213000 195288
rect 213052 195276 213058 195288
rect 217318 195276 217324 195288
rect 213052 195248 217324 195276
rect 213052 195236 213058 195248
rect 217318 195236 217324 195248
rect 217376 195236 217382 195288
rect 210878 193128 210884 193180
rect 210936 193168 210942 193180
rect 216766 193168 216772 193180
rect 210936 193140 216772 193168
rect 210936 193128 210942 193140
rect 216766 193128 216772 193140
rect 216824 193128 216830 193180
rect 215846 189388 215852 189440
rect 215904 189428 215910 189440
rect 218514 189428 218520 189440
rect 215904 189400 218520 189428
rect 215904 189388 215910 189400
rect 218514 189388 218520 189400
rect 218572 189388 218578 189440
rect 3510 188980 3516 189032
rect 3568 189020 3574 189032
rect 206278 189020 206284 189032
rect 3568 188992 206284 189020
rect 3568 188980 3574 188992
rect 206278 188980 206284 188992
rect 206336 188980 206342 189032
rect 210970 188980 210976 189032
rect 211028 189020 211034 189032
rect 216674 189020 216680 189032
rect 211028 188992 216680 189020
rect 211028 188980 211034 188992
rect 216674 188980 216680 188992
rect 216732 188980 216738 189032
rect 577498 179324 577504 179376
rect 577556 179364 577562 179376
rect 579706 179364 579712 179376
rect 577556 179336 579712 179364
rect 577556 179324 577562 179336
rect 579706 179324 579712 179336
rect 579764 179324 579770 179376
rect 212074 159876 212080 159928
rect 212132 159916 212138 159928
rect 256694 159916 256700 159928
rect 212132 159888 256700 159916
rect 212132 159876 212138 159888
rect 256694 159876 256700 159888
rect 256752 159876 256758 159928
rect 218790 159808 218796 159860
rect 218848 159848 218854 159860
rect 264974 159848 264980 159860
rect 218848 159820 264980 159848
rect 218848 159808 218854 159820
rect 264974 159808 264980 159820
rect 265032 159808 265038 159860
rect 216306 159740 216312 159792
rect 216364 159780 216370 159792
rect 263594 159780 263600 159792
rect 216364 159752 263600 159780
rect 216364 159740 216370 159752
rect 263594 159740 263600 159752
rect 263652 159740 263658 159792
rect 213454 159672 213460 159724
rect 213512 159712 213518 159724
rect 260834 159712 260840 159724
rect 213512 159684 260840 159712
rect 213512 159672 213518 159684
rect 260834 159672 260840 159684
rect 260892 159672 260898 159724
rect 213086 159604 213092 159656
rect 213144 159644 213150 159656
rect 269114 159644 269120 159656
rect 213144 159616 269120 159644
rect 213144 159604 213150 159616
rect 269114 159604 269120 159616
rect 269172 159604 269178 159656
rect 217134 159536 217140 159588
rect 217192 159576 217198 159588
rect 276198 159576 276204 159588
rect 217192 159548 276204 159576
rect 217192 159536 217198 159548
rect 276198 159536 276204 159548
rect 276256 159536 276262 159588
rect 313458 159536 313464 159588
rect 313516 159576 313522 159588
rect 373258 159576 373264 159588
rect 313516 159548 373264 159576
rect 313516 159536 313522 159548
rect 373258 159536 373264 159548
rect 373316 159536 373322 159588
rect 215938 159468 215944 159520
rect 215996 159508 216002 159520
rect 276014 159508 276020 159520
rect 215996 159480 276020 159508
rect 215996 159468 216002 159480
rect 276014 159468 276020 159480
rect 276072 159468 276078 159520
rect 298462 159468 298468 159520
rect 298520 159508 298526 159520
rect 358170 159508 358176 159520
rect 298520 159480 358176 159508
rect 298520 159468 298526 159480
rect 358170 159468 358176 159480
rect 358228 159468 358234 159520
rect 217870 159400 217876 159452
rect 217928 159440 217934 159452
rect 278774 159440 278780 159452
rect 217928 159412 278780 159440
rect 217928 159400 217934 159412
rect 278774 159400 278780 159412
rect 278832 159400 278838 159452
rect 310974 159400 310980 159452
rect 311032 159440 311038 159452
rect 371602 159440 371608 159452
rect 311032 159412 371608 159440
rect 311032 159400 311038 159412
rect 371602 159400 371608 159412
rect 371660 159400 371666 159452
rect 214466 159332 214472 159384
rect 214524 159372 214530 159384
rect 282914 159372 282920 159384
rect 214524 159344 282920 159372
rect 214524 159332 214530 159344
rect 282914 159332 282920 159344
rect 282972 159332 282978 159384
rect 303522 159332 303528 159384
rect 303580 159372 303586 159384
rect 369210 159372 369216 159384
rect 303580 159344 369216 159372
rect 303580 159332 303586 159344
rect 369210 159332 369216 159344
rect 369268 159332 369274 159384
rect 295886 159264 295892 159316
rect 295944 159304 295950 159316
rect 369118 159304 369124 159316
rect 295944 159276 369124 159304
rect 295944 159264 295950 159276
rect 369118 159264 369124 159276
rect 369176 159264 369182 159316
rect 293494 159196 293500 159248
rect 293552 159236 293558 159248
rect 370682 159236 370688 159248
rect 293552 159208 370688 159236
rect 293552 159196 293558 159208
rect 370682 159196 370688 159208
rect 370740 159196 370746 159248
rect 276106 159128 276112 159180
rect 276164 159168 276170 159180
rect 363690 159168 363696 159180
rect 276164 159140 363696 159168
rect 276164 159128 276170 159140
rect 363690 159128 363696 159140
rect 363748 159128 363754 159180
rect 278498 159060 278504 159112
rect 278556 159100 278562 159112
rect 367922 159100 367928 159112
rect 278556 159072 367928 159100
rect 278556 159060 278562 159072
rect 367922 159060 367928 159072
rect 367980 159060 367986 159112
rect 273622 158992 273628 159044
rect 273680 159032 273686 159044
rect 367830 159032 367836 159044
rect 273680 159004 367836 159032
rect 273680 158992 273686 159004
rect 367830 158992 367836 159004
rect 367888 158992 367894 159044
rect 213270 158924 213276 158976
rect 213328 158964 213334 158976
rect 238202 158964 238208 158976
rect 213328 158936 238208 158964
rect 213328 158924 213334 158936
rect 238202 158924 238208 158936
rect 238260 158924 238266 158976
rect 265342 158924 265348 158976
rect 265400 158964 265406 158976
rect 359642 158964 359648 158976
rect 265400 158936 359648 158964
rect 265400 158924 265406 158936
rect 359642 158924 359648 158936
rect 359700 158924 359706 158976
rect 213178 158856 213184 158908
rect 213236 158896 213242 158908
rect 239582 158896 239588 158908
rect 213236 158868 239588 158896
rect 213236 158856 213242 158868
rect 239582 158856 239588 158868
rect 239640 158856 239646 158908
rect 263962 158856 263968 158908
rect 264020 158896 264026 158908
rect 363598 158896 363604 158908
rect 264020 158868 363604 158896
rect 264020 158856 264026 158868
rect 363598 158856 363604 158868
rect 363656 158856 363662 158908
rect 213362 158788 213368 158840
rect 213420 158828 213426 158840
rect 241698 158828 241704 158840
rect 213420 158800 241704 158828
rect 213420 158788 213426 158800
rect 241698 158788 241704 158800
rect 241756 158788 241762 158840
rect 262858 158788 262864 158840
rect 262916 158828 262922 158840
rect 364610 158828 364616 158840
rect 262916 158800 364616 158828
rect 262916 158788 262922 158800
rect 364610 158788 364616 158800
rect 364668 158788 364674 158840
rect 211982 158720 211988 158772
rect 212040 158760 212046 158772
rect 240502 158760 240508 158772
rect 212040 158732 240508 158760
rect 212040 158720 212046 158732
rect 240502 158720 240508 158732
rect 240560 158720 240566 158772
rect 259546 158720 259552 158772
rect 259604 158760 259610 158772
rect 364702 158760 364708 158772
rect 259604 158732 364708 158760
rect 259604 158720 259610 158732
rect 364702 158720 364708 158732
rect 364760 158720 364766 158772
rect 219066 158652 219072 158704
rect 219124 158692 219130 158704
rect 234614 158692 234620 158704
rect 219124 158664 234620 158692
rect 219124 158652 219130 158664
rect 234614 158652 234620 158664
rect 234672 158652 234678 158704
rect 248322 158652 248328 158704
rect 248380 158692 248386 158704
rect 365162 158692 365168 158704
rect 248380 158664 365168 158692
rect 248380 158652 248386 158664
rect 365162 158652 365168 158664
rect 365220 158652 365226 158704
rect 216122 158584 216128 158636
rect 216180 158624 216186 158636
rect 233234 158624 233240 158636
rect 216180 158596 233240 158624
rect 216180 158584 216186 158596
rect 233234 158584 233240 158596
rect 233292 158584 233298 158636
rect 256050 158584 256056 158636
rect 256108 158624 256114 158636
rect 371786 158624 371792 158636
rect 256108 158596 371792 158624
rect 256108 158584 256114 158596
rect 371786 158584 371792 158596
rect 371844 158584 371850 158636
rect 214834 158516 214840 158568
rect 214892 158556 214898 158568
rect 235994 158556 236000 158568
rect 214892 158528 236000 158556
rect 214892 158516 214898 158528
rect 235994 158516 236000 158528
rect 236052 158516 236058 158568
rect 261202 158516 261208 158568
rect 261260 158556 261266 158568
rect 373166 158556 373172 158568
rect 261260 158528 373172 158556
rect 261260 158516 261266 158528
rect 373166 158516 373172 158528
rect 373224 158516 373230 158568
rect 211890 158448 211896 158500
rect 211948 158488 211954 158500
rect 234706 158488 234712 158500
rect 211948 158460 234712 158488
rect 211948 158448 211954 158460
rect 234706 158448 234712 158460
rect 234764 158448 234770 158500
rect 255958 158448 255964 158500
rect 256016 158488 256022 158500
rect 364426 158488 364432 158500
rect 256016 158460 364432 158488
rect 256016 158448 256022 158460
rect 364426 158448 364432 158460
rect 364484 158448 364490 158500
rect 218974 158380 218980 158432
rect 219032 158420 219038 158432
rect 242986 158420 242992 158432
rect 219032 158392 242992 158420
rect 219032 158380 219038 158392
rect 242986 158380 242992 158392
rect 243044 158380 243050 158432
rect 257154 158380 257160 158432
rect 257212 158420 257218 158432
rect 364334 158420 364340 158432
rect 257212 158392 364340 158420
rect 257212 158380 257218 158392
rect 364334 158380 364340 158392
rect 364392 158380 364398 158432
rect 214650 158312 214656 158364
rect 214708 158352 214714 158364
rect 242894 158352 242900 158364
rect 214708 158324 242900 158352
rect 214708 158312 214714 158324
rect 242894 158312 242900 158324
rect 242952 158312 242958 158364
rect 254578 158312 254584 158364
rect 254636 158352 254642 158364
rect 360930 158352 360936 158364
rect 254636 158324 360936 158352
rect 254636 158312 254642 158324
rect 360930 158312 360936 158324
rect 360988 158312 360994 158364
rect 214926 158244 214932 158296
rect 214984 158284 214990 158296
rect 245654 158284 245660 158296
rect 214984 158256 245660 158284
rect 214984 158244 214990 158256
rect 245654 158244 245660 158256
rect 245712 158244 245718 158296
rect 258258 158244 258264 158296
rect 258316 158284 258322 158296
rect 364518 158284 364524 158296
rect 258316 158256 364524 158284
rect 258316 158244 258322 158256
rect 364518 158244 364524 158256
rect 364576 158244 364582 158296
rect 216214 158176 216220 158228
rect 216272 158216 216278 158228
rect 247034 158216 247040 158228
rect 216272 158188 247040 158216
rect 216272 158176 216278 158188
rect 247034 158176 247040 158188
rect 247092 158176 247098 158228
rect 265986 158176 265992 158228
rect 266044 158216 266050 158228
rect 369302 158216 369308 158228
rect 266044 158188 369308 158216
rect 266044 158176 266050 158188
rect 369302 158176 369308 158188
rect 369360 158176 369366 158228
rect 216398 158108 216404 158160
rect 216456 158148 216462 158160
rect 249794 158148 249800 158160
rect 216456 158120 249800 158148
rect 216456 158108 216462 158120
rect 249794 158108 249800 158120
rect 249852 158108 249858 158160
rect 291010 158108 291016 158160
rect 291068 158148 291074 158160
rect 370590 158148 370596 158160
rect 291068 158120 370596 158148
rect 291068 158108 291074 158120
rect 370590 158108 370596 158120
rect 370648 158108 370654 158160
rect 218882 158040 218888 158092
rect 218940 158080 218946 158092
rect 252554 158080 252560 158092
rect 218940 158052 252560 158080
rect 218940 158040 218946 158052
rect 252554 158040 252560 158052
rect 252612 158040 252618 158092
rect 300946 158040 300952 158092
rect 301004 158080 301010 158092
rect 370498 158080 370504 158092
rect 301004 158052 370504 158080
rect 301004 158040 301010 158052
rect 370498 158040 370504 158052
rect 370556 158040 370562 158092
rect 211614 157972 211620 158024
rect 211672 158012 211678 158024
rect 273254 158012 273260 158024
rect 211672 157984 273260 158012
rect 211672 157972 211678 157984
rect 273254 157972 273260 157984
rect 273312 157972 273318 158024
rect 308674 157972 308680 158024
rect 308732 158012 308738 158024
rect 372982 158012 372988 158024
rect 308732 157984 372988 158012
rect 308732 157972 308738 157984
rect 372982 157972 372988 157984
rect 373040 157972 373046 158024
rect 216030 157904 216036 157956
rect 216088 157944 216094 157956
rect 230474 157944 230480 157956
rect 216088 157916 230480 157944
rect 216088 157904 216094 157916
rect 230474 157904 230480 157916
rect 230532 157904 230538 157956
rect 321094 157904 321100 157956
rect 321152 157944 321158 157956
rect 371694 157944 371700 157956
rect 321152 157916 371700 157944
rect 321152 157904 321158 157916
rect 371694 157904 371700 157916
rect 371752 157904 371758 157956
rect 214742 157836 214748 157888
rect 214800 157876 214806 157888
rect 229094 157876 229100 157888
rect 214800 157848 229100 157876
rect 214800 157836 214806 157848
rect 229094 157836 229100 157848
rect 229152 157836 229158 157888
rect 323394 157836 323400 157888
rect 323452 157876 323458 157888
rect 371878 157876 371884 157888
rect 323452 157848 371884 157876
rect 323452 157836 323458 157848
rect 371878 157836 371884 157848
rect 371936 157836 371942 157888
rect 219158 157768 219164 157820
rect 219216 157808 219222 157820
rect 227714 157808 227720 157820
rect 219216 157780 227720 157808
rect 219216 157768 219222 157780
rect 227714 157768 227720 157780
rect 227772 157768 227778 157820
rect 325970 157768 325976 157820
rect 326028 157808 326034 157820
rect 373074 157808 373080 157820
rect 326028 157780 373080 157808
rect 326028 157768 326034 157780
rect 373074 157768 373080 157780
rect 373132 157768 373138 157820
rect 250162 157292 250168 157344
rect 250220 157332 250226 157344
rect 368566 157332 368572 157344
rect 250220 157304 368572 157332
rect 250220 157292 250226 157304
rect 368566 157292 368572 157304
rect 368624 157292 368630 157344
rect 251450 157224 251456 157276
rect 251508 157264 251514 157276
rect 368842 157264 368848 157276
rect 251508 157236 368848 157264
rect 251508 157224 251514 157236
rect 368842 157224 368848 157236
rect 368900 157224 368906 157276
rect 267642 157156 267648 157208
rect 267700 157196 267706 157208
rect 367370 157196 367376 157208
rect 267700 157168 367376 157196
rect 267700 157156 267706 157168
rect 367370 157156 367376 157168
rect 367428 157156 367434 157208
rect 268746 157088 268752 157140
rect 268804 157128 268810 157140
rect 367646 157128 367652 157140
rect 268804 157100 367652 157128
rect 268804 157088 268810 157100
rect 367646 157088 367652 157100
rect 367704 157088 367710 157140
rect 271138 157020 271144 157072
rect 271196 157060 271202 157072
rect 367738 157060 367744 157072
rect 271196 157032 367744 157060
rect 271196 157020 271202 157032
rect 367738 157020 367744 157032
rect 367796 157020 367802 157072
rect 266814 156952 266820 157004
rect 266872 156992 266878 157004
rect 363506 156992 363512 157004
rect 266872 156964 363512 156992
rect 266872 156952 266878 156964
rect 363506 156952 363512 156964
rect 363564 156952 363570 157004
rect 269850 156884 269856 156936
rect 269908 156924 269914 156936
rect 365898 156924 365904 156936
rect 269908 156896 365904 156924
rect 269908 156884 269914 156896
rect 365898 156884 365904 156896
rect 365956 156884 365962 156936
rect 272242 156816 272248 156868
rect 272300 156856 272306 156868
rect 366266 156856 366272 156868
rect 272300 156828 366272 156856
rect 272300 156816 272306 156828
rect 366266 156816 366272 156828
rect 366324 156816 366330 156868
rect 274174 156748 274180 156800
rect 274232 156788 274238 156800
rect 367554 156788 367560 156800
rect 274232 156760 367560 156788
rect 274232 156748 274238 156760
rect 367554 156748 367560 156760
rect 367612 156748 367618 156800
rect 274450 156680 274456 156732
rect 274508 156720 274514 156732
rect 366358 156720 366364 156732
rect 274508 156692 366364 156720
rect 274508 156680 274514 156692
rect 366358 156680 366364 156692
rect 366416 156680 366422 156732
rect 275922 156612 275928 156664
rect 275980 156652 275986 156664
rect 367278 156652 367284 156664
rect 275980 156624 367284 156652
rect 275980 156612 275986 156624
rect 367278 156612 367284 156624
rect 367336 156612 367342 156664
rect 277118 156544 277124 156596
rect 277176 156584 277182 156596
rect 366082 156584 366088 156596
rect 277176 156556 366088 156584
rect 277176 156544 277182 156556
rect 366082 156544 366088 156556
rect 366140 156544 366146 156596
rect 279970 156476 279976 156528
rect 280028 156516 280034 156528
rect 366174 156516 366180 156528
rect 280028 156488 366180 156516
rect 280028 156476 280034 156488
rect 366174 156476 366180 156488
rect 366232 156476 366238 156528
rect 278130 156408 278136 156460
rect 278188 156448 278194 156460
rect 361114 156448 361120 156460
rect 278188 156420 361120 156448
rect 278188 156408 278194 156420
rect 361114 156408 361120 156420
rect 361172 156408 361178 156460
rect 252370 155864 252376 155916
rect 252428 155904 252434 155916
rect 368658 155904 368664 155916
rect 252428 155876 368664 155904
rect 252428 155864 252434 155876
rect 368658 155864 368664 155876
rect 368716 155864 368722 155916
rect 251082 155796 251088 155848
rect 251140 155836 251146 155848
rect 366450 155836 366456 155848
rect 251140 155808 366456 155836
rect 251140 155796 251146 155808
rect 366450 155796 366456 155808
rect 366508 155796 366514 155848
rect 213546 155728 213552 155780
rect 213604 155768 213610 155780
rect 237374 155768 237380 155780
rect 213604 155740 237380 155768
rect 213604 155728 213610 155740
rect 237374 155728 237380 155740
rect 237432 155728 237438 155780
rect 253566 155728 253572 155780
rect 253624 155768 253630 155780
rect 367462 155768 367468 155780
rect 253624 155740 367468 155768
rect 253624 155728 253630 155740
rect 367462 155728 367468 155740
rect 367520 155728 367526 155780
rect 211798 155660 211804 155712
rect 211856 155700 211862 155712
rect 241514 155700 241520 155712
rect 211856 155672 241520 155700
rect 211856 155660 211862 155672
rect 241514 155660 241520 155672
rect 241572 155660 241578 155712
rect 268930 155660 268936 155712
rect 268988 155700 268994 155712
rect 365070 155700 365076 155712
rect 268988 155672 365076 155700
rect 268988 155660 268994 155672
rect 365070 155660 365076 155672
rect 365128 155660 365134 155712
rect 214558 155592 214564 155644
rect 214616 155632 214622 155644
rect 248414 155632 248420 155644
rect 214616 155604 248420 155632
rect 214616 155592 214622 155604
rect 248414 155592 248420 155604
rect 248472 155592 248478 155644
rect 281074 155592 281080 155644
rect 281132 155632 281138 155644
rect 370222 155632 370228 155644
rect 281132 155604 370228 155632
rect 281132 155592 281138 155604
rect 370222 155592 370228 155604
rect 370280 155592 370286 155644
rect 211062 155524 211068 155576
rect 211120 155564 211126 155576
rect 255314 155564 255320 155576
rect 211120 155536 255320 155564
rect 211120 155524 211126 155536
rect 255314 155524 255320 155536
rect 255372 155524 255378 155576
rect 283742 155524 283748 155576
rect 283800 155564 283806 155576
rect 370038 155564 370044 155576
rect 283800 155536 370044 155564
rect 283800 155524 283806 155536
rect 370038 155524 370044 155536
rect 370096 155524 370102 155576
rect 211706 155456 211712 155508
rect 211764 155496 211770 155508
rect 259546 155496 259552 155508
rect 211764 155468 259552 155496
rect 211764 155456 211770 155468
rect 259546 155456 259552 155468
rect 259604 155456 259610 155508
rect 286502 155456 286508 155508
rect 286560 155496 286566 155508
rect 370130 155496 370136 155508
rect 286560 155468 370136 155496
rect 286560 155456 286566 155468
rect 370130 155456 370136 155468
rect 370188 155456 370194 155508
rect 218606 155388 218612 155440
rect 218664 155428 218670 155440
rect 280154 155428 280160 155440
rect 218664 155400 280160 155428
rect 218664 155388 218670 155400
rect 280154 155388 280160 155400
rect 280212 155388 280218 155440
rect 348510 155388 348516 155440
rect 348568 155428 348574 155440
rect 369026 155428 369032 155440
rect 348568 155400 369032 155428
rect 348568 155388 348574 155400
rect 369026 155388 369032 155400
rect 369084 155388 369090 155440
rect 218514 155320 218520 155372
rect 218572 155360 218578 155372
rect 284386 155360 284392 155372
rect 218572 155332 284392 155360
rect 218572 155320 218578 155332
rect 284386 155320 284392 155332
rect 284444 155320 284450 155372
rect 292574 155320 292580 155372
rect 292632 155360 292638 155372
rect 357986 155360 357992 155372
rect 292632 155332 357992 155360
rect 292632 155320 292638 155332
rect 357986 155320 357992 155332
rect 358044 155320 358050 155372
rect 217502 155252 217508 155304
rect 217560 155292 217566 155304
rect 285674 155292 285680 155304
rect 217560 155264 285680 155292
rect 217560 155252 217566 155264
rect 285674 155252 285680 155264
rect 285732 155252 285738 155304
rect 292666 155252 292672 155304
rect 292724 155292 292730 155304
rect 363782 155292 363788 155304
rect 292724 155264 363788 155292
rect 292724 155252 292730 155264
rect 363782 155252 363788 155264
rect 363840 155252 363846 155304
rect 215754 155184 215760 155236
rect 215812 155224 215818 155236
rect 284294 155224 284300 155236
rect 215812 155196 284300 155224
rect 215812 155184 215818 155196
rect 284294 155184 284300 155196
rect 284352 155184 284358 155236
rect 289814 155184 289820 155236
rect 289872 155224 289878 155236
rect 370406 155224 370412 155236
rect 289872 155196 370412 155224
rect 289872 155184 289878 155196
rect 370406 155184 370412 155196
rect 370464 155184 370470 155236
rect 348418 155116 348424 155168
rect 348476 155156 348482 155168
rect 366542 155156 366548 155168
rect 348476 155128 366548 155156
rect 348476 155116 348482 155128
rect 366542 155116 366548 155128
rect 366600 155116 366606 155168
rect 253658 154504 253664 154556
rect 253716 154544 253722 154556
rect 372890 154544 372896 154556
rect 253716 154516 372896 154544
rect 253716 154504 253722 154516
rect 372890 154504 372896 154516
rect 372948 154504 372954 154556
rect 258626 154436 258632 154488
rect 258684 154476 258690 154488
rect 370314 154476 370320 154488
rect 258684 154448 370320 154476
rect 258684 154436 258690 154448
rect 370314 154436 370320 154448
rect 370372 154436 370378 154488
rect 263962 154368 263968 154420
rect 264020 154408 264026 154420
rect 371418 154408 371424 154420
rect 264020 154380 371424 154408
rect 264020 154368 264026 154380
rect 371418 154368 371424 154380
rect 371476 154368 371482 154420
rect 271046 154300 271052 154352
rect 271104 154340 271110 154352
rect 372798 154340 372804 154352
rect 271104 154312 372804 154340
rect 271104 154300 271110 154312
rect 372798 154300 372804 154312
rect 372856 154300 372862 154352
rect 288250 154232 288256 154284
rect 288308 154272 288314 154284
rect 369946 154272 369952 154284
rect 288308 154244 369952 154272
rect 288308 154232 288314 154244
rect 369946 154232 369952 154244
rect 370004 154232 370010 154284
rect 306098 154164 306104 154216
rect 306156 154204 306162 154216
rect 371326 154204 371332 154216
rect 306156 154176 371332 154204
rect 306156 154164 306162 154176
rect 371326 154164 371332 154176
rect 371384 154164 371390 154216
rect 315850 154096 315856 154148
rect 315908 154136 315914 154148
rect 371510 154136 371516 154148
rect 315908 154108 371516 154136
rect 315908 154096 315914 154108
rect 371510 154096 371516 154108
rect 371568 154096 371574 154148
rect 318610 154028 318616 154080
rect 318668 154068 318674 154080
rect 372706 154068 372712 154080
rect 318668 154040 372712 154068
rect 318668 154028 318674 154040
rect 372706 154028 372712 154040
rect 372764 154028 372770 154080
rect 3510 150356 3516 150408
rect 3568 150396 3574 150408
rect 210418 150396 210424 150408
rect 3568 150368 210424 150396
rect 3568 150356 3574 150368
rect 210418 150356 210424 150368
rect 210476 150356 210482 150408
rect 3510 137912 3516 137964
rect 3568 137952 3574 137964
rect 203518 137952 203524 137964
rect 3568 137924 203524 137952
rect 3568 137912 3574 137924
rect 203518 137912 203524 137924
rect 203576 137912 203582 137964
rect 3510 97928 3516 97980
rect 3568 97968 3574 97980
rect 197998 97968 198004 97980
rect 3568 97940 198004 97968
rect 3568 97928 3574 97940
rect 197998 97928 198004 97940
rect 198056 97928 198062 97980
rect 3510 85484 3516 85536
rect 3568 85524 3574 85536
rect 200758 85524 200764 85536
rect 3568 85496 200764 85524
rect 3568 85484 3574 85496
rect 200758 85484 200764 85496
rect 200816 85484 200822 85536
rect 3510 71680 3516 71732
rect 3568 71720 3574 71732
rect 207658 71720 207664 71732
rect 3568 71692 207664 71720
rect 3568 71680 3574 71692
rect 207658 71680 207664 71692
rect 207716 71680 207722 71732
rect 3510 59304 3516 59356
rect 3568 59344 3574 59356
rect 25498 59344 25504 59356
rect 3568 59316 25504 59344
rect 3568 59304 3574 59316
rect 25498 59304 25504 59316
rect 25556 59304 25562 59356
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 196618 20652 196624 20664
rect 3476 20624 196624 20652
rect 3476 20612 3482 20624
rect 196618 20612 196624 20624
rect 196676 20612 196682 20664
rect 160094 11704 160100 11756
rect 160152 11744 160158 11756
rect 161290 11744 161296 11756
rect 160152 11716 161296 11744
rect 160152 11704 160158 11716
rect 161290 11704 161296 11716
rect 161348 11704 161354 11756
rect 201494 11704 201500 11756
rect 201552 11744 201558 11756
rect 202690 11744 202696 11756
rect 201552 11716 202696 11744
rect 201552 11704 201558 11716
rect 202690 11704 202696 11716
rect 202748 11704 202754 11756
rect 234614 11704 234620 11756
rect 234672 11744 234678 11756
rect 235810 11744 235816 11756
rect 234672 11716 235816 11744
rect 234672 11704 234678 11716
rect 235810 11704 235816 11716
rect 235868 11704 235874 11756
rect 242894 11704 242900 11756
rect 242952 11744 242958 11756
rect 244090 11744 244096 11756
rect 242952 11716 244096 11744
rect 242952 11704 242958 11716
rect 244090 11704 244096 11716
rect 244148 11704 244154 11756
rect 316218 9324 316224 9376
rect 316276 9364 316282 9376
rect 363414 9364 363420 9376
rect 316276 9336 363420 9364
rect 316276 9324 316282 9336
rect 363414 9324 363420 9336
rect 363472 9324 363478 9376
rect 312630 9256 312636 9308
rect 312688 9296 312694 9308
rect 360286 9296 360292 9308
rect 312688 9268 360292 9296
rect 312688 9256 312694 9268
rect 360286 9256 360292 9268
rect 360344 9256 360350 9308
rect 298462 9188 298468 9240
rect 298520 9228 298526 9240
rect 357894 9228 357900 9240
rect 298520 9200 357900 9228
rect 298520 9188 298526 9200
rect 357894 9188 357900 9200
rect 357952 9188 357958 9240
rect 301958 9120 301964 9172
rect 302016 9160 302022 9172
rect 362126 9160 362132 9172
rect 302016 9132 362132 9160
rect 302016 9120 302022 9132
rect 362126 9120 362132 9132
rect 362184 9120 362190 9172
rect 300762 9052 300768 9104
rect 300820 9092 300826 9104
rect 360838 9092 360844 9104
rect 300820 9064 360844 9092
rect 300820 9052 300826 9064
rect 360838 9052 360844 9064
rect 360896 9052 360902 9104
rect 304350 8984 304356 9036
rect 304408 9024 304414 9036
rect 365806 9024 365812 9036
rect 304408 8996 365812 9024
rect 304408 8984 304414 8996
rect 365806 8984 365812 8996
rect 365864 8984 365870 9036
rect 297266 8916 297272 8968
rect 297324 8956 297330 8968
rect 359458 8956 359464 8968
rect 297324 8928 359464 8956
rect 297324 8916 297330 8928
rect 359458 8916 359464 8928
rect 359516 8916 359522 8968
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 88978 6848 88984 6860
rect 3476 6820 88984 6848
rect 3476 6808 3482 6820
rect 88978 6808 88984 6820
rect 89036 6808 89042 6860
rect 317322 6808 317328 6860
rect 317380 6848 317386 6860
rect 358814 6848 358820 6860
rect 317380 6820 358820 6848
rect 317380 6808 317386 6820
rect 358814 6808 358820 6820
rect 358872 6808 358878 6860
rect 322106 6740 322112 6792
rect 322164 6780 322170 6792
rect 368474 6780 368480 6792
rect 322164 6752 368480 6780
rect 322164 6740 322170 6752
rect 368474 6740 368480 6752
rect 368532 6740 368538 6792
rect 320910 6672 320916 6724
rect 320968 6712 320974 6724
rect 367094 6712 367100 6724
rect 320968 6684 367100 6712
rect 320968 6672 320974 6684
rect 367094 6672 367100 6684
rect 367152 6672 367158 6724
rect 315022 6604 315028 6656
rect 315080 6644 315086 6656
rect 361574 6644 361580 6656
rect 315080 6616 361580 6644
rect 315080 6604 315086 6616
rect 361574 6604 361580 6616
rect 361632 6604 361638 6656
rect 313826 6536 313832 6588
rect 313884 6576 313890 6588
rect 360654 6576 360660 6588
rect 313884 6548 360660 6576
rect 313884 6536 313890 6548
rect 360654 6536 360660 6548
rect 360712 6536 360718 6588
rect 318518 6468 318524 6520
rect 318576 6508 318582 6520
rect 365714 6508 365720 6520
rect 318576 6480 365720 6508
rect 318576 6468 318582 6480
rect 365714 6468 365720 6480
rect 365772 6468 365778 6520
rect 310238 6400 310244 6452
rect 310296 6440 310302 6452
rect 357802 6440 357808 6452
rect 310296 6412 357808 6440
rect 310296 6400 310302 6412
rect 357802 6400 357808 6412
rect 357860 6400 357866 6452
rect 311434 6332 311440 6384
rect 311492 6372 311498 6384
rect 359366 6372 359372 6384
rect 311492 6344 359372 6372
rect 311492 6332 311498 6344
rect 359366 6332 359372 6344
rect 359424 6332 359430 6384
rect 307938 6264 307944 6316
rect 307996 6304 308002 6316
rect 356790 6304 356796 6316
rect 307996 6276 356796 6304
rect 307996 6264 308002 6276
rect 356790 6264 356796 6276
rect 356848 6264 356854 6316
rect 306742 6196 306748 6248
rect 306800 6236 306806 6248
rect 367186 6236 367192 6248
rect 306800 6208 367192 6236
rect 306800 6196 306806 6208
rect 367186 6196 367192 6208
rect 367244 6196 367250 6248
rect 303154 6128 303160 6180
rect 303212 6168 303218 6180
rect 363322 6168 363328 6180
rect 303212 6140 363328 6168
rect 303212 6128 303218 6140
rect 363322 6128 363328 6140
rect 363380 6128 363386 6180
rect 326798 6060 326804 6112
rect 326856 6100 326862 6112
rect 360746 6100 360752 6112
rect 326856 6072 360752 6100
rect 326856 6060 326862 6072
rect 360746 6060 360752 6072
rect 360804 6060 360810 6112
rect 323302 5992 323308 6044
rect 323360 6032 323366 6044
rect 357710 6032 357716 6044
rect 323360 6004 357716 6032
rect 323360 5992 323366 6004
rect 357710 5992 357716 6004
rect 357768 5992 357774 6044
rect 330386 5924 330392 5976
rect 330444 5964 330450 5976
rect 363138 5964 363144 5976
rect 330444 5936 363144 5964
rect 330444 5924 330450 5936
rect 363138 5924 363144 5936
rect 363196 5924 363202 5976
rect 44266 4088 44272 4140
rect 44324 4128 44330 4140
rect 46198 4128 46204 4140
rect 44324 4100 46204 4128
rect 44324 4088 44330 4100
rect 46198 4088 46204 4100
rect 46256 4088 46262 4140
rect 213822 4088 213828 4140
rect 213880 4128 213886 4140
rect 260650 4128 260656 4140
rect 213880 4100 260656 4128
rect 213880 4088 213886 4100
rect 260650 4088 260656 4100
rect 260708 4088 260714 4140
rect 332686 4088 332692 4140
rect 332744 4128 332750 4140
rect 360470 4128 360476 4140
rect 332744 4100 360476 4128
rect 332744 4088 332750 4100
rect 360470 4088 360476 4100
rect 360528 4088 360534 4140
rect 467098 4088 467104 4140
rect 467156 4128 467162 4140
rect 467650 4128 467656 4140
rect 467156 4100 467656 4128
rect 467156 4088 467162 4100
rect 467650 4088 467656 4100
rect 467708 4088 467714 4140
rect 219342 4020 219348 4072
rect 219400 4060 219406 4072
rect 266538 4060 266544 4072
rect 219400 4032 266544 4060
rect 219400 4020 219406 4032
rect 266538 4020 266544 4032
rect 266596 4020 266602 4072
rect 327994 4020 328000 4072
rect 328052 4060 328058 4072
rect 359182 4060 359188 4072
rect 328052 4032 359188 4060
rect 328052 4020 328058 4032
rect 359182 4020 359188 4032
rect 359240 4020 359246 4072
rect 177850 3952 177856 4004
rect 177908 3992 177914 4004
rect 181438 3992 181444 4004
rect 177908 3964 181444 3992
rect 177908 3952 177914 3964
rect 181438 3952 181444 3964
rect 181496 3952 181502 4004
rect 216582 3952 216588 4004
rect 216640 3992 216646 4004
rect 267734 3992 267740 4004
rect 216640 3964 267740 3992
rect 216640 3952 216646 3964
rect 267734 3952 267740 3964
rect 267792 3952 267798 4004
rect 324406 3952 324412 4004
rect 324464 3992 324470 4004
rect 357526 3992 357532 4004
rect 324464 3964 357532 3992
rect 324464 3952 324470 3964
rect 357526 3952 357532 3964
rect 357584 3952 357590 4004
rect 215202 3884 215208 3936
rect 215260 3924 215266 3936
rect 262950 3924 262956 3936
rect 215260 3896 262956 3924
rect 215260 3884 215266 3896
rect 262950 3884 262956 3896
rect 263008 3884 263014 3936
rect 329190 3884 329196 3936
rect 329248 3924 329254 3936
rect 361850 3924 361856 3936
rect 329248 3896 361856 3924
rect 329248 3884 329254 3896
rect 361850 3884 361856 3896
rect 361908 3884 361914 3936
rect 4062 3816 4068 3868
rect 4120 3856 4126 3868
rect 7558 3856 7564 3868
rect 4120 3828 7564 3856
rect 4120 3816 4126 3828
rect 7558 3816 7564 3828
rect 7616 3816 7622 3868
rect 213730 3816 213736 3868
rect 213788 3856 213794 3868
rect 268838 3856 268844 3868
rect 213788 3828 268844 3856
rect 213788 3816 213794 3828
rect 268838 3816 268844 3828
rect 268896 3816 268902 3868
rect 325602 3816 325608 3868
rect 325660 3856 325666 3868
rect 358998 3856 359004 3868
rect 325660 3828 359004 3856
rect 325660 3816 325666 3828
rect 358998 3816 359004 3828
rect 359056 3816 359062 3868
rect 69106 3748 69112 3800
rect 69164 3788 69170 3800
rect 71038 3788 71044 3800
rect 69164 3760 71044 3788
rect 69164 3748 69170 3760
rect 71038 3748 71044 3760
rect 71096 3748 71102 3800
rect 135254 3748 135260 3800
rect 135312 3788 135318 3800
rect 136450 3788 136456 3800
rect 135312 3760 136456 3788
rect 135312 3748 135318 3760
rect 136450 3748 136456 3760
rect 136508 3748 136514 3800
rect 170766 3748 170772 3800
rect 170824 3788 170830 3800
rect 174538 3788 174544 3800
rect 170824 3760 174544 3788
rect 170824 3748 170830 3760
rect 174538 3748 174544 3760
rect 174596 3748 174602 3800
rect 212442 3748 212448 3800
rect 212500 3788 212506 3800
rect 271230 3788 271236 3800
rect 212500 3760 271236 3788
rect 212500 3748 212506 3760
rect 271230 3748 271236 3760
rect 271288 3748 271294 3800
rect 309042 3748 309048 3800
rect 309100 3788 309106 3800
rect 356698 3788 356704 3800
rect 309100 3760 356704 3788
rect 309100 3748 309106 3760
rect 356698 3748 356704 3760
rect 356756 3748 356762 3800
rect 357342 3748 357348 3800
rect 357400 3788 357406 3800
rect 362034 3788 362040 3800
rect 357400 3760 362040 3788
rect 357400 3748 357406 3760
rect 362034 3748 362040 3760
rect 362092 3748 362098 3800
rect 25314 3680 25320 3732
rect 25372 3720 25378 3732
rect 171870 3720 171876 3732
rect 25372 3692 171876 3720
rect 25372 3680 25378 3692
rect 171870 3680 171876 3692
rect 171928 3680 171934 3732
rect 217962 3680 217968 3732
rect 218020 3720 218026 3732
rect 278314 3720 278320 3732
rect 218020 3692 278320 3720
rect 218020 3680 218026 3692
rect 278314 3680 278320 3692
rect 278372 3680 278378 3732
rect 294874 3680 294880 3732
rect 294932 3720 294938 3732
rect 348510 3720 348516 3732
rect 294932 3692 348516 3720
rect 294932 3680 294938 3692
rect 348510 3680 348516 3692
rect 348568 3680 348574 3732
rect 349246 3680 349252 3732
rect 349304 3720 349310 3732
rect 357618 3720 357624 3732
rect 349304 3692 357624 3720
rect 349304 3680 349310 3692
rect 357618 3680 357624 3692
rect 357676 3680 357682 3732
rect 14458 3652 14464 3664
rect 6886 3624 14464 3652
rect 1670 3544 1676 3596
rect 1728 3584 1734 3596
rect 6886 3584 6914 3624
rect 14458 3612 14464 3624
rect 14516 3612 14522 3664
rect 14734 3612 14740 3664
rect 14792 3652 14798 3664
rect 25590 3652 25596 3664
rect 14792 3624 25596 3652
rect 14792 3612 14798 3624
rect 25590 3612 25596 3624
rect 25648 3612 25654 3664
rect 33594 3612 33600 3664
rect 33652 3652 33658 3664
rect 39390 3652 39396 3664
rect 33652 3624 39396 3652
rect 33652 3612 33658 3624
rect 39390 3612 39396 3624
rect 39448 3612 39454 3664
rect 52546 3612 52552 3664
rect 52604 3652 52610 3664
rect 204898 3652 204904 3664
rect 52604 3624 204904 3652
rect 52604 3612 52610 3624
rect 204898 3612 204904 3624
rect 204956 3612 204962 3664
rect 212258 3612 212264 3664
rect 212316 3652 212322 3664
rect 272426 3652 272432 3664
rect 212316 3624 272432 3652
rect 212316 3612 212322 3624
rect 272426 3612 272432 3624
rect 272484 3612 272490 3664
rect 291378 3612 291384 3664
rect 291436 3652 291442 3664
rect 348418 3652 348424 3664
rect 291436 3624 348424 3652
rect 291436 3612 291442 3624
rect 348418 3612 348424 3624
rect 348476 3612 348482 3664
rect 350442 3612 350448 3664
rect 350500 3652 350506 3664
rect 361942 3652 361948 3664
rect 350500 3624 361948 3652
rect 350500 3612 350506 3624
rect 361942 3612 361948 3624
rect 362000 3612 362006 3664
rect 1728 3556 6914 3584
rect 1728 3544 1734 3556
rect 12342 3544 12348 3596
rect 12400 3584 12406 3596
rect 13078 3584 13084 3596
rect 12400 3556 13084 3584
rect 12400 3544 12406 3556
rect 13078 3544 13084 3556
rect 13136 3544 13142 3596
rect 15930 3544 15936 3596
rect 15988 3584 15994 3596
rect 170398 3584 170404 3596
rect 15988 3556 170404 3584
rect 15988 3544 15994 3556
rect 170398 3544 170404 3556
rect 170456 3544 170462 3596
rect 193214 3544 193220 3596
rect 193272 3584 193278 3596
rect 194410 3584 194416 3596
rect 193272 3556 194416 3584
rect 193272 3544 193278 3556
rect 194410 3544 194416 3556
rect 194468 3544 194474 3596
rect 215018 3544 215024 3596
rect 215076 3584 215082 3596
rect 274818 3584 274824 3596
rect 215076 3556 274824 3584
rect 215076 3544 215082 3556
rect 274818 3544 274824 3556
rect 274876 3544 274882 3596
rect 292574 3544 292580 3596
rect 292632 3584 292638 3596
rect 293310 3584 293316 3596
rect 292632 3556 293316 3584
rect 292632 3544 292638 3556
rect 293310 3544 293316 3556
rect 293368 3544 293374 3596
rect 296070 3544 296076 3596
rect 296128 3584 296134 3596
rect 353938 3584 353944 3596
rect 296128 3556 353944 3584
rect 296128 3544 296134 3556
rect 353938 3544 353944 3556
rect 353996 3544 354002 3596
rect 357526 3544 357532 3596
rect 357584 3584 357590 3596
rect 369302 3584 369308 3596
rect 357584 3556 369308 3584
rect 357584 3544 357590 3556
rect 369302 3544 369308 3556
rect 369360 3544 369366 3596
rect 413278 3544 413284 3596
rect 413336 3584 413342 3596
rect 426158 3584 426164 3596
rect 413336 3556 426164 3584
rect 413336 3544 413342 3556
rect 426158 3544 426164 3556
rect 426216 3544 426222 3596
rect 475378 3544 475384 3596
rect 475436 3584 475442 3596
rect 476942 3584 476948 3596
rect 475436 3556 476948 3584
rect 475436 3544 475442 3556
rect 476942 3544 476948 3556
rect 477000 3544 477006 3596
rect 496078 3544 496084 3596
rect 496136 3584 496142 3596
rect 497090 3584 497096 3596
rect 496136 3556 497096 3584
rect 496136 3544 496142 3556
rect 497090 3544 497096 3556
rect 497148 3544 497154 3596
rect 498194 3544 498200 3596
rect 498252 3584 498258 3596
rect 499022 3584 499028 3596
rect 498252 3556 499028 3584
rect 498252 3544 498258 3556
rect 499022 3544 499028 3556
rect 499080 3544 499086 3596
rect 504358 3544 504364 3596
rect 504416 3584 504422 3596
rect 507670 3584 507676 3596
rect 504416 3556 507676 3584
rect 504416 3544 504422 3556
rect 507670 3544 507676 3556
rect 507728 3544 507734 3596
rect 511258 3544 511264 3596
rect 511316 3584 511322 3596
rect 513558 3584 513564 3596
rect 511316 3556 513564 3584
rect 511316 3544 511322 3556
rect 513558 3544 513564 3556
rect 513616 3544 513622 3596
rect 514018 3544 514024 3596
rect 514076 3584 514082 3596
rect 514754 3584 514760 3596
rect 514076 3556 514760 3584
rect 514076 3544 514082 3556
rect 514754 3544 514760 3556
rect 514812 3544 514818 3596
rect 538858 3544 538864 3596
rect 538916 3584 538922 3596
rect 551462 3584 551468 3596
rect 538916 3556 551468 3584
rect 538916 3544 538922 3556
rect 551462 3544 551468 3556
rect 551520 3544 551526 3596
rect 564434 3544 564440 3596
rect 564492 3584 564498 3596
rect 565262 3584 565268 3596
rect 564492 3556 565268 3584
rect 564492 3544 564498 3556
rect 565262 3544 565268 3556
rect 565320 3544 565326 3596
rect 6454 3476 6460 3528
rect 6512 3516 6518 3528
rect 172054 3516 172060 3528
rect 6512 3488 172060 3516
rect 6512 3476 6518 3488
rect 172054 3476 172060 3488
rect 172112 3476 172118 3528
rect 217318 3476 217324 3528
rect 217376 3516 217382 3528
rect 281902 3516 281908 3528
rect 217376 3488 281908 3516
rect 217376 3476 217382 3488
rect 281902 3476 281908 3488
rect 281960 3476 281966 3528
rect 299658 3476 299664 3528
rect 299716 3516 299722 3528
rect 357342 3516 357348 3528
rect 299716 3488 357348 3516
rect 299716 3476 299722 3488
rect 357342 3476 357348 3488
rect 357400 3476 357406 3528
rect 357434 3476 357440 3528
rect 357492 3516 357498 3528
rect 358722 3516 358728 3528
rect 357492 3488 358728 3516
rect 357492 3476 357498 3488
rect 358722 3476 358728 3488
rect 358780 3476 358786 3528
rect 373994 3476 374000 3528
rect 374052 3516 374058 3528
rect 375282 3516 375288 3528
rect 374052 3488 375288 3516
rect 374052 3476 374058 3488
rect 375282 3476 375288 3488
rect 375340 3476 375346 3528
rect 390554 3476 390560 3528
rect 390612 3516 390618 3528
rect 391842 3516 391848 3528
rect 390612 3488 391848 3516
rect 390612 3476 390618 3488
rect 391842 3476 391848 3488
rect 391900 3476 391906 3528
rect 415486 3476 415492 3528
rect 415544 3516 415550 3528
rect 416682 3516 416688 3528
rect 415544 3488 416688 3516
rect 415544 3476 415550 3488
rect 416682 3476 416688 3488
rect 416740 3476 416746 3528
rect 422938 3476 422944 3528
rect 422996 3516 423002 3528
rect 424962 3516 424968 3528
rect 422996 3488 424968 3516
rect 422996 3476 423002 3488
rect 424962 3476 424968 3488
rect 425020 3476 425026 3528
rect 428550 3476 428556 3528
rect 428608 3516 428614 3528
rect 429654 3516 429660 3528
rect 428608 3488 429660 3516
rect 428608 3476 428614 3488
rect 429654 3476 429660 3488
rect 429712 3476 429718 3528
rect 431954 3476 431960 3528
rect 432012 3516 432018 3528
rect 433242 3516 433248 3528
rect 432012 3488 433248 3516
rect 432012 3476 432018 3488
rect 433242 3476 433248 3488
rect 433300 3476 433306 3528
rect 440326 3476 440332 3528
rect 440384 3516 440390 3528
rect 441522 3516 441528 3528
rect 440384 3488 441528 3516
rect 440384 3476 440390 3488
rect 441522 3476 441528 3488
rect 441580 3476 441586 3528
rect 448606 3476 448612 3528
rect 448664 3516 448670 3528
rect 449802 3516 449808 3528
rect 448664 3488 449808 3516
rect 448664 3476 448670 3488
rect 449802 3476 449808 3488
rect 449860 3476 449866 3528
rect 465074 3476 465080 3528
rect 465132 3516 465138 3528
rect 465902 3516 465908 3528
rect 465132 3488 465908 3516
rect 465132 3476 465138 3488
rect 465902 3476 465908 3488
rect 465960 3476 465966 3528
rect 471238 3476 471244 3528
rect 471296 3516 471302 3528
rect 473446 3516 473452 3528
rect 471296 3488 473452 3516
rect 471296 3476 471302 3488
rect 473446 3476 473452 3488
rect 473504 3476 473510 3528
rect 480898 3476 480904 3528
rect 480956 3516 480962 3528
rect 580994 3516 581000 3528
rect 480956 3488 581000 3516
rect 480956 3476 480962 3488
rect 580994 3476 581000 3488
rect 581052 3476 581058 3528
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 171778 3448 171784 3460
rect 624 3420 171784 3448
rect 624 3408 630 3420
rect 171778 3408 171784 3420
rect 171836 3408 171842 3460
rect 173158 3408 173164 3460
rect 173216 3448 173222 3460
rect 184198 3448 184204 3460
rect 173216 3420 184204 3448
rect 173216 3408 173222 3420
rect 184198 3408 184204 3420
rect 184256 3408 184262 3460
rect 219158 3408 219164 3460
rect 219216 3448 219222 3460
rect 287790 3448 287796 3460
rect 219216 3420 287796 3448
rect 219216 3408 219222 3420
rect 287790 3408 287796 3420
rect 287848 3408 287854 3460
rect 288986 3408 288992 3460
rect 289044 3448 289050 3460
rect 354122 3448 354128 3460
rect 289044 3420 354128 3448
rect 289044 3408 289050 3420
rect 354122 3408 354128 3420
rect 354180 3408 354186 3460
rect 356330 3408 356336 3460
rect 356388 3448 356394 3460
rect 369854 3448 369860 3460
rect 356388 3420 369860 3448
rect 356388 3408 356394 3420
rect 369854 3408 369860 3420
rect 369912 3408 369918 3460
rect 378778 3408 378784 3460
rect 378836 3448 378842 3460
rect 572714 3448 572720 3460
rect 378836 3420 572720 3448
rect 378836 3408 378842 3420
rect 572714 3408 572720 3420
rect 572772 3408 572778 3460
rect 38378 3340 38384 3392
rect 38436 3380 38442 3392
rect 39298 3380 39304 3392
rect 38436 3352 39304 3380
rect 38436 3340 38442 3352
rect 39298 3340 39304 3352
rect 39356 3340 39362 3392
rect 93854 3340 93860 3392
rect 93912 3380 93918 3392
rect 94774 3380 94780 3392
rect 93912 3352 94780 3380
rect 93912 3340 93918 3352
rect 94774 3340 94780 3352
rect 94832 3340 94838 3392
rect 110414 3340 110420 3392
rect 110472 3380 110478 3392
rect 111610 3380 111616 3392
rect 110472 3352 111616 3380
rect 110472 3340 110478 3352
rect 111610 3340 111616 3352
rect 111668 3340 111674 3392
rect 213638 3340 213644 3392
rect 213696 3380 213702 3392
rect 258258 3380 258264 3392
rect 213696 3352 258264 3380
rect 213696 3340 213702 3352
rect 258258 3340 258264 3352
rect 258316 3340 258322 3392
rect 331582 3340 331588 3392
rect 331640 3380 331646 3392
rect 358906 3380 358912 3392
rect 331640 3352 358912 3380
rect 331640 3340 331646 3352
rect 358906 3340 358912 3352
rect 358964 3340 358970 3392
rect 171962 3272 171968 3324
rect 172020 3312 172026 3324
rect 175918 3312 175924 3324
rect 172020 3284 175924 3312
rect 172020 3272 172026 3284
rect 175918 3272 175924 3284
rect 175976 3272 175982 3324
rect 212074 3272 212080 3324
rect 212132 3312 212138 3324
rect 254670 3312 254676 3324
rect 212132 3284 254676 3312
rect 212132 3272 212138 3284
rect 254670 3272 254676 3284
rect 254728 3272 254734 3324
rect 336274 3272 336280 3324
rect 336332 3312 336338 3324
rect 356146 3312 356152 3324
rect 336332 3284 356152 3312
rect 336332 3272 336338 3284
rect 356146 3272 356152 3284
rect 356204 3272 356210 3324
rect 212350 3204 212356 3256
rect 212408 3244 212414 3256
rect 245194 3244 245200 3256
rect 212408 3216 245200 3244
rect 212408 3204 212414 3216
rect 245194 3204 245200 3216
rect 245252 3204 245258 3256
rect 335078 3204 335084 3256
rect 335136 3244 335142 3256
rect 359274 3244 359280 3256
rect 335136 3216 359280 3244
rect 335136 3204 335142 3216
rect 359274 3204 359280 3216
rect 359332 3204 359338 3256
rect 567838 3204 567844 3256
rect 567896 3244 567902 3256
rect 571518 3244 571524 3256
rect 567896 3216 571524 3244
rect 567896 3204 567902 3216
rect 571518 3204 571524 3216
rect 571576 3204 571582 3256
rect 354030 3136 354036 3188
rect 354088 3176 354094 3188
rect 360930 3176 360936 3188
rect 354088 3148 360936 3176
rect 354088 3136 354094 3148
rect 360930 3136 360936 3148
rect 360988 3136 360994 3188
rect 356146 3068 356152 3120
rect 356204 3108 356210 3120
rect 361666 3108 361672 3120
rect 356204 3080 361672 3108
rect 356204 3068 356210 3080
rect 361666 3068 361672 3080
rect 361724 3068 361730 3120
rect 476758 3068 476764 3120
rect 476816 3108 476822 3120
rect 479334 3108 479340 3120
rect 476816 3080 479340 3108
rect 476816 3068 476822 3080
rect 479334 3068 479340 3080
rect 479392 3068 479398 3120
rect 30098 3000 30104 3052
rect 30156 3040 30162 3052
rect 32398 3040 32404 3052
rect 30156 3012 32404 3040
rect 30156 3000 30162 3012
rect 32398 3000 32404 3012
rect 32456 3000 32462 3052
rect 355226 3000 355232 3052
rect 355284 3040 355290 3052
rect 362218 3040 362224 3052
rect 355284 3012 362224 3040
rect 355284 3000 355290 3012
rect 362218 3000 362224 3012
rect 362276 3000 362282 3052
rect 467650 3000 467656 3052
rect 467708 3040 467714 3052
rect 471054 3040 471060 3052
rect 467708 3012 471060 3040
rect 467708 3000 467714 3012
rect 471054 3000 471060 3012
rect 471112 3000 471118 3052
rect 571978 3000 571984 3052
rect 572036 3040 572042 3052
rect 573910 3040 573916 3052
rect 572036 3012 573916 3040
rect 572036 3000 572042 3012
rect 573910 3000 573916 3012
rect 573968 3000 573974 3052
rect 20622 2864 20628 2916
rect 20680 2904 20686 2916
rect 22738 2904 22744 2916
rect 20680 2876 22744 2904
rect 20680 2864 20686 2876
rect 22738 2864 22744 2876
rect 22796 2864 22802 2916
rect 398834 2184 398840 2236
rect 398892 2224 398898 2236
rect 400122 2224 400128 2236
rect 398892 2196 400128 2224
rect 398892 2184 398898 2196
rect 400122 2184 400128 2196
rect 400180 2184 400186 2236
rect 407114 2184 407120 2236
rect 407172 2224 407178 2236
rect 408402 2224 408408 2236
rect 407172 2196 408408 2224
rect 407172 2184 407178 2196
rect 408402 2184 408408 2196
rect 408460 2184 408466 2236
rect 456794 2184 456800 2236
rect 456852 2224 456858 2236
rect 458082 2224 458088 2236
rect 456852 2196 458088 2224
rect 456852 2184 456858 2196
rect 458082 2184 458088 2196
rect 458140 2184 458146 2236
rect 382274 1912 382280 1964
rect 382332 1952 382338 1964
rect 383562 1952 383568 1964
rect 382332 1924 383568 1952
rect 382332 1912 382338 1924
rect 383562 1912 383568 1924
rect 383620 1912 383626 1964
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 219348 700408 219400 700460
rect 267648 700408 267700 700460
rect 8116 700340 8168 700392
rect 13084 700340 13136 700392
rect 137836 700340 137888 700392
rect 138664 700340 138716 700392
rect 217968 700340 218020 700392
rect 283840 700340 283892 700392
rect 348792 700340 348844 700392
rect 357440 700340 357492 700392
rect 105452 700272 105504 700324
rect 206284 700272 206336 700324
rect 219256 700272 219308 700324
rect 300124 700272 300176 700324
rect 332508 700272 332560 700324
rect 358820 700272 358872 700324
rect 367744 700272 367796 700324
rect 559656 700272 559708 700324
rect 24308 699660 24360 699712
rect 25504 699660 25556 699712
rect 396724 699660 396776 699712
rect 397460 699660 397512 699712
rect 428464 699660 428516 699712
rect 429844 699660 429896 699712
rect 371884 696940 371936 696992
rect 580172 696940 580224 696992
rect 3424 683136 3476 683188
rect 10324 683136 10376 683188
rect 3516 670692 3568 670744
rect 180064 670692 180116 670744
rect 360844 670692 360896 670744
rect 580172 670692 580224 670744
rect 3424 656888 3476 656940
rect 14464 656888 14516 656940
rect 369124 643084 369176 643136
rect 580172 643084 580224 643136
rect 3424 632068 3476 632120
rect 8944 632068 8996 632120
rect 377404 630640 377456 630692
rect 579988 630640 580040 630692
rect 3148 618264 3200 618316
rect 182824 618264 182876 618316
rect 432604 616836 432656 616888
rect 580172 616836 580224 616888
rect 3424 606024 3476 606076
rect 7564 606024 7616 606076
rect 363604 590656 363656 590708
rect 580172 590656 580224 590708
rect 3332 579640 3384 579692
rect 32404 579640 32456 579692
rect 373264 576852 373316 576904
rect 580172 576852 580224 576904
rect 3424 565836 3476 565888
rect 21364 565836 21416 565888
rect 217876 565088 217928 565140
rect 234620 565088 234672 565140
rect 359464 563048 359516 563100
rect 580172 563048 580224 563100
rect 3424 553392 3476 553444
rect 17224 553392 17276 553444
rect 576124 536800 576176 536852
rect 579896 536800 579948 536852
rect 2780 527144 2832 527196
rect 4804 527144 4856 527196
rect 570604 524424 570656 524476
rect 580172 524424 580224 524476
rect 3056 500964 3108 501016
rect 18604 500964 18656 501016
rect 574744 484372 574796 484424
rect 580172 484372 580224 484424
rect 219256 478524 219308 478576
rect 266452 478524 266504 478576
rect 217968 478456 218020 478508
rect 267740 478456 267792 478508
rect 217416 478388 217468 478440
rect 302240 478388 302292 478440
rect 266360 478320 266412 478372
rect 357440 478320 357492 478372
rect 218888 478252 218940 478304
rect 310520 478252 310572 478304
rect 264980 478184 265032 478236
rect 358820 478184 358872 478236
rect 18604 478116 18656 478168
rect 281540 478116 281592 478168
rect 241428 476756 241480 476808
rect 309140 476756 309192 476808
rect 242808 476688 242860 476740
rect 311900 476688 311952 476740
rect 238484 476620 238536 476672
rect 305000 476620 305052 476672
rect 306104 476620 306156 476672
rect 322204 476620 322256 476672
rect 264888 476552 264940 476604
rect 317420 476552 317472 476604
rect 269028 476484 269080 476536
rect 321560 476484 321612 476536
rect 259368 476416 259420 476468
rect 314660 476416 314712 476468
rect 253848 476348 253900 476400
rect 309232 476348 309284 476400
rect 318708 476348 318760 476400
rect 327724 476348 327776 476400
rect 303528 476280 303580 476332
rect 320824 476280 320876 476332
rect 321468 476280 321520 476332
rect 329104 476280 329156 476332
rect 309048 476212 309100 476264
rect 323584 476212 323636 476264
rect 324228 476212 324280 476264
rect 338764 476212 338816 476264
rect 240048 476144 240100 476196
rect 307760 476144 307812 476196
rect 311808 476076 311860 476128
rect 324964 476076 325016 476128
rect 326988 476076 327040 476128
rect 331864 476076 331916 476128
rect 302148 475532 302200 475584
rect 336740 475532 336792 475584
rect 281448 475464 281500 475516
rect 327080 475464 327132 475516
rect 237288 475396 237340 475448
rect 305092 475396 305144 475448
rect 217600 475328 217652 475380
rect 316132 475328 316184 475380
rect 3424 474716 3476 474768
rect 282920 474716 282972 474768
rect 274548 474172 274600 474224
rect 324320 474172 324372 474224
rect 237380 474104 237432 474156
rect 303620 474104 303672 474156
rect 255228 474036 255280 474088
rect 323032 474036 323084 474088
rect 17224 473968 17276 474020
rect 280160 473968 280212 474020
rect 314568 473968 314620 474020
rect 343640 473968 343692 474020
rect 252376 472744 252428 472796
rect 318800 472744 318852 472796
rect 218980 472676 219032 472728
rect 307852 472676 307904 472728
rect 315948 472676 316000 472728
rect 345204 472676 345256 472728
rect 255320 472608 255372 472660
rect 373264 472608 373316 472660
rect 217508 471316 217560 471368
rect 300860 471316 300912 471368
rect 3516 471248 3568 471300
rect 283012 471248 283064 471300
rect 284208 471248 284260 471300
rect 328460 471248 328512 471300
rect 251824 470568 251876 470620
rect 580172 470568 580224 470620
rect 274456 469956 274508 470008
rect 342352 469956 342404 470008
rect 219072 469888 219124 469940
rect 313280 469888 313332 469940
rect 25504 469820 25556 469872
rect 274640 469820 274692 469872
rect 299388 469820 299440 469872
rect 335360 469820 335412 469872
rect 218060 468596 218112 468648
rect 269304 468596 269356 468648
rect 271696 468596 271748 468648
rect 289084 468596 289136 468648
rect 291108 468596 291160 468648
rect 332600 468596 332652 468648
rect 217692 468528 217744 468580
rect 318892 468528 318944 468580
rect 263600 468460 263652 468512
rect 396724 468460 396776 468512
rect 270408 467236 270460 467288
rect 339592 467236 339644 467288
rect 21364 467168 21416 467220
rect 280252 467168 280304 467220
rect 252560 467100 252612 467152
rect 576124 467100 576176 467152
rect 266176 465876 266228 465928
rect 297364 465876 297416 465928
rect 217784 465808 217836 465860
rect 320364 465808 320416 465860
rect 88340 465740 88392 465792
rect 273260 465740 273312 465792
rect 259460 465672 259512 465724
rect 527180 465672 527232 465724
rect 267556 464448 267608 464500
rect 335452 464448 335504 464500
rect 180064 464380 180116 464432
rect 277400 464380 277452 464432
rect 251180 464312 251232 464364
rect 574744 464312 574796 464364
rect 259276 462952 259328 463004
rect 327172 462952 327224 463004
rect 3240 462340 3292 462392
rect 284484 462340 284536 462392
rect 256516 461796 256568 461848
rect 311992 461796 312044 461848
rect 278596 461728 278648 461780
rect 347780 461728 347832 461780
rect 4804 461660 4856 461712
rect 281632 461660 281684 461712
rect 258080 461592 258132 461644
rect 580264 461592 580316 461644
rect 250996 460368 251048 460420
rect 306380 460368 306432 460420
rect 277216 460300 277268 460352
rect 346492 460300 346544 460352
rect 256700 460232 256752 460284
rect 377404 460232 377456 460284
rect 32404 460164 32456 460216
rect 278780 460164 278832 460216
rect 262036 459008 262088 459060
rect 298744 459008 298796 459060
rect 273168 458940 273220 458992
rect 341064 458940 341116 458992
rect 8944 458872 8996 458924
rect 277492 458872 277544 458924
rect 253940 458804 253992 458856
rect 570604 458804 570656 458856
rect 260656 457512 260708 457564
rect 328552 457512 328604 457564
rect 153200 457444 153252 457496
rect 271880 457444 271932 457496
rect 249800 456764 249852 456816
rect 580172 456764 580224 456816
rect 251088 456152 251140 456204
rect 317512 456152 317564 456204
rect 262220 456084 262272 456136
rect 462320 456084 462372 456136
rect 10324 456016 10376 456068
rect 276020 456016 276072 456068
rect 280068 456016 280120 456068
rect 349252 456016 349304 456068
rect 252468 454792 252520 454844
rect 320272 454792 320324 454844
rect 256792 454724 256844 454776
rect 369124 454724 369176 454776
rect 40040 454656 40092 454708
rect 274732 454656 274784 454708
rect 275928 454656 275980 454708
rect 345112 454656 345164 454708
rect 249064 453432 249116 453484
rect 305184 453432 305236 453484
rect 169760 453364 169812 453416
rect 270500 453364 270552 453416
rect 271788 453364 271840 453416
rect 340972 453364 341024 453416
rect 254032 453296 254084 453348
rect 363604 453296 363656 453348
rect 246304 452004 246356 452056
rect 309324 452004 309376 452056
rect 265072 451936 265124 451988
rect 364340 451936 364392 451988
rect 7564 451868 7616 451920
rect 278872 451868 278924 451920
rect 288348 451868 288400 451920
rect 331220 451868 331272 451920
rect 253756 450712 253808 450764
rect 321652 450712 321704 450764
rect 217324 450644 217376 450696
rect 302332 450644 302384 450696
rect 263692 450576 263744 450628
rect 428464 450576 428516 450628
rect 13084 450508 13136 450560
rect 274824 450508 274876 450560
rect 293868 449284 293920 449336
rect 333980 449284 334032 449336
rect 247684 449216 247736 449268
rect 310612 449216 310664 449268
rect 258172 449148 258224 449200
rect 371884 449148 371936 449200
rect 3148 448536 3200 448588
rect 284392 448536 284444 448588
rect 256608 447924 256660 447976
rect 324412 447924 324464 447976
rect 71780 447856 71832 447908
rect 273352 447856 273404 447908
rect 296628 447856 296680 447908
rect 335544 447856 335596 447908
rect 260840 447788 260892 447840
rect 494060 447788 494112 447840
rect 260748 446496 260800 446548
rect 330024 446496 330076 446548
rect 259552 446428 259604 446480
rect 367744 446428 367796 446480
rect 138664 446360 138716 446412
rect 270592 446360 270644 446412
rect 206284 445136 206336 445188
rect 271972 445136 272024 445188
rect 257988 445068 258040 445120
rect 325700 445068 325752 445120
rect 258264 445000 258316 445052
rect 360844 445000 360896 445052
rect 201500 443776 201552 443828
rect 269212 443776 269264 443828
rect 278688 443776 278740 443828
rect 325792 443776 325844 443828
rect 219164 443708 219216 443760
rect 314752 443708 314804 443760
rect 255412 443640 255464 443692
rect 432604 443640 432656 443692
rect 277308 442416 277360 442468
rect 325884 442416 325936 442468
rect 249708 442348 249760 442400
rect 314844 442348 314896 442400
rect 182824 442280 182876 442332
rect 278964 442280 279016 442332
rect 254124 442212 254176 442264
rect 359464 442212 359516 442264
rect 248236 440988 248288 441040
rect 314108 440988 314160 441040
rect 14464 440920 14516 440972
rect 277032 440920 277084 440972
rect 286968 440920 287020 440972
rect 330576 440920 330628 440972
rect 252744 440852 252796 440904
rect 578884 440852 578936 440904
rect 245476 439832 245528 439884
rect 306840 439832 306892 439884
rect 266268 439764 266320 439816
rect 334808 439764 334860 439816
rect 264796 439696 264848 439748
rect 333612 439696 333664 439748
rect 263508 439628 263560 439680
rect 332324 439628 332376 439680
rect 268936 439560 268988 439612
rect 338396 439560 338448 439612
rect 267648 439492 267700 439544
rect 337200 439492 337252 439544
rect 338764 439492 338816 439544
rect 348792 439492 348844 439544
rect 244188 438268 244240 438320
rect 304356 438268 304408 438320
rect 262128 438200 262180 438252
rect 331128 438200 331180 438252
rect 274364 438132 274416 438184
rect 344560 438132 344612 438184
rect 264888 437044 264940 437096
rect 219348 436908 219400 436960
rect 267924 436908 267976 436960
rect 258172 436840 258224 436892
rect 258540 436840 258592 436892
rect 273260 436908 273312 436960
rect 273628 436908 273680 436960
rect 274640 436908 274692 436960
rect 275468 436908 275520 436960
rect 278780 436908 278832 436960
rect 279700 436908 279752 436960
rect 281540 436908 281592 436960
rect 282092 436908 282144 436960
rect 282920 436908 282972 436960
rect 283380 436908 283432 436960
rect 311900 436908 311952 436960
rect 312636 436908 312688 436960
rect 317420 436908 317472 436960
rect 317972 436908 318024 436960
rect 318800 436908 318852 436960
rect 319260 436908 319312 436960
rect 320272 436908 320324 436960
rect 321100 436908 321152 436960
rect 325792 436908 325844 436960
rect 326620 436908 326672 436960
rect 327080 436908 327132 436960
rect 327724 436908 327776 436960
rect 328460 436908 328512 436960
rect 329012 436908 329064 436960
rect 345112 436908 345164 436960
rect 345388 436908 345440 436960
rect 412640 436840 412692 436892
rect 254032 436772 254084 436824
rect 254860 436772 254912 436824
rect 256700 436772 256752 436824
rect 257252 436772 257304 436824
rect 258080 436772 258132 436824
rect 259092 436772 259144 436824
rect 259460 436772 259512 436824
rect 260380 436772 260432 436824
rect 268568 436772 268620 436824
rect 477500 436772 477552 436824
rect 263784 436704 263836 436756
rect 542360 436704 542412 436756
rect 231216 436636 231268 436688
rect 286140 436636 286192 436688
rect 325700 436636 325752 436688
rect 325976 436636 326028 436688
rect 210424 436568 210476 436620
rect 295892 436568 295944 436620
rect 203524 436500 203576 436552
rect 295248 436500 295300 436552
rect 198004 436432 198056 436484
rect 297732 436432 297784 436484
rect 244832 436364 244884 436416
rect 353944 436364 353996 436416
rect 244188 436296 244240 436348
rect 355324 436296 355376 436348
rect 88984 436228 89036 436280
rect 300768 436228 300820 436280
rect 14556 436160 14608 436212
rect 291660 436160 291712 436212
rect 8944 436092 8996 436144
rect 292212 436092 292264 436144
rect 263048 435752 263100 435804
rect 268568 435752 268620 435804
rect 261208 435684 261260 435736
rect 263784 435684 263836 435736
rect 98644 435208 98696 435260
rect 289176 435208 289228 435260
rect 225604 435140 225656 435192
rect 291016 435140 291068 435192
rect 207664 435072 207716 435124
rect 298284 435072 298336 435124
rect 246028 435004 246080 435056
rect 356704 435004 356756 435056
rect 100024 434936 100076 434988
rect 287336 434936 287388 434988
rect 7564 434868 7616 434920
rect 285496 434868 285548 434920
rect 285680 434868 285732 434920
rect 580908 434868 580960 434920
rect 282184 434800 282236 434852
rect 580540 434800 580592 434852
rect 241152 434732 241204 434784
rect 577504 434732 577556 434784
rect 309140 434596 309192 434648
rect 310060 434596 310112 434648
rect 335636 434596 335688 434648
rect 336004 434596 336056 434648
rect 263600 434528 263652 434580
rect 263876 434528 263928 434580
rect 264980 434528 265032 434580
rect 265716 434528 265768 434580
rect 302240 434528 302292 434580
rect 302884 434528 302936 434580
rect 305092 434528 305144 434580
rect 305828 434528 305880 434580
rect 309232 434528 309284 434580
rect 309508 434528 309560 434580
rect 335360 434528 335412 434580
rect 336372 434528 336424 434580
rect 243544 434460 243596 434512
rect 352564 434460 352616 434512
rect 327816 434392 327868 434444
rect 346308 434392 346360 434444
rect 329104 434324 329156 434376
rect 347596 434324 347648 434376
rect 331864 434256 331916 434308
rect 349988 434256 350040 434308
rect 94504 434188 94556 434240
rect 290372 434188 290424 434240
rect 324964 434188 325016 434240
rect 342720 434188 342772 434240
rect 246672 434120 246724 434172
rect 285680 434120 285732 434172
rect 298744 434120 298796 434172
rect 316592 434120 316644 434172
rect 322388 434120 322440 434172
rect 340236 434120 340288 434172
rect 238760 434052 238812 434104
rect 282184 434052 282236 434104
rect 297364 434052 297416 434104
rect 320180 434052 320232 434104
rect 320824 434052 320876 434104
rect 339040 434052 339092 434104
rect 217876 433984 217928 434036
rect 269120 433984 269172 434036
rect 240508 433848 240560 433900
rect 279976 433984 280028 434036
rect 289084 433984 289136 434036
rect 323216 433984 323268 434036
rect 323584 433984 323636 434036
rect 341524 433984 341576 434036
rect 269396 433916 269448 433968
rect 287980 433916 288032 433968
rect 248420 433780 248472 433832
rect 289728 433780 289780 433832
rect 242348 433712 242400 433764
rect 282920 433712 282972 433764
rect 229744 433644 229796 433696
rect 286784 433644 286836 433696
rect 231124 433576 231176 433628
rect 288624 433576 288676 433628
rect 209044 433508 209096 433560
rect 292856 433508 292908 433560
rect 199384 433440 199436 433492
rect 294052 433440 294104 433492
rect 350632 433440 350684 433492
rect 480904 433440 480956 433492
rect 247868 433372 247920 433424
rect 262680 433372 262732 433424
rect 351184 433372 351236 433424
rect 581092 433372 581144 433424
rect 249708 433304 249760 433356
rect 272248 433304 272300 433356
rect 280068 433304 280120 433356
rect 289820 433304 289872 433356
rect 304908 433304 304960 433356
rect 305184 433304 305236 433356
rect 351828 433304 351880 433356
rect 582380 433304 582432 433356
rect 289728 432760 289780 432812
rect 580172 432760 580224 432812
rect 3608 432692 3660 432744
rect 269396 432692 269448 432744
rect 279976 432692 280028 432744
rect 3516 432624 3568 432676
rect 280068 432624 280120 432676
rect 282920 432692 282972 432744
rect 580632 432692 580684 432744
rect 580724 432624 580776 432676
rect 3424 432556 3476 432608
rect 253204 432556 253256 432608
rect 262680 432556 262732 432608
rect 580080 432556 580132 432608
rect 97908 432488 97960 432540
rect 251824 432488 251876 432540
rect 206284 432420 206336 432472
rect 293408 432420 293460 432472
rect 200764 432352 200816 432404
rect 297088 432352 297140 432404
rect 196624 432284 196676 432336
rect 301044 432284 301096 432336
rect 140780 432216 140832 432268
rect 249432 432216 249484 432268
rect 352840 432216 352892 432268
rect 247592 432148 247644 432200
rect 352748 432148 352800 432200
rect 242072 432080 242124 432132
rect 358084 432080 358136 432132
rect 245568 432012 245620 432064
rect 352656 432012 352708 432064
rect 233608 431944 233660 431996
rect 580356 431944 580408 431996
rect 272248 431876 272300 431928
rect 579896 431876 579948 431928
rect 250536 431740 250588 431792
rect 355416 430584 355468 430636
rect 580724 427320 580776 427372
rect 579988 427116 580040 427168
rect 580632 427116 580684 427168
rect 580724 427116 580776 427168
rect 3332 423580 3384 423632
rect 7564 423580 7616 423632
rect 355416 419432 355468 419484
rect 579988 419432 580040 419484
rect 3332 411204 3384 411256
rect 229744 411204 229796 411256
rect 352840 405628 352892 405680
rect 579988 405628 580040 405680
rect 3332 398760 3384 398812
rect 231216 398760 231268 398812
rect 3700 375980 3752 376032
rect 231124 375980 231176 376032
rect 167644 374892 167696 374944
rect 174636 374892 174688 374944
rect 121276 374824 121328 374876
rect 170772 374824 170824 374876
rect 108396 374756 108448 374808
rect 229744 374756 229796 374808
rect 131580 374688 131632 374740
rect 171876 374688 171928 374740
rect 147036 374620 147088 374672
rect 170404 374620 170456 374672
rect 139308 374552 139360 374604
rect 170864 374552 170916 374604
rect 116124 374484 116176 374536
rect 173256 374484 173308 374536
rect 110972 374416 111024 374468
rect 170956 374416 171008 374468
rect 165528 374348 165580 374400
rect 226984 374348 227036 374400
rect 162492 374280 162544 374332
rect 228364 374280 228416 374332
rect 157340 374212 157392 374264
rect 230020 374212 230072 374264
rect 129004 374144 129056 374196
rect 229836 374144 229888 374196
rect 113548 374076 113600 374128
rect 231216 374076 231268 374128
rect 14464 373056 14516 373108
rect 165068 373056 165120 373108
rect 165528 373056 165580 373108
rect 136732 372988 136784 373040
rect 170680 372988 170732 373040
rect 144460 372920 144512 372972
rect 188344 372920 188396 372972
rect 126428 372852 126480 372904
rect 173164 372852 173216 372904
rect 100668 372784 100720 372836
rect 174544 372784 174596 372836
rect 152188 372716 152240 372768
rect 231124 372716 231176 372768
rect 103244 372648 103296 372700
rect 229928 372648 229980 372700
rect 149612 372580 149664 372632
rect 170588 372580 170640 372632
rect 3332 372512 3384 372564
rect 100024 372512 100076 372564
rect 99840 371764 99892 371816
rect 97724 371492 97776 371544
rect 97816 371424 97868 371476
rect 106096 371560 106148 371612
rect 118332 371560 118384 371612
rect 118976 371560 119028 371612
rect 119068 371560 119120 371612
rect 155040 371696 155092 371748
rect 170036 371696 170088 371748
rect 173440 371628 173492 371680
rect 124128 371560 124180 371612
rect 173348 371560 173400 371612
rect 230112 371492 230164 371544
rect 231308 371424 231360 371476
rect 173624 371356 173676 371408
rect 170036 371288 170088 371340
rect 231400 371288 231452 371340
rect 228456 371220 228508 371272
rect 172336 368500 172388 368552
rect 231584 368500 231636 368552
rect 169944 367888 169996 367940
rect 170496 367888 170548 367940
rect 172336 362924 172388 362976
rect 230204 362924 230256 362976
rect 172428 357416 172480 357468
rect 230296 357416 230348 357468
rect 172428 354696 172480 354748
rect 230388 354696 230440 354748
rect 352748 353200 352800 353252
rect 580172 353200 580224 353252
rect 172428 351908 172480 351960
rect 220084 351908 220136 351960
rect 172428 346400 172480 346452
rect 224224 346400 224276 346452
rect 172428 342252 172480 342304
rect 232228 342252 232280 342304
rect 172428 339464 172480 339516
rect 231676 339464 231728 339516
rect 172428 336744 172480 336796
rect 182824 336744 182876 336796
rect 172428 331236 172480 331288
rect 231768 331236 231820 331288
rect 172428 328448 172480 328500
rect 227076 328448 227128 328500
rect 356704 325592 356756 325644
rect 580172 325592 580224 325644
rect 171324 322940 171376 322992
rect 228548 322940 228600 322992
rect 171508 320152 171560 320204
rect 231032 320152 231084 320204
rect 3332 320084 3384 320136
rect 98644 320084 98696 320136
rect 171508 317432 171560 317484
rect 231952 317432 232004 317484
rect 172428 314644 172480 314696
rect 232136 314644 232188 314696
rect 231860 313216 231912 313268
rect 232044 313216 232096 313268
rect 172428 311856 172480 311908
rect 232044 311856 232096 311908
rect 172336 311244 172388 311296
rect 230940 311244 230992 311296
rect 172244 311176 172296 311228
rect 232228 311176 232280 311228
rect 170864 311108 170916 311160
rect 232320 311108 232372 311160
rect 172152 310700 172204 310752
rect 171968 310632 172020 310684
rect 222292 310632 222344 310684
rect 172060 310564 172112 310616
rect 232228 310564 232280 310616
rect 230204 310428 230256 310480
rect 232320 310496 232372 310548
rect 232596 310496 232648 310548
rect 232964 310496 233016 310548
rect 233148 310564 233200 310616
rect 233700 310564 233752 310616
rect 233516 310428 233568 310480
rect 232228 310360 232280 310412
rect 222292 310292 222344 310344
rect 231860 310292 231912 310344
rect 232136 310292 232188 310344
rect 235172 310292 235224 310344
rect 248328 310292 248380 310344
rect 232044 310224 232096 310276
rect 235908 310224 235960 310276
rect 230388 310156 230440 310208
rect 238208 310156 238260 310208
rect 230940 310088 230992 310140
rect 232044 310088 232096 310140
rect 231768 310020 231820 310072
rect 241060 310020 241112 310072
rect 172428 309952 172480 310004
rect 235540 309952 235592 310004
rect 231676 309612 231728 309664
rect 244740 309612 244792 309664
rect 228548 309544 228600 309596
rect 238944 309544 238996 309596
rect 230296 309476 230348 309528
rect 242072 309476 242124 309528
rect 297180 309476 297232 309528
rect 356796 309544 356848 309596
rect 231584 309408 231636 309460
rect 247776 309408 247828 309460
rect 297364 309408 297416 309460
rect 356704 309408 356756 309460
rect 231032 309340 231084 309392
rect 248512 309340 248564 309392
rect 298652 309340 298704 309392
rect 358820 309340 358872 309392
rect 231952 309272 232004 309324
rect 251364 309272 251416 309324
rect 298284 309272 298336 309324
rect 361580 309272 361632 309324
rect 182824 309204 182876 309256
rect 238392 309204 238444 309256
rect 297916 309204 297968 309256
rect 360292 309204 360344 309256
rect 170496 309136 170548 309188
rect 233976 309136 234028 309188
rect 299204 309136 299256 309188
rect 367100 309136 367152 309188
rect 171784 309068 171836 309120
rect 232412 309068 232464 309120
rect 233700 309068 233752 309120
rect 238024 309068 238076 309120
rect 347228 309068 347280 309120
rect 363604 309068 363656 309120
rect 230112 309000 230164 309052
rect 233424 309000 233476 309052
rect 346860 309000 346912 309052
rect 364616 309000 364668 309052
rect 233148 308932 233200 308984
rect 240876 308932 240928 308984
rect 261208 308932 261260 308984
rect 261484 308932 261536 308984
rect 346492 308932 346544 308984
rect 364984 308932 365036 308984
rect 229836 308864 229888 308916
rect 241428 308864 241480 308916
rect 345020 308864 345072 308916
rect 364340 308864 364392 308916
rect 231400 308796 231452 308848
rect 239128 308796 239180 308848
rect 188344 308728 188396 308780
rect 237656 308728 237708 308780
rect 228456 308660 228508 308712
rect 249064 308796 249116 308848
rect 345388 308796 345440 308848
rect 364524 308796 364576 308848
rect 170588 308592 170640 308644
rect 246948 308728 247000 308780
rect 258080 308728 258132 308780
rect 346124 308728 346176 308780
rect 364892 308728 364944 308780
rect 250904 308660 250956 308712
rect 245660 308592 245712 308644
rect 305184 308660 305236 308712
rect 305460 308660 305512 308712
rect 348240 308660 348292 308712
rect 352472 308660 352524 308712
rect 352748 308660 352800 308712
rect 364708 308660 364760 308712
rect 267648 308592 267700 308644
rect 314660 308592 314712 308644
rect 315856 308592 315908 308644
rect 316224 308592 316276 308644
rect 318248 308592 318300 308644
rect 320364 308592 320416 308644
rect 320640 308592 320692 308644
rect 344744 308592 344796 308644
rect 364432 308592 364484 308644
rect 173164 308524 173216 308576
rect 243728 308524 243780 308576
rect 252284 308524 252336 308576
rect 170680 308388 170732 308440
rect 236644 308456 236696 308508
rect 270224 308524 270276 308576
rect 275284 308524 275336 308576
rect 294604 308524 294656 308576
rect 294788 308524 294840 308576
rect 313280 308524 313332 308576
rect 314200 308524 314252 308576
rect 314752 308524 314804 308576
rect 315212 308524 315264 308576
rect 316132 308524 316184 308576
rect 316500 308524 316552 308576
rect 317512 308524 317564 308576
rect 317972 308524 318024 308576
rect 339408 308524 339460 308576
rect 364800 308524 364852 308576
rect 268660 308456 268712 308508
rect 304448 308456 304500 308508
rect 347136 308456 347188 308508
rect 350724 308456 350776 308508
rect 352472 308456 352524 308508
rect 367376 308456 367428 308508
rect 231124 308388 231176 308440
rect 239588 308388 239640 308440
rect 173348 308320 173400 308372
rect 241612 308320 241664 308372
rect 243544 308184 243596 308236
rect 251824 308184 251876 308236
rect 232044 308116 232096 308168
rect 243452 308116 243504 308168
rect 246856 308116 246908 308168
rect 252744 308116 252796 308168
rect 231860 308048 231912 308100
rect 246396 308048 246448 308100
rect 250536 308048 250588 308100
rect 269212 308388 269264 308440
rect 295984 308388 296036 308440
rect 349896 308388 349948 308440
rect 367284 308388 367336 308440
rect 312360 308320 312412 308372
rect 313188 308320 313240 308372
rect 313648 308320 313700 308372
rect 314016 308320 314068 308372
rect 314844 308320 314896 308372
rect 315304 308320 315356 308372
rect 316408 308320 316460 308372
rect 317052 308320 317104 308372
rect 317420 308320 317472 308372
rect 317696 308320 317748 308372
rect 317880 308320 317932 308372
rect 318340 308320 318392 308372
rect 318800 308320 318852 308372
rect 319260 308320 319312 308372
rect 319444 308320 319496 308372
rect 319904 308320 319956 308372
rect 320548 308320 320600 308372
rect 321100 308320 321152 308372
rect 340972 308320 341024 308372
rect 343364 308320 343416 308372
rect 344376 308320 344428 308372
rect 360936 308320 360988 308372
rect 273168 308252 273220 308304
rect 273720 308252 273772 308304
rect 311900 308252 311952 308304
rect 312636 308252 312688 308304
rect 313372 308252 313424 308304
rect 313924 308252 313976 308304
rect 314936 308252 314988 308304
rect 315120 308252 315172 308304
rect 316316 308252 316368 308304
rect 317236 308252 317288 308304
rect 319168 308252 319220 308304
rect 320180 308252 320232 308304
rect 321284 308252 321336 308304
rect 350540 308252 350592 308304
rect 350908 308252 350960 308304
rect 312084 308184 312136 308236
rect 312544 308184 312596 308236
rect 313556 308184 313608 308236
rect 314568 308184 314620 308236
rect 314752 308184 314804 308236
rect 315488 308184 315540 308236
rect 316040 308184 316092 308236
rect 316500 308184 316552 308236
rect 317420 308184 317472 308236
rect 318524 308184 318576 308236
rect 318800 308184 318852 308236
rect 350724 308184 350776 308236
rect 351276 308184 351328 308236
rect 312176 308116 312228 308168
rect 313004 308116 313056 308168
rect 313372 308116 313424 308168
rect 314384 308116 314436 308168
rect 314936 308116 314988 308168
rect 315672 308116 315724 308168
rect 319168 308116 319220 308168
rect 319720 308116 319772 308168
rect 350908 308116 350960 308168
rect 351828 308116 351880 308168
rect 318984 308048 319036 308100
rect 319536 308048 319588 308100
rect 347872 308048 347924 308100
rect 363512 308252 363564 308304
rect 250720 307980 250772 308032
rect 254676 307980 254728 308032
rect 275284 307980 275336 308032
rect 280344 307980 280396 308032
rect 311256 307980 311308 308032
rect 312636 307980 312688 308032
rect 316132 307980 316184 308032
rect 316868 307980 316920 308032
rect 319076 307980 319128 308032
rect 320088 307980 320140 308032
rect 249064 307912 249116 307964
rect 255964 307912 256016 307964
rect 270592 307912 270644 307964
rect 271144 307912 271196 307964
rect 242808 307844 242860 307896
rect 250996 307844 251048 307896
rect 257436 307844 257488 307896
rect 263416 307844 263468 307896
rect 272524 307844 272576 307896
rect 278596 307912 278648 307964
rect 318616 307912 318668 307964
rect 319536 307912 319588 307964
rect 330024 307912 330076 307964
rect 331864 307912 331916 307964
rect 345756 307912 345808 307964
rect 352748 307912 352800 307964
rect 278320 307844 278372 307896
rect 280896 307844 280948 307896
rect 325792 307844 325844 307896
rect 329012 307844 329064 307896
rect 347504 307844 347556 307896
rect 359648 307844 359700 307896
rect 237380 307776 237432 307828
rect 240692 307776 240744 307828
rect 247040 307776 247092 307828
rect 250444 307776 250496 307828
rect 251824 307776 251876 307828
rect 259092 307776 259144 307828
rect 270040 307776 270092 307828
rect 270500 307776 270552 307828
rect 275376 307776 275428 307828
rect 277400 307776 277452 307828
rect 278136 307776 278188 307828
rect 278780 307776 278832 307828
rect 306932 307776 306984 307828
rect 308680 307776 308732 307828
rect 309048 307776 309100 307828
rect 310060 307776 310112 307828
rect 321836 307776 321888 307828
rect 323676 307776 323728 307828
rect 324136 307776 324188 307828
rect 325148 307776 325200 307828
rect 325240 307776 325292 307828
rect 327816 307776 327868 307828
rect 328368 307776 328420 307828
rect 329380 307776 329432 307828
rect 331220 307776 331272 307828
rect 333428 307776 333480 307828
rect 341616 307776 341668 307828
rect 342444 307776 342496 307828
rect 229744 307708 229796 307760
rect 243912 307708 243964 307760
rect 227076 307640 227128 307692
rect 241244 307640 241296 307692
rect 172428 307572 172480 307624
rect 245844 307572 245896 307624
rect 220084 307504 220136 307556
rect 242716 307504 242768 307556
rect 228364 307436 228416 307488
rect 248696 307436 248748 307488
rect 224224 307368 224276 307420
rect 241796 307368 241848 307420
rect 170404 307300 170456 307352
rect 249156 307300 249208 307352
rect 170496 307232 170548 307284
rect 236828 307232 236880 307284
rect 323308 307232 323360 307284
rect 323492 307232 323544 307284
rect 215208 307164 215260 307216
rect 290464 307164 290516 307216
rect 316684 307164 316736 307216
rect 437480 307164 437532 307216
rect 210976 307096 211028 307148
rect 339960 307096 340012 307148
rect 350632 307096 350684 307148
rect 351644 307096 351696 307148
rect 195980 307028 196032 307080
rect 280528 307028 280580 307080
rect 326252 307028 326304 307080
rect 500960 307028 501012 307080
rect 171876 306960 171928 307012
rect 251548 306960 251600 307012
rect 269396 306960 269448 307012
rect 269672 306960 269724 307012
rect 325884 306960 325936 307012
rect 326160 306960 326212 307012
rect 337108 306960 337160 307012
rect 246028 306892 246080 306944
rect 251456 306756 251508 306808
rect 261392 306824 261444 306876
rect 283196 306824 283248 306876
rect 283656 306824 283708 306876
rect 294052 306824 294104 306876
rect 263876 306688 263928 306740
rect 264152 306688 264204 306740
rect 337200 306756 337252 306808
rect 332692 306688 332744 306740
rect 333060 306688 333112 306740
rect 261392 306620 261444 306672
rect 294052 306620 294104 306672
rect 263876 306552 263928 306604
rect 264060 306552 264112 306604
rect 300860 306552 300912 306604
rect 301320 306552 301372 306604
rect 252744 306484 252796 306536
rect 253664 306484 253716 306536
rect 263600 306484 263652 306536
rect 264612 306484 264664 306536
rect 282736 306484 282788 306536
rect 289084 306484 289136 306536
rect 309140 306484 309192 306536
rect 309600 306484 309652 306536
rect 329932 306484 329984 306536
rect 330576 306484 330628 306536
rect 248604 306416 248656 306468
rect 249524 306416 249576 306468
rect 252652 306416 252704 306468
rect 253296 306416 253348 306468
rect 255596 306416 255648 306468
rect 255872 306416 255924 306468
rect 258172 306416 258224 306468
rect 258724 306416 258776 306468
rect 262220 306416 262272 306468
rect 262864 306416 262916 306468
rect 263784 306416 263836 306468
rect 264796 306416 264848 306468
rect 264980 306416 265032 306468
rect 265440 306416 265492 306468
rect 266636 306416 266688 306468
rect 266912 306416 266964 306468
rect 269764 306416 269816 306468
rect 271604 306416 271656 306468
rect 272064 306416 272116 306468
rect 272156 306416 272208 306468
rect 272800 306416 272852 306468
rect 273260 306416 273312 306468
rect 273628 306416 273680 306468
rect 276204 306416 276256 306468
rect 276480 306416 276532 306468
rect 277492 306416 277544 306468
rect 278412 306416 278464 306468
rect 280528 306416 280580 306468
rect 281448 306416 281500 306468
rect 281724 306416 281776 306468
rect 282184 306416 282236 306468
rect 233332 306348 233384 306400
rect 234160 306348 234212 306400
rect 241704 306348 241756 306400
rect 242624 306348 242676 306400
rect 247132 306348 247184 306400
rect 247960 306348 248012 306400
rect 248696 306348 248748 306400
rect 249340 306348 249392 306400
rect 251272 306348 251324 306400
rect 252376 306348 252428 306400
rect 252560 306348 252612 306400
rect 253204 306348 253256 306400
rect 256700 306348 256752 306400
rect 257344 306348 257396 306400
rect 258356 306348 258408 306400
rect 258908 306348 258960 306400
rect 259552 306348 259604 306400
rect 259828 306348 259880 306400
rect 259920 306348 259972 306400
rect 260564 306348 260616 306400
rect 262404 306348 262456 306400
rect 263048 306348 263100 306400
rect 263692 306348 263744 306400
rect 264152 306348 264204 306400
rect 269304 306348 269356 306400
rect 270868 306348 270920 306400
rect 271328 306348 271380 306400
rect 272340 306348 272392 306400
rect 273076 306348 273128 306400
rect 273536 306348 273588 306400
rect 273812 306348 273864 306400
rect 275008 306348 275060 306400
rect 275468 306348 275520 306400
rect 276020 306348 276072 306400
rect 277216 306348 277268 306400
rect 277676 306348 277728 306400
rect 278044 306348 278096 306400
rect 278872 306348 278924 306400
rect 279516 306348 279568 306400
rect 280436 306348 280488 306400
rect 281264 306348 281316 306400
rect 3332 306280 3384 306332
rect 94504 306280 94556 306332
rect 218980 306280 219032 306332
rect 287428 306416 287480 306468
rect 307852 306416 307904 306468
rect 308496 306416 308548 306468
rect 309324 306416 309376 306468
rect 309784 306416 309836 306468
rect 310520 306416 310572 306468
rect 310888 306416 310940 306468
rect 322940 306416 322992 306468
rect 327172 306416 327224 306468
rect 327448 306416 327500 306468
rect 330116 306416 330168 306468
rect 330392 306416 330444 306468
rect 291384 306348 291436 306400
rect 291752 306348 291804 306400
rect 295340 306348 295392 306400
rect 296352 306348 296404 306400
rect 296720 306348 296772 306400
rect 297180 306348 297232 306400
rect 301136 306348 301188 306400
rect 301320 306348 301372 306400
rect 303988 306348 304040 306400
rect 304816 306348 304868 306400
rect 305000 306348 305052 306400
rect 305552 306348 305604 306400
rect 321836 306348 321888 306400
rect 322572 306348 322624 306400
rect 286048 306280 286100 306332
rect 286784 306280 286836 306332
rect 289912 306280 289964 306332
rect 290372 306280 290424 306332
rect 291476 306280 291528 306332
rect 292396 306280 292448 306332
rect 292856 306280 292908 306332
rect 293316 306280 293368 306332
rect 293960 306280 294012 306332
rect 294236 306280 294288 306332
rect 295524 306280 295576 306332
rect 296168 306280 296220 306332
rect 299480 306280 299532 306332
rect 299756 306280 299808 306332
rect 303896 306280 303948 306332
rect 304264 306280 304316 306332
rect 305092 306280 305144 306332
rect 305736 306280 305788 306332
rect 306380 306280 306432 306332
rect 307116 306280 307168 306332
rect 321652 306280 321704 306332
rect 322112 306280 322164 306332
rect 218888 306212 218940 306264
rect 282736 306212 282788 306264
rect 283012 306212 283064 306264
rect 283932 306212 283984 306264
rect 288900 306212 288952 306264
rect 289452 306212 289504 306264
rect 290188 306212 290240 306264
rect 290832 306212 290884 306264
rect 291568 306212 291620 306264
rect 292120 306212 292172 306264
rect 296720 306212 296772 306264
rect 297088 306212 297140 306264
rect 302516 306212 302568 306264
rect 303068 306212 303120 306264
rect 303712 306212 303764 306264
rect 304172 306212 304224 306264
rect 305276 306212 305328 306264
rect 305920 306212 305972 306264
rect 309508 306212 309560 306264
rect 310152 306212 310204 306264
rect 310704 306212 310756 306264
rect 310980 306212 311032 306264
rect 321560 306212 321612 306264
rect 322756 306212 322808 306264
rect 169944 306144 169996 306196
rect 238392 306144 238444 306196
rect 239036 306144 239088 306196
rect 239496 306144 239548 306196
rect 242992 306144 243044 306196
rect 244096 306144 244148 306196
rect 244556 306144 244608 306196
rect 245108 306144 245160 306196
rect 250076 306144 250128 306196
rect 250628 306144 250680 306196
rect 251548 306144 251600 306196
rect 252192 306144 252244 306196
rect 252836 306144 252888 306196
rect 253848 306144 253900 306196
rect 254032 306144 254084 306196
rect 255044 306144 255096 306196
rect 255688 306144 255740 306196
rect 256424 306144 256476 306196
rect 256976 306144 257028 306196
rect 257712 306144 257764 306196
rect 258264 306144 258316 306196
rect 258632 306144 258684 306196
rect 259460 306144 259512 306196
rect 259828 306144 259880 306196
rect 261300 306144 261352 306196
rect 261944 306144 261996 306196
rect 263692 306144 263744 306196
rect 264244 306144 264296 306196
rect 265072 306144 265124 306196
rect 265716 306144 265768 306196
rect 266728 306144 266780 306196
rect 267096 306144 267148 306196
rect 269488 306144 269540 306196
rect 270132 306144 270184 306196
rect 271972 306144 272024 306196
rect 272984 306144 273036 306196
rect 273812 306144 273864 306196
rect 274548 306144 274600 306196
rect 274640 306144 274692 306196
rect 275100 306144 275152 306196
rect 278044 306144 278096 306196
rect 278320 306144 278372 306196
rect 280252 306144 280304 306196
rect 280712 306144 280764 306196
rect 282092 306144 282144 306196
rect 282552 306144 282604 306196
rect 216404 306076 216456 306128
rect 288532 306144 288584 306196
rect 290280 306144 290332 306196
rect 291016 306144 291068 306196
rect 293132 306144 293184 306196
rect 293684 306144 293736 306196
rect 294236 306144 294288 306196
rect 294880 306144 294932 306196
rect 298100 306144 298152 306196
rect 299388 306144 299440 306196
rect 299572 306144 299624 306196
rect 300216 306144 300268 306196
rect 302332 306144 302384 306196
rect 303436 306144 303488 306196
rect 303620 306144 303672 306196
rect 304632 306144 304684 306196
rect 305368 306144 305420 306196
rect 306104 306144 306156 306196
rect 309416 306144 309468 306196
rect 310336 306144 310388 306196
rect 321744 306144 321796 306196
rect 322204 306144 322256 306196
rect 333520 306416 333572 306468
rect 337016 306416 337068 306468
rect 337292 306416 337344 306468
rect 349712 306416 349764 306468
rect 332784 306348 332836 306400
rect 336832 306348 336884 306400
rect 337660 306348 337712 306400
rect 324504 306280 324556 306332
rect 327080 306280 327132 306332
rect 327724 306280 327776 306332
rect 328460 306280 328512 306332
rect 329104 306280 329156 306332
rect 330024 306280 330076 306332
rect 330852 306280 330904 306332
rect 333244 306280 333296 306332
rect 333704 306280 333756 306332
rect 334348 306280 334400 306332
rect 334624 306280 334676 306332
rect 336740 306280 336792 306332
rect 337292 306280 337344 306332
rect 341156 306280 341208 306332
rect 341708 306280 341760 306332
rect 343640 306280 343692 306332
rect 344192 306280 344244 306332
rect 366272 306280 366324 306332
rect 323308 306212 323360 306264
rect 323768 306212 323820 306264
rect 323400 306144 323452 306196
rect 283196 306076 283248 306128
rect 283748 306076 283800 306128
rect 292948 306076 293000 306128
rect 293868 306076 293920 306128
rect 294144 306076 294196 306128
rect 295248 306076 295300 306128
rect 299480 306076 299532 306128
rect 300768 306076 300820 306128
rect 301228 306076 301280 306128
rect 301964 306076 302016 306128
rect 305000 306076 305052 306128
rect 306288 306076 306340 306128
rect 306564 306076 306616 306128
rect 307668 306076 307720 306128
rect 310704 306076 310756 306128
rect 311532 306076 311584 306128
rect 321652 306076 321704 306128
rect 322388 306076 322440 306128
rect 323032 306076 323084 306128
rect 323584 306076 323636 306128
rect 325976 306212 326028 306264
rect 326620 306212 326672 306264
rect 327540 306212 327592 306264
rect 328092 306212 328144 306264
rect 329840 306212 329892 306264
rect 330392 306212 330444 306264
rect 336924 306212 336976 306264
rect 337752 306212 337804 306264
rect 340972 306212 341024 306264
rect 341892 306212 341944 306264
rect 342352 306212 342404 306264
rect 342904 306212 342956 306264
rect 349160 306212 349212 306264
rect 350172 306212 350224 306264
rect 350356 306212 350408 306264
rect 366364 306212 366416 306264
rect 325884 306144 325936 306196
rect 326436 306144 326488 306196
rect 327264 306144 327316 306196
rect 327908 306144 327960 306196
rect 331680 306144 331732 306196
rect 332508 306144 332560 306196
rect 332968 306144 333020 306196
rect 333336 306144 333388 306196
rect 335268 306144 335320 306196
rect 335636 306144 335688 306196
rect 335820 306144 335872 306196
rect 336372 306144 336424 306196
rect 336740 306144 336792 306196
rect 337936 306144 337988 306196
rect 338120 306144 338172 306196
rect 214932 306008 214984 306060
rect 172244 305940 172296 305992
rect 244924 305940 244976 305992
rect 254308 305940 254360 305992
rect 255228 305940 255280 305992
rect 255412 305940 255464 305992
rect 256332 305940 256384 305992
rect 257160 305940 257212 305992
rect 257896 305940 257948 305992
rect 258264 305940 258316 305992
rect 259276 305940 259328 305992
rect 259644 305940 259696 305992
rect 260380 305940 260432 305992
rect 261116 305940 261168 305992
rect 261760 305940 261812 305992
rect 263968 305940 264020 305992
rect 264428 305940 264480 305992
rect 265256 305940 265308 305992
rect 265900 305940 265952 305992
rect 266360 305940 266412 305992
rect 266820 305940 266872 305992
rect 269396 305940 269448 305992
rect 270316 305940 270368 305992
rect 270960 305940 271012 305992
rect 271512 305940 271564 305992
rect 273444 306008 273496 306060
rect 273996 306008 274048 306060
rect 274824 306008 274876 306060
rect 275560 306008 275612 306060
rect 276388 306008 276440 306060
rect 277032 306008 277084 306060
rect 277768 306008 277820 306060
rect 278228 306008 278280 306060
rect 279148 306008 279200 306060
rect 279700 306008 279752 306060
rect 281816 306008 281868 306060
rect 282368 306008 282420 306060
rect 287980 306008 288032 306060
rect 292764 306008 292816 306060
rect 293500 306008 293552 306060
rect 296812 306008 296864 306060
rect 297732 306008 297784 306060
rect 300860 306008 300912 306060
rect 301872 306008 301924 306060
rect 323216 306008 323268 306060
rect 323952 306008 324004 306060
rect 324596 306076 324648 306128
rect 325424 306076 325476 306128
rect 327356 306076 327408 306128
rect 328184 306076 328236 306128
rect 328828 306076 328880 306128
rect 329472 306076 329524 306128
rect 331496 306076 331548 306128
rect 331956 306076 332008 306128
rect 334440 306076 334492 306128
rect 334992 306076 335044 306128
rect 335452 306076 335504 306128
rect 336188 306076 336240 306128
rect 328920 306008 328972 306060
rect 329288 306008 329340 306060
rect 331404 306008 331456 306060
rect 332140 306008 332192 306060
rect 334164 306008 334216 306060
rect 334808 306008 334860 306060
rect 349988 306144 350040 306196
rect 367560 306144 367612 306196
rect 348976 306076 349028 306128
rect 365904 306076 365956 306128
rect 349344 306008 349396 306060
rect 367744 306008 367796 306060
rect 296904 305940 296956 305992
rect 297548 305940 297600 305992
rect 324412 305940 324464 305992
rect 324504 305940 324556 305992
rect 325608 305940 325660 305992
rect 328552 305940 328604 305992
rect 329012 305940 329064 305992
rect 329932 305940 329984 305992
rect 331036 305940 331088 305992
rect 334256 305940 334308 305992
rect 335176 305940 335228 305992
rect 338212 305940 338264 305992
rect 348608 305940 348660 305992
rect 367652 305940 367704 305992
rect 216312 305872 216364 305924
rect 290648 305872 290700 305924
rect 324228 305872 324280 305924
rect 324872 305872 324924 305924
rect 331772 305872 331824 305924
rect 332324 305872 332376 305924
rect 344008 305872 344060 305924
rect 367468 305872 367520 305924
rect 216588 305804 216640 305856
rect 291200 305804 291252 305856
rect 328552 305804 328604 305856
rect 329656 305804 329708 305856
rect 332784 305804 332836 305856
rect 333888 305804 333940 305856
rect 344560 305804 344612 305856
rect 367836 305804 367888 305856
rect 213828 305736 213880 305788
rect 290096 305736 290148 305788
rect 342628 305736 342680 305788
rect 368572 305736 368624 305788
rect 212080 305668 212132 305720
rect 289636 305668 289688 305720
rect 343088 305668 343140 305720
rect 368848 305668 368900 305720
rect 175924 305600 175976 305652
rect 274640 305600 274692 305652
rect 274916 305600 274968 305652
rect 275928 305600 275980 305652
rect 278964 305600 279016 305652
rect 279424 305600 279476 305652
rect 282000 305600 282052 305652
rect 282828 305600 282880 305652
rect 298192 305600 298244 305652
rect 299020 305600 299072 305652
rect 342076 305600 342128 305652
rect 368940 305600 368992 305652
rect 219072 305532 219124 305584
rect 286416 305532 286468 305584
rect 350908 305532 350960 305584
rect 366180 305532 366232 305584
rect 219164 305464 219216 305516
rect 285312 305464 285364 305516
rect 351000 305464 351052 305516
rect 366088 305464 366140 305516
rect 172612 305396 172664 305448
rect 236276 305396 236328 305448
rect 238944 305396 238996 305448
rect 239956 305396 240008 305448
rect 254216 305396 254268 305448
rect 254584 305396 254636 305448
rect 256792 305396 256844 305448
rect 257252 305396 257304 305448
rect 259460 305396 259512 305448
rect 260012 305396 260064 305448
rect 260932 305396 260984 305448
rect 261576 305396 261628 305448
rect 265348 305396 265400 305448
rect 266176 305396 266228 305448
rect 266636 305396 266688 305448
rect 267280 305396 267332 305448
rect 267832 305396 267884 305448
rect 268292 305396 268344 305448
rect 273720 305396 273772 305448
rect 274180 305396 274232 305448
rect 274640 305396 274692 305448
rect 276848 305396 276900 305448
rect 278964 305396 279016 305448
rect 280068 305396 280120 305448
rect 281724 305396 281776 305448
rect 282644 305396 282696 305448
rect 351460 305396 351512 305448
rect 361028 305396 361080 305448
rect 238668 305328 238720 305380
rect 239772 305328 239824 305380
rect 267740 305328 267792 305380
rect 268200 305328 268252 305380
rect 238392 305260 238444 305312
rect 242256 305260 242308 305312
rect 256792 305260 256844 305312
rect 257528 305260 257580 305312
rect 267832 305260 267884 305312
rect 268844 305260 268896 305312
rect 97172 305192 97224 305244
rect 97540 305192 97592 305244
rect 307944 305192 307996 305244
rect 308772 305192 308824 305244
rect 97540 305056 97592 305108
rect 97816 305056 97868 305108
rect 262496 304988 262548 305040
rect 262864 304988 262916 305040
rect 172336 304920 172388 304972
rect 244280 304920 244332 304972
rect 247224 304920 247276 304972
rect 249708 304920 249760 304972
rect 262312 304920 262364 304972
rect 262772 304920 262824 304972
rect 262496 304852 262548 304904
rect 263508 304852 263560 304904
rect 325700 304852 325752 304904
rect 326804 304852 326856 304904
rect 301412 304648 301464 304700
rect 302148 304648 302200 304700
rect 169852 304444 169904 304496
rect 237840 304444 237892 304496
rect 342444 304444 342496 304496
rect 342720 304444 342772 304496
rect 171692 304376 171744 304428
rect 244372 304376 244424 304428
rect 308128 304376 308180 304428
rect 308956 304376 309008 304428
rect 170036 304308 170088 304360
rect 247592 304308 247644 304360
rect 171876 304240 171928 304292
rect 254860 304240 254912 304292
rect 271052 304240 271104 304292
rect 271696 304240 271748 304292
rect 236092 304172 236144 304224
rect 236276 304172 236328 304224
rect 255780 304104 255832 304156
rect 256148 304104 256200 304156
rect 310612 304104 310664 304156
rect 310888 304104 310940 304156
rect 337108 304104 337160 304156
rect 337476 304104 337528 304156
rect 310612 303968 310664 304020
rect 311440 303968 311492 304020
rect 302424 303696 302476 303748
rect 302884 303696 302936 303748
rect 216128 303560 216180 303612
rect 285956 303560 286008 303612
rect 349252 303560 349304 303612
rect 371332 303560 371384 303612
rect 214748 303492 214800 303544
rect 285496 303492 285548 303544
rect 349804 303492 349856 303544
rect 371608 303492 371660 303544
rect 216496 303424 216548 303476
rect 287152 303424 287204 303476
rect 348424 303424 348476 303476
rect 370504 303424 370556 303476
rect 216220 303356 216272 303408
rect 288164 303356 288216 303408
rect 347688 303356 347740 303408
rect 369124 303356 369176 303408
rect 214840 303288 214892 303340
rect 286600 303288 286652 303340
rect 346676 303288 346728 303340
rect 369952 303288 370004 303340
rect 214656 303220 214708 303272
rect 287612 303220 287664 303272
rect 349528 303220 349580 303272
rect 372988 303220 373040 303272
rect 215024 303152 215076 303204
rect 292304 303152 292356 303204
rect 347320 303152 347372 303204
rect 370688 303152 370740 303204
rect 213460 303084 213512 303136
rect 290464 303084 290516 303136
rect 347044 303084 347096 303136
rect 370596 303084 370648 303136
rect 212448 303016 212500 303068
rect 291844 303016 291896 303068
rect 346308 303016 346360 303068
rect 370136 303016 370188 303068
rect 171968 302948 172020 303000
rect 252008 302948 252060 303000
rect 345940 302948 345992 303000
rect 370044 302948 370096 303000
rect 175280 302880 175332 302932
rect 275376 302880 275428 302932
rect 345572 302880 345624 302932
rect 370228 302880 370280 302932
rect 216036 302812 216088 302864
rect 285680 302812 285732 302864
rect 348792 302812 348844 302864
rect 369216 302812 369268 302864
rect 215116 302744 215168 302796
rect 285128 302744 285180 302796
rect 352012 302744 352064 302796
rect 373080 302744 373132 302796
rect 172336 302676 172388 302728
rect 234804 302676 234856 302728
rect 236460 302676 236512 302728
rect 237288 302676 237340 302728
rect 348056 302676 348108 302728
rect 358176 302676 358228 302728
rect 261024 302472 261076 302524
rect 262128 302472 262180 302524
rect 339960 302268 340012 302320
rect 340604 302268 340656 302320
rect 172428 302132 172480 302184
rect 238668 302132 238720 302184
rect 219348 301588 219400 301640
rect 290280 301588 290332 301640
rect 211988 301520 212040 301572
rect 340420 301520 340472 301572
rect 213368 301452 213420 301504
rect 341064 301452 341116 301504
rect 251364 301316 251416 301368
rect 251640 301316 251692 301368
rect 97448 300772 97500 300824
rect 248880 300772 248932 300824
rect 343732 300772 343784 300824
rect 365076 300772 365128 300824
rect 97264 300704 97316 300756
rect 247040 300704 247092 300756
rect 350540 300704 350592 300756
rect 372712 300704 372764 300756
rect 99380 300636 99432 300688
rect 248604 300636 248656 300688
rect 349160 300636 349212 300688
rect 373264 300636 373316 300688
rect 97724 300568 97776 300620
rect 244556 300568 244608 300620
rect 342628 300568 342680 300620
rect 369308 300568 369360 300620
rect 97816 300500 97868 300552
rect 242808 300500 242860 300552
rect 342444 300500 342496 300552
rect 371424 300500 371476 300552
rect 99012 300432 99064 300484
rect 243084 300432 243136 300484
rect 341156 300432 341208 300484
rect 370320 300432 370372 300484
rect 97632 300364 97684 300416
rect 241980 300364 242032 300416
rect 343640 300364 343692 300416
rect 372804 300364 372856 300416
rect 99472 300296 99524 300348
rect 240600 300296 240652 300348
rect 342536 300296 342588 300348
rect 373172 300296 373224 300348
rect 97356 300228 97408 300280
rect 237380 300228 237432 300280
rect 343364 300228 343416 300280
rect 371792 300228 371844 300280
rect 99840 300160 99892 300212
rect 238944 300160 238996 300212
rect 339684 300160 339736 300212
rect 372896 300160 372948 300212
rect 99196 300092 99248 300144
rect 237196 300092 237248 300144
rect 294144 300092 294196 300144
rect 369032 300092 369084 300144
rect 98920 300024 98972 300076
rect 233424 300024 233476 300076
rect 350632 300024 350684 300076
rect 371884 300024 371936 300076
rect 217968 299956 218020 300008
rect 292672 299956 292724 300008
rect 350724 299956 350776 300008
rect 371700 299956 371752 300008
rect 213552 299888 213604 299940
rect 286048 299888 286100 299940
rect 350816 299888 350868 299940
rect 371516 299888 371568 299940
rect 271144 299752 271196 299804
rect 271604 299752 271656 299804
rect 97908 299412 97960 299464
rect 241704 299412 241756 299464
rect 352656 299412 352708 299464
rect 580172 299412 580224 299464
rect 98644 299344 98696 299396
rect 239312 299344 239364 299396
rect 98828 299276 98880 299328
rect 237472 299276 237524 299328
rect 98552 299208 98604 299260
rect 236184 299208 236236 299260
rect 104532 299140 104584 299192
rect 234712 299140 234764 299192
rect 114836 299072 114888 299124
rect 242992 299072 243044 299124
rect 119988 299004 120040 299056
rect 246120 299004 246172 299056
rect 125140 298936 125192 298988
rect 239128 298936 239180 298988
rect 140596 298868 140648 298920
rect 249892 298868 249944 298920
rect 156052 298800 156104 298852
rect 250076 298800 250128 298852
rect 146944 298732 146996 298784
rect 248696 298732 248748 298784
rect 333244 298732 333296 298784
rect 538864 298732 538916 298784
rect 145748 298664 145800 298716
rect 236276 298664 236328 298716
rect 161204 298596 161256 298648
rect 247316 298596 247368 298648
rect 163780 298528 163832 298580
rect 234528 298528 234580 298580
rect 158628 298052 158680 298104
rect 169944 298052 169996 298104
rect 132868 297916 132920 297968
rect 247224 297916 247276 297968
rect 122564 297848 122616 297900
rect 236368 297848 236420 297900
rect 138020 297780 138072 297832
rect 237564 297780 237616 297832
rect 130292 297712 130344 297764
rect 146944 297712 146996 297764
rect 148324 297712 148376 297764
rect 234804 297712 234856 297764
rect 100024 297644 100076 297696
rect 172244 297644 172296 297696
rect 213736 297644 213788 297696
rect 291752 297644 291804 297696
rect 107108 297576 107160 297628
rect 170496 297576 170548 297628
rect 211712 297576 211764 297628
rect 290372 297576 290424 297628
rect 109684 297508 109736 297560
rect 170036 297508 170088 297560
rect 213276 297508 213328 297560
rect 338396 297508 338448 297560
rect 112260 297440 112312 297492
rect 172612 297440 172664 297492
rect 213184 297440 213236 297492
rect 339592 297440 339644 297492
rect 135444 297372 135496 297424
rect 171692 297372 171744 297424
rect 212264 297372 212316 297424
rect 291936 297372 291988 297424
rect 337292 297372 337344 297424
rect 567844 297372 567896 297424
rect 143172 297304 143224 297356
rect 172336 297304 172388 297356
rect 213644 297304 213696 297356
rect 290004 297304 290056 297356
rect 215944 297236 215996 297288
rect 291476 297236 291528 297288
rect 218796 297168 218848 297220
rect 290188 297168 290240 297220
rect 98736 297100 98788 297152
rect 245844 297100 245896 297152
rect 101956 297032 102008 297084
rect 247500 297032 247552 297084
rect 99104 296624 99156 296676
rect 240324 296624 240376 296676
rect 117320 296556 117372 296608
rect 243176 296556 243228 296608
rect 126980 296488 127032 296540
rect 247132 296488 247184 296540
rect 153200 296420 153252 296472
rect 247408 296420 247460 296472
rect 149060 296080 149112 296132
rect 273352 296080 273404 296132
rect 143540 296012 143592 296064
rect 272616 296012 272668 296064
rect 125600 295944 125652 295996
rect 269672 295944 269724 295996
rect 210884 295196 210936 295248
rect 283288 295196 283340 295248
rect 217876 295128 217928 295180
rect 293040 295128 293092 295180
rect 215852 295060 215904 295112
rect 292948 295060 293000 295112
rect 214380 294992 214432 295044
rect 292580 294992 292632 295044
rect 213092 294924 213144 294976
rect 291660 294924 291712 294976
rect 214472 294856 214524 294908
rect 292764 294856 292816 294908
rect 211620 294788 211672 294840
rect 291568 294788 291620 294840
rect 213000 294720 213052 294772
rect 292856 294720 292908 294772
rect 164240 294652 164292 294704
rect 275468 294652 275520 294704
rect 139400 294584 139452 294636
rect 271144 294584 271196 294636
rect 321928 294584 321980 294636
rect 471244 294584 471296 294636
rect 217692 293360 217744 293412
rect 341524 293360 341576 293412
rect 150440 293292 150492 293344
rect 273260 293292 273312 293344
rect 333152 293292 333204 293344
rect 543740 293292 543792 293344
rect 64880 293224 64932 293276
rect 260840 293224 260892 293276
rect 337200 293224 337252 293276
rect 571984 293224 572036 293276
rect 184204 291864 184256 291916
rect 276388 291864 276440 291916
rect 315212 291864 315264 291916
rect 422944 291864 422996 291916
rect 128360 291796 128412 291848
rect 269764 291796 269816 291848
rect 333060 291796 333112 291848
rect 547880 291796 547932 291848
rect 132500 290504 132552 290556
rect 271236 290504 271288 290556
rect 22744 290436 22796 290488
rect 254400 290436 254452 290488
rect 316500 290436 316552 290488
rect 431960 290436 432012 290488
rect 312452 289416 312504 289468
rect 407120 289416 407172 289468
rect 315120 289348 315172 289400
rect 413284 289348 413336 289400
rect 312544 289280 312596 289332
rect 411260 289280 411312 289332
rect 313924 289212 313976 289264
rect 415400 289212 415452 289264
rect 313832 289144 313884 289196
rect 418160 289144 418212 289196
rect 135260 289076 135312 289128
rect 270960 289076 271012 289128
rect 337108 289076 337160 289128
rect 575480 289076 575532 289128
rect 308312 287988 308364 288040
rect 382280 287988 382332 288040
rect 309784 287920 309836 287972
rect 386420 287920 386472 287972
rect 312636 287852 312688 287904
rect 400220 287852 400272 287904
rect 146300 287784 146352 287836
rect 272340 287784 272392 287836
rect 311072 287784 311124 287836
rect 404360 287784 404412 287836
rect 71044 287716 71096 287768
rect 261392 287716 261444 287768
rect 323676 287716 323728 287768
rect 471980 287716 472032 287768
rect 39304 287648 39356 287700
rect 257252 287648 257304 287700
rect 324872 287648 324924 287700
rect 488540 287648 488592 287700
rect 306932 286628 306984 286680
rect 375380 286628 375432 286680
rect 310980 286560 311032 286612
rect 397460 286560 397512 286612
rect 313740 286492 313792 286544
rect 416780 286492 416832 286544
rect 217784 286424 217836 286476
rect 338212 286424 338264 286476
rect 153200 286356 153252 286408
rect 273720 286356 273772 286408
rect 324780 286356 324832 286408
rect 492680 286356 492732 286408
rect 12440 286288 12492 286340
rect 253020 286288 253072 286340
rect 327632 286288 327684 286340
rect 509240 286288 509292 286340
rect 308496 285200 308548 285252
rect 372620 285200 372672 285252
rect 309692 285132 309744 285184
rect 391940 285132 391992 285184
rect 157340 285064 157392 285116
rect 275100 285064 275152 285116
rect 310888 285064 310940 285116
rect 396080 285064 396132 285116
rect 135352 284996 135404 285048
rect 270868 284996 270920 285048
rect 310796 284996 310848 285048
rect 398840 284996 398892 285048
rect 103520 284928 103572 284980
rect 266912 284928 266964 284980
rect 312360 284928 312412 284980
rect 414020 284928 414072 284980
rect 218428 283772 218480 283824
rect 283012 283772 283064 283824
rect 126980 283704 127032 283756
rect 269488 283704 269540 283756
rect 308220 283704 308272 283756
rect 378140 283704 378192 283756
rect 111800 283636 111852 283688
rect 268292 283636 268344 283688
rect 308128 283636 308180 283688
rect 385040 283636 385092 283688
rect 31760 283568 31812 283620
rect 249064 283568 249116 283620
rect 309600 283568 309652 283620
rect 389180 283568 389232 283620
rect 306748 282548 306800 282600
rect 371240 282548 371292 282600
rect 306840 282480 306892 282532
rect 374000 282480 374052 282532
rect 310704 282412 310756 282464
rect 402980 282412 403032 282464
rect 217416 282344 217468 282396
rect 342352 282344 342404 282396
rect 161480 282276 161532 282328
rect 275008 282276 275060 282328
rect 321836 282276 321888 282328
rect 475384 282276 475436 282328
rect 131120 282208 131172 282260
rect 270776 282208 270828 282260
rect 330392 282208 330444 282260
rect 524420 282208 524472 282260
rect 44180 282140 44232 282192
rect 257160 282140 257212 282192
rect 337016 282140 337068 282192
rect 574100 282140 574152 282192
rect 165620 280984 165672 281036
rect 274916 280984 274968 281036
rect 315028 280984 315080 281036
rect 426440 280984 426492 281036
rect 218704 280916 218756 280968
rect 339960 280916 340012 280968
rect 140780 280848 140832 280900
rect 272248 280848 272300 280900
rect 316408 280848 316460 280900
rect 440240 280848 440292 280900
rect 110420 280780 110472 280832
rect 268200 280780 268252 280832
rect 323492 280780 323544 280832
rect 481640 280780 481692 280832
rect 181444 279692 181496 279744
rect 277860 279692 277912 279744
rect 303988 279692 304040 279744
rect 357440 279692 357492 279744
rect 168472 279624 168524 279676
rect 276296 279624 276348 279676
rect 314936 279624 314988 279676
rect 430580 279624 430632 279676
rect 102140 279556 102192 279608
rect 266820 279556 266872 279608
rect 324688 279556 324740 279608
rect 491300 279556 491352 279608
rect 45560 279488 45612 279540
rect 246396 279488 246448 279540
rect 332968 279488 333020 279540
rect 547972 279488 548024 279540
rect 13084 279420 13136 279472
rect 252928 279420 252980 279472
rect 334532 279420 334584 279472
rect 556160 279420 556212 279472
rect 308036 278196 308088 278248
rect 382372 278196 382424 278248
rect 316316 278128 316368 278180
rect 440332 278128 440384 278180
rect 147680 278060 147732 278112
rect 273628 278060 273680 278112
rect 333336 278060 333388 278112
rect 534080 278060 534132 278112
rect 117320 277992 117372 278044
rect 251916 277992 251968 278044
rect 331772 277992 331824 278044
rect 540980 277992 541032 278044
rect 318156 276972 318208 277024
rect 433340 276972 433392 277024
rect 326160 276904 326212 276956
rect 506572 276904 506624 276956
rect 151820 276836 151872 276888
rect 273536 276836 273588 276888
rect 327540 276836 327592 276888
rect 511264 276836 511316 276888
rect 106280 276768 106332 276820
rect 266728 276768 266780 276820
rect 330300 276768 330352 276820
rect 531320 276768 531372 276820
rect 84200 276700 84252 276752
rect 264152 276700 264204 276752
rect 331680 276700 331732 276752
rect 542360 276700 542412 276752
rect 71780 276632 71832 276684
rect 261300 276632 261352 276684
rect 332876 276632 332928 276684
rect 546500 276632 546552 276684
rect 309508 275612 309560 275664
rect 393320 275612 393372 275664
rect 313648 275544 313700 275596
rect 419540 275544 419592 275596
rect 313556 275476 313608 275528
rect 423772 275476 423824 275528
rect 316224 275408 316276 275460
rect 434720 275408 434772 275460
rect 184940 275340 184992 275392
rect 278136 275340 278188 275392
rect 326068 275340 326120 275392
rect 498200 275340 498252 275392
rect 129740 275272 129792 275324
rect 270684 275272 270736 275324
rect 330208 275272 330260 275324
rect 527180 275272 527232 275324
rect 313464 274252 313516 274304
rect 415492 274252 415544 274304
rect 320824 274184 320876 274236
rect 469220 274184 469272 274236
rect 321744 274116 321796 274168
rect 473452 274116 473504 274168
rect 127072 274048 127124 274100
rect 269396 274048 269448 274100
rect 323400 274048 323452 274100
rect 476764 274048 476816 274100
rect 85580 273980 85632 274032
rect 264060 273980 264112 274032
rect 329012 273980 329064 274032
rect 516140 273980 516192 274032
rect 39396 273912 39448 273964
rect 255780 273912 255832 273964
rect 331588 273912 331640 273964
rect 538220 273912 538272 273964
rect 355324 273164 355376 273216
rect 579988 273164 580040 273216
rect 167000 272688 167052 272740
rect 276204 272688 276256 272740
rect 312268 272688 312320 272740
rect 407212 272688 407264 272740
rect 88340 272620 88392 272672
rect 263968 272620 264020 272672
rect 312176 272620 312228 272672
rect 412640 272620 412692 272672
rect 66260 272552 66312 272604
rect 261208 272552 261260 272604
rect 319536 272552 319588 272604
rect 449900 272552 449952 272604
rect 2780 272484 2832 272536
rect 251456 272484 251508 272536
rect 336004 272484 336056 272536
rect 569960 272484 570012 272536
rect 209780 271396 209832 271448
rect 282092 271396 282144 271448
rect 312084 271396 312136 271448
rect 408500 271396 408552 271448
rect 205640 271328 205692 271380
rect 282184 271328 282236 271380
rect 320732 271328 320784 271380
rect 465080 271328 465132 271380
rect 151912 271260 151964 271312
rect 273444 271260 273496 271312
rect 323308 271260 323360 271312
rect 484400 271260 484452 271312
rect 143632 271192 143684 271244
rect 272156 271192 272208 271244
rect 330116 271192 330168 271244
rect 528560 271192 528612 271244
rect 81440 271124 81492 271176
rect 257344 271124 257396 271176
rect 332784 271124 332836 271176
rect 552020 271124 552072 271176
rect 198740 270172 198792 270224
rect 278044 270172 278096 270224
rect 194600 270104 194652 270156
rect 275284 270104 275336 270156
rect 310612 270104 310664 270156
rect 401600 270104 401652 270156
rect 133880 270036 133932 270088
rect 270592 270036 270644 270088
rect 319444 270036 319496 270088
rect 458180 270036 458232 270088
rect 124220 269968 124272 270020
rect 269304 269968 269356 270020
rect 320640 269968 320692 270020
rect 465172 269968 465224 270020
rect 107660 269900 107712 269952
rect 266636 269900 266688 269952
rect 324596 269900 324648 269952
rect 495440 269900 495492 269952
rect 99380 269832 99432 269884
rect 265624 269832 265676 269884
rect 327448 269832 327500 269884
rect 504364 269832 504416 269884
rect 17960 269764 18012 269816
rect 252836 269764 252888 269816
rect 334440 269764 334492 269816
rect 558920 269764 558972 269816
rect 201500 268676 201552 268728
rect 280528 268676 280580 268728
rect 310520 268676 310572 268728
rect 398932 268676 398984 268728
rect 191840 268608 191892 268660
rect 279332 268608 279384 268660
rect 317972 268608 318024 268660
rect 447140 268608 447192 268660
rect 136640 268540 136692 268592
rect 271052 268540 271104 268592
rect 319352 268540 319404 268592
rect 455420 268540 455472 268592
rect 115940 268472 115992 268524
rect 268108 268472 268160 268524
rect 325884 268472 325936 268524
rect 502340 268472 502392 268524
rect 95240 268404 95292 268456
rect 265532 268404 265584 268456
rect 325976 268404 326028 268456
rect 503720 268404 503772 268456
rect 92480 268336 92532 268388
rect 265440 268336 265492 268388
rect 335912 268336 335964 268388
rect 565820 268336 565872 268388
rect 3516 267656 3568 267708
rect 225604 267656 225656 267708
rect 309324 267248 309376 267300
rect 390560 267248 390612 267300
rect 187700 267180 187752 267232
rect 279240 267180 279292 267232
rect 309416 267180 309468 267232
rect 394700 267180 394752 267232
rect 122840 267112 122892 267164
rect 269212 267112 269264 267164
rect 314844 267112 314896 267164
rect 427820 267112 427872 267164
rect 114560 267044 114612 267096
rect 268016 267044 268068 267096
rect 319260 267044 319312 267096
rect 451280 267044 451332 267096
rect 63500 266976 63552 267028
rect 260104 266976 260156 267028
rect 327356 266976 327408 267028
rect 514024 266976 514076 267028
rect 162860 265888 162912 265940
rect 274824 265888 274876 265940
rect 307944 265888 307996 265940
rect 383660 265888 383712 265940
rect 138020 265820 138072 265872
rect 272064 265820 272116 265872
rect 309232 265820 309284 265872
rect 387800 265820 387852 265872
rect 70400 265752 70452 265804
rect 261116 265752 261168 265804
rect 311992 265752 312044 265804
rect 405740 265752 405792 265804
rect 60740 265684 60792 265736
rect 260012 265684 260064 265736
rect 316132 265684 316184 265736
rect 438860 265684 438912 265736
rect 40040 265616 40092 265668
rect 257068 265616 257120 265668
rect 330024 265616 330076 265668
rect 531412 265616 531464 265668
rect 208400 264596 208452 264648
rect 281816 264596 281868 264648
rect 204260 264528 204312 264580
rect 281908 264528 281960 264580
rect 306564 264528 306616 264580
rect 376760 264528 376812 264580
rect 174544 264460 174596 264512
rect 276572 264460 276624 264512
rect 307852 264460 307904 264512
rect 380900 264460 380952 264512
rect 144920 264392 144972 264444
rect 271972 264392 272024 264444
rect 317880 264392 317932 264444
rect 448520 264392 448572 264444
rect 100760 264324 100812 264376
rect 265348 264324 265400 264376
rect 325792 264324 325844 264376
rect 499580 264324 499632 264376
rect 74540 264256 74592 264308
rect 262772 264256 262824 264308
rect 328920 264256 328972 264308
rect 521660 264256 521712 264308
rect 46204 264188 46256 264240
rect 256976 264188 257028 264240
rect 331496 264188 331548 264240
rect 539600 264188 539652 264240
rect 201592 263168 201644 263220
rect 280436 263168 280488 263220
rect 154580 263100 154632 263152
rect 273904 263100 273956 263152
rect 306380 263100 306432 263152
rect 374092 263100 374144 263152
rect 113180 263032 113232 263084
rect 267924 263032 267976 263084
rect 317696 263032 317748 263084
rect 441620 263032 441672 263084
rect 104900 262964 104952 263016
rect 266544 262964 266596 263016
rect 317788 262964 317840 263016
rect 444380 262964 444432 263016
rect 52460 262896 52512 262948
rect 251824 262896 251876 262948
rect 320548 262896 320600 262948
rect 466460 262896 466512 262948
rect 16580 262828 16632 262880
rect 252744 262828 252796 262880
rect 336924 262828 336976 262880
rect 578240 262828 578292 262880
rect 197360 261876 197412 261928
rect 280252 261876 280304 261928
rect 193220 261808 193272 261860
rect 280344 261808 280396 261860
rect 180800 261740 180852 261792
rect 277768 261740 277820 261792
rect 98000 261672 98052 261724
rect 265256 261672 265308 261724
rect 320456 261672 320508 261724
rect 462320 261672 462372 261724
rect 85672 261604 85724 261656
rect 263876 261604 263928 261656
rect 320364 261604 320416 261656
rect 463700 261604 463752 261656
rect 49700 261536 49752 261588
rect 258540 261536 258592 261588
rect 321652 261536 321704 261588
rect 474740 261536 474792 261588
rect 25596 261468 25648 261520
rect 252652 261468 252704 261520
rect 324504 261468 324556 261520
rect 496084 261468 496136 261520
rect 190460 260516 190512 260568
rect 279148 260516 279200 260568
rect 186320 260448 186372 260500
rect 279056 260448 279108 260500
rect 217600 260380 217652 260432
rect 338120 260380 338172 260432
rect 110512 260312 110564 260364
rect 250628 260312 250680 260364
rect 329932 260312 329984 260364
rect 532700 260312 532752 260364
rect 27620 260244 27672 260296
rect 254308 260244 254360 260296
rect 331312 260244 331364 260296
rect 536840 260244 536892 260296
rect 9680 260176 9732 260228
rect 253204 260176 253256 260228
rect 331404 260176 331456 260228
rect 539692 260176 539744 260228
rect 7564 260108 7616 260160
rect 251364 260108 251416 260160
rect 335820 260108 335872 260160
rect 568580 260108 568632 260160
rect 353944 259360 353996 259412
rect 579804 259360 579856 259412
rect 183560 258884 183612 258936
rect 272524 258884 272576 258936
rect 179420 258816 179472 258868
rect 277676 258816 277728 258868
rect 176660 258748 176712 258800
rect 277584 258748 277636 258800
rect 331956 258748 332008 258800
rect 525800 258748 525852 258800
rect 93860 258680 93912 258732
rect 265164 258680 265216 258732
rect 329840 258680 329892 258732
rect 529940 258680 529992 258732
rect 209872 257660 209924 257712
rect 281724 257660 281776 257712
rect 96620 257592 96672 257644
rect 265072 257592 265124 257644
rect 42800 257524 42852 257576
rect 256792 257524 256844 257576
rect 38660 257456 38712 257508
rect 256884 257456 256936 257508
rect 329196 257456 329248 257508
rect 514852 257456 514904 257508
rect 35900 257388 35952 257440
rect 255688 257388 255740 257440
rect 328828 257388 328880 257440
rect 523040 257388 523092 257440
rect 22100 257320 22152 257372
rect 254216 257320 254268 257372
rect 335728 257320 335780 257372
rect 564440 257320 564492 257372
rect 207020 256368 207072 256420
rect 281632 256368 281684 256420
rect 313372 256368 313424 256420
rect 422300 256368 422352 256420
rect 217140 256300 217192 256352
rect 342904 256300 342956 256352
rect 80060 256232 80112 256284
rect 262680 256232 262732 256284
rect 314752 256232 314804 256284
rect 428464 256232 428516 256284
rect 41420 256164 41472 256216
rect 256700 256164 256752 256216
rect 316040 256164 316092 256216
rect 436100 256164 436152 256216
rect 34520 256096 34572 256148
rect 255412 256096 255464 256148
rect 317604 256096 317656 256148
rect 443000 256096 443052 256148
rect 30380 256028 30432 256080
rect 255596 256028 255648 256080
rect 325700 256028 325752 256080
rect 505100 256028 505152 256080
rect 27712 255960 27764 256012
rect 255504 255960 255556 256012
rect 327264 255960 327316 256012
rect 512000 255960 512052 256012
rect 3516 255144 3568 255196
rect 8944 255144 8996 255196
rect 202880 254940 202932 254992
rect 281540 254940 281592 254992
rect 200120 254872 200172 254924
rect 280620 254872 280672 254924
rect 307760 254872 307812 254924
rect 379520 254872 379572 254924
rect 102232 254804 102284 254856
rect 266452 254804 266504 254856
rect 309140 254804 309192 254856
rect 390652 254804 390704 254856
rect 93952 254736 94004 254788
rect 264980 254736 265032 254788
rect 320272 254736 320324 254788
rect 460940 254736 460992 254788
rect 91100 254668 91152 254720
rect 263784 254668 263836 254720
rect 329104 254668 329156 254720
rect 498292 254668 498344 254720
rect 77300 254600 77352 254652
rect 262588 254600 262640 254652
rect 334348 254600 334400 254652
rect 556252 254600 556304 254652
rect 73160 254532 73212 254584
rect 261024 254532 261076 254584
rect 334256 254532 334308 254584
rect 560300 254532 560352 254584
rect 193312 253648 193364 253700
rect 278964 253648 279016 253700
rect 217048 253580 217100 253632
rect 340972 253580 341024 253632
rect 121460 253512 121512 253564
rect 269580 253512 269632 253564
rect 319168 253512 319220 253564
rect 456800 253512 456852 253564
rect 118700 253444 118752 253496
rect 267832 253444 267884 253496
rect 323216 253444 323268 253496
rect 485780 253444 485832 253496
rect 82820 253376 82872 253428
rect 262496 253376 262548 253428
rect 324412 253376 324464 253428
rect 489920 253376 489972 253428
rect 69020 253308 69072 253360
rect 260932 253308 260984 253360
rect 327172 253308 327224 253360
rect 507860 253308 507912 253360
rect 62120 253240 62172 253292
rect 259920 253240 259972 253292
rect 331220 253240 331272 253292
rect 535460 253240 535512 253292
rect 23480 253172 23532 253224
rect 250536 253172 250588 253224
rect 335636 253172 335688 253224
rect 561680 253172 561732 253224
rect 218520 252152 218572 252204
rect 341432 252152 341484 252204
rect 86960 252084 87012 252136
rect 263692 252084 263744 252136
rect 313280 252084 313332 252136
rect 420920 252084 420972 252136
rect 78680 252016 78732 252068
rect 262404 252016 262456 252068
rect 319076 252016 319128 252068
rect 459560 252016 459612 252068
rect 26240 251948 26292 252000
rect 254032 251948 254084 252000
rect 328736 251948 328788 252000
rect 518900 251948 518952 252000
rect 19340 251880 19392 251932
rect 254124 251880 254176 251932
rect 332692 251880 332744 251932
rect 549260 251880 549312 251932
rect 8300 251812 8352 251864
rect 251272 251812 251324 251864
rect 335544 251812 335596 251864
rect 564532 251812 564584 251864
rect 301504 251132 301556 251184
rect 363052 251132 363104 251184
rect 301320 251064 301372 251116
rect 362960 251064 363012 251116
rect 301412 250996 301464 251048
rect 363236 250996 363288 251048
rect 298284 250928 298336 250980
rect 360660 250928 360712 250980
rect 300032 250860 300084 250912
rect 363144 250860 363196 250912
rect 311900 250792 311952 250844
rect 409880 250792 409932 250844
rect 142160 250724 142212 250776
rect 272432 250724 272484 250776
rect 317512 250724 317564 250776
rect 445760 250724 445812 250776
rect 77392 250656 77444 250708
rect 262312 250656 262364 250708
rect 325056 250656 325108 250708
rect 487160 250656 487212 250708
rect 75920 250588 75972 250640
rect 262864 250588 262916 250640
rect 327816 250588 327868 250640
rect 494060 250588 494112 250640
rect 55220 250520 55272 250572
rect 259828 250520 259880 250572
rect 328644 250520 328696 250572
rect 517520 250520 517572 250572
rect 11060 250452 11112 250504
rect 246304 250452 246356 250504
rect 336832 250452 336884 250504
rect 576860 250452 576912 250504
rect 189080 249364 189132 249416
rect 278872 249364 278924 249416
rect 89720 249296 89772 249348
rect 263600 249296 263652 249348
rect 318892 249296 318944 249348
rect 452660 249296 452712 249348
rect 60832 249228 60884 249280
rect 259644 249228 259696 249280
rect 318984 249228 319036 249280
rect 456892 249228 456944 249280
rect 56600 249160 56652 249212
rect 259736 249160 259788 249212
rect 324320 249160 324372 249212
rect 490012 249160 490064 249212
rect 48320 249092 48372 249144
rect 258448 249092 258500 249144
rect 328552 249092 328604 249144
rect 523132 249092 523184 249144
rect 4160 249024 4212 249076
rect 243544 249024 243596 249076
rect 335452 249024 335504 249076
rect 567200 249024 567252 249076
rect 303804 248344 303856 248396
rect 361948 248344 362000 248396
rect 302608 248276 302660 248328
rect 361764 248276 361816 248328
rect 301228 248208 301280 248260
rect 360568 248208 360620 248260
rect 204904 248140 204956 248192
rect 258356 248140 258408 248192
rect 301044 248140 301096 248192
rect 360476 248140 360528 248192
rect 185032 248072 185084 248124
rect 279424 248072 279476 248124
rect 301136 248072 301188 248124
rect 361672 248072 361724 248124
rect 182180 248004 182232 248056
rect 277492 248004 277544 248056
rect 299848 248004 299900 248056
rect 360752 248004 360804 248056
rect 173900 247936 173952 247988
rect 276020 247936 276072 247988
rect 299940 247936 299992 247988
rect 361856 247936 361908 247988
rect 155960 247868 156012 247920
rect 273812 247868 273864 247920
rect 297088 247868 297140 247920
rect 365812 247868 365864 247920
rect 67640 247800 67692 247852
rect 261484 247800 261536 247852
rect 317420 247800 317472 247852
rect 448612 247800 448664 247852
rect 57980 247732 58032 247784
rect 259552 247732 259604 247784
rect 318800 247732 318852 247784
rect 454040 247732 454092 247784
rect 20720 247664 20772 247716
rect 254492 247664 254544 247716
rect 321560 247664 321612 247716
rect 477500 247664 477552 247716
rect 299756 247596 299808 247648
rect 357716 247596 357768 247648
rect 302516 247528 302568 247580
rect 360384 247528 360436 247580
rect 347136 247460 347188 247512
rect 369860 247460 369912 247512
rect 178040 246644 178092 246696
rect 277952 246644 278004 246696
rect 118792 246576 118844 246628
rect 268384 246576 268436 246628
rect 327080 246576 327132 246628
rect 510620 246576 510672 246628
rect 59360 246508 59412 246560
rect 259460 246508 259512 246560
rect 333980 246508 334032 246560
rect 553400 246508 553452 246560
rect 53840 246440 53892 246492
rect 258264 246440 258316 246492
rect 334072 246440 334124 246492
rect 554780 246440 554832 246492
rect 51080 246372 51132 246424
rect 258172 246372 258224 246424
rect 335360 246372 335412 246424
rect 563060 246372 563112 246424
rect 6920 246304 6972 246356
rect 251548 246304 251600 246356
rect 352564 246304 352616 246356
rect 580172 246304 580224 246356
rect 300952 245556 301004 245608
rect 359280 245556 359332 245608
rect 362500 245556 362552 245608
rect 365720 245556 365772 245608
rect 299664 245488 299716 245540
rect 359004 245488 359056 245540
rect 299480 245420 299532 245472
rect 358912 245420 358964 245472
rect 299572 245352 299624 245404
rect 359188 245352 359240 245404
rect 160192 245284 160244 245336
rect 275192 245284 275244 245336
rect 296904 245284 296956 245336
rect 357808 245284 357860 245336
rect 158720 245216 158772 245268
rect 274732 245216 274784 245268
rect 296812 245216 296864 245268
rect 359372 245216 359424 245268
rect 217232 245148 217284 245200
rect 336740 245148 336792 245200
rect 349896 245148 349948 245200
rect 362040 245148 362092 245200
rect 120080 245080 120132 245132
rect 250444 245080 250496 245132
rect 295800 245080 295852 245132
rect 363328 245080 363380 245132
rect 109040 245012 109092 245064
rect 267004 245012 267056 245064
rect 298100 245012 298152 245064
rect 368480 245012 368532 245064
rect 46940 244944 46992 244996
rect 258632 244944 258684 244996
rect 296720 244944 296772 244996
rect 367192 244944 367244 244996
rect 35992 244876 36044 244928
rect 255964 244876 256016 244928
rect 314660 244876 314712 244928
rect 432052 244876 432104 244928
rect 300860 244808 300912 244860
rect 359096 244808 359148 244860
rect 302332 244740 302384 244792
rect 357624 244740 357676 244792
rect 355416 244468 355468 244520
rect 363420 244468 363472 244520
rect 218612 243720 218664 243772
rect 293224 243720 293276 243772
rect 295708 243720 295760 243772
rect 357900 243720 357952 243772
rect 219256 243652 219308 243704
rect 293960 243652 294012 243704
rect 295616 243652 295668 243704
rect 359464 243652 359516 243704
rect 217508 243584 217560 243636
rect 294052 243584 294104 243636
rect 295524 243584 295576 243636
rect 360844 243584 360896 243636
rect 215760 243516 215812 243568
rect 293132 243516 293184 243568
rect 295340 243516 295392 243568
rect 362132 243516 362184 243568
rect 3516 241408 3568 241460
rect 14556 241408 14608 241460
rect 577596 219172 577648 219224
rect 579712 219172 579764 219224
rect 3332 215228 3384 215280
rect 209044 215228 209096 215280
rect 358084 206932 358136 206984
rect 579620 206932 579672 206984
rect 358360 204824 358412 204876
rect 363788 204824 363840 204876
rect 358268 204688 358320 204740
rect 363788 204688 363840 204740
rect 3056 202784 3108 202836
rect 199384 202784 199436 202836
rect 214380 195508 214432 195560
rect 217140 195508 217192 195560
rect 213000 195236 213052 195288
rect 217324 195236 217376 195288
rect 210884 193128 210936 193180
rect 216772 193128 216824 193180
rect 215852 189388 215904 189440
rect 218520 189388 218572 189440
rect 3516 188980 3568 189032
rect 206284 188980 206336 189032
rect 210976 188980 211028 189032
rect 216680 188980 216732 189032
rect 577504 179324 577556 179376
rect 579712 179324 579764 179376
rect 212080 159876 212132 159928
rect 256700 159876 256752 159928
rect 218796 159808 218848 159860
rect 264980 159808 265032 159860
rect 216312 159740 216364 159792
rect 263600 159740 263652 159792
rect 213460 159672 213512 159724
rect 260840 159672 260892 159724
rect 213092 159604 213144 159656
rect 269120 159604 269172 159656
rect 217140 159536 217192 159588
rect 276204 159536 276256 159588
rect 313464 159536 313516 159588
rect 373264 159536 373316 159588
rect 215944 159468 215996 159520
rect 276020 159468 276072 159520
rect 298468 159468 298520 159520
rect 358176 159468 358228 159520
rect 217876 159400 217928 159452
rect 278780 159400 278832 159452
rect 310980 159400 311032 159452
rect 371608 159400 371660 159452
rect 214472 159332 214524 159384
rect 282920 159332 282972 159384
rect 303528 159332 303580 159384
rect 369216 159332 369268 159384
rect 295892 159264 295944 159316
rect 369124 159264 369176 159316
rect 293500 159196 293552 159248
rect 370688 159196 370740 159248
rect 276112 159128 276164 159180
rect 363696 159128 363748 159180
rect 278504 159060 278556 159112
rect 367928 159060 367980 159112
rect 273628 158992 273680 159044
rect 367836 158992 367888 159044
rect 213276 158924 213328 158976
rect 238208 158924 238260 158976
rect 265348 158924 265400 158976
rect 359648 158924 359700 158976
rect 213184 158856 213236 158908
rect 239588 158856 239640 158908
rect 263968 158856 264020 158908
rect 363604 158856 363656 158908
rect 213368 158788 213420 158840
rect 241704 158788 241756 158840
rect 262864 158788 262916 158840
rect 364616 158788 364668 158840
rect 211988 158720 212040 158772
rect 240508 158720 240560 158772
rect 259552 158720 259604 158772
rect 364708 158720 364760 158772
rect 219072 158652 219124 158704
rect 234620 158652 234672 158704
rect 248328 158652 248380 158704
rect 365168 158652 365220 158704
rect 216128 158584 216180 158636
rect 233240 158584 233292 158636
rect 256056 158584 256108 158636
rect 371792 158584 371844 158636
rect 214840 158516 214892 158568
rect 236000 158516 236052 158568
rect 261208 158516 261260 158568
rect 373172 158516 373224 158568
rect 211896 158448 211948 158500
rect 234712 158448 234764 158500
rect 255964 158448 256016 158500
rect 364432 158448 364484 158500
rect 218980 158380 219032 158432
rect 242992 158380 243044 158432
rect 257160 158380 257212 158432
rect 364340 158380 364392 158432
rect 214656 158312 214708 158364
rect 242900 158312 242952 158364
rect 254584 158312 254636 158364
rect 360936 158312 360988 158364
rect 214932 158244 214984 158296
rect 245660 158244 245712 158296
rect 258264 158244 258316 158296
rect 364524 158244 364576 158296
rect 216220 158176 216272 158228
rect 247040 158176 247092 158228
rect 265992 158176 266044 158228
rect 369308 158176 369360 158228
rect 216404 158108 216456 158160
rect 249800 158108 249852 158160
rect 291016 158108 291068 158160
rect 370596 158108 370648 158160
rect 218888 158040 218940 158092
rect 252560 158040 252612 158092
rect 300952 158040 301004 158092
rect 370504 158040 370556 158092
rect 211620 157972 211672 158024
rect 273260 157972 273312 158024
rect 308680 157972 308732 158024
rect 372988 157972 373040 158024
rect 216036 157904 216088 157956
rect 230480 157904 230532 157956
rect 321100 157904 321152 157956
rect 371700 157904 371752 157956
rect 214748 157836 214800 157888
rect 229100 157836 229152 157888
rect 323400 157836 323452 157888
rect 371884 157836 371936 157888
rect 219164 157768 219216 157820
rect 227720 157768 227772 157820
rect 325976 157768 326028 157820
rect 373080 157768 373132 157820
rect 250168 157292 250220 157344
rect 368572 157292 368624 157344
rect 251456 157224 251508 157276
rect 368848 157224 368900 157276
rect 267648 157156 267700 157208
rect 367376 157156 367428 157208
rect 268752 157088 268804 157140
rect 367652 157088 367704 157140
rect 271144 157020 271196 157072
rect 367744 157020 367796 157072
rect 266820 156952 266872 157004
rect 363512 156952 363564 157004
rect 269856 156884 269908 156936
rect 365904 156884 365956 156936
rect 272248 156816 272300 156868
rect 366272 156816 366324 156868
rect 274180 156748 274232 156800
rect 367560 156748 367612 156800
rect 274456 156680 274508 156732
rect 366364 156680 366416 156732
rect 275928 156612 275980 156664
rect 367284 156612 367336 156664
rect 277124 156544 277176 156596
rect 366088 156544 366140 156596
rect 279976 156476 280028 156528
rect 366180 156476 366232 156528
rect 278136 156408 278188 156460
rect 361120 156408 361172 156460
rect 252376 155864 252428 155916
rect 368664 155864 368716 155916
rect 251088 155796 251140 155848
rect 366456 155796 366508 155848
rect 213552 155728 213604 155780
rect 237380 155728 237432 155780
rect 253572 155728 253624 155780
rect 367468 155728 367520 155780
rect 211804 155660 211856 155712
rect 241520 155660 241572 155712
rect 268936 155660 268988 155712
rect 365076 155660 365128 155712
rect 214564 155592 214616 155644
rect 248420 155592 248472 155644
rect 281080 155592 281132 155644
rect 370228 155592 370280 155644
rect 211068 155524 211120 155576
rect 255320 155524 255372 155576
rect 283748 155524 283800 155576
rect 370044 155524 370096 155576
rect 211712 155456 211764 155508
rect 259552 155456 259604 155508
rect 286508 155456 286560 155508
rect 370136 155456 370188 155508
rect 218612 155388 218664 155440
rect 280160 155388 280212 155440
rect 348516 155388 348568 155440
rect 369032 155388 369084 155440
rect 218520 155320 218572 155372
rect 284392 155320 284444 155372
rect 292580 155320 292632 155372
rect 357992 155320 358044 155372
rect 217508 155252 217560 155304
rect 285680 155252 285732 155304
rect 292672 155252 292724 155304
rect 363788 155252 363840 155304
rect 215760 155184 215812 155236
rect 284300 155184 284352 155236
rect 289820 155184 289872 155236
rect 370412 155184 370464 155236
rect 348424 155116 348476 155168
rect 366548 155116 366600 155168
rect 253664 154504 253716 154556
rect 372896 154504 372948 154556
rect 258632 154436 258684 154488
rect 370320 154436 370372 154488
rect 263968 154368 264020 154420
rect 371424 154368 371476 154420
rect 271052 154300 271104 154352
rect 372804 154300 372856 154352
rect 288256 154232 288308 154284
rect 369952 154232 370004 154284
rect 306104 154164 306156 154216
rect 371332 154164 371384 154216
rect 315856 154096 315908 154148
rect 371516 154096 371568 154148
rect 318616 154028 318668 154080
rect 372712 154028 372764 154080
rect 3516 150356 3568 150408
rect 210424 150356 210476 150408
rect 3516 137912 3568 137964
rect 203524 137912 203576 137964
rect 3516 97928 3568 97980
rect 198004 97928 198056 97980
rect 3516 85484 3568 85536
rect 200764 85484 200816 85536
rect 3516 71680 3568 71732
rect 207664 71680 207716 71732
rect 3516 59304 3568 59356
rect 25504 59304 25556 59356
rect 3424 20612 3476 20664
rect 196624 20612 196676 20664
rect 160100 11704 160152 11756
rect 161296 11704 161348 11756
rect 201500 11704 201552 11756
rect 202696 11704 202748 11756
rect 234620 11704 234672 11756
rect 235816 11704 235868 11756
rect 242900 11704 242952 11756
rect 244096 11704 244148 11756
rect 316224 9324 316276 9376
rect 363420 9324 363472 9376
rect 312636 9256 312688 9308
rect 360292 9256 360344 9308
rect 298468 9188 298520 9240
rect 357900 9188 357952 9240
rect 301964 9120 302016 9172
rect 362132 9120 362184 9172
rect 300768 9052 300820 9104
rect 360844 9052 360896 9104
rect 304356 8984 304408 9036
rect 365812 8984 365864 9036
rect 297272 8916 297324 8968
rect 359464 8916 359516 8968
rect 3424 6808 3476 6860
rect 88984 6808 89036 6860
rect 317328 6808 317380 6860
rect 358820 6808 358872 6860
rect 322112 6740 322164 6792
rect 368480 6740 368532 6792
rect 320916 6672 320968 6724
rect 367100 6672 367152 6724
rect 315028 6604 315080 6656
rect 361580 6604 361632 6656
rect 313832 6536 313884 6588
rect 360660 6536 360712 6588
rect 318524 6468 318576 6520
rect 365720 6468 365772 6520
rect 310244 6400 310296 6452
rect 357808 6400 357860 6452
rect 311440 6332 311492 6384
rect 359372 6332 359424 6384
rect 307944 6264 307996 6316
rect 356796 6264 356848 6316
rect 306748 6196 306800 6248
rect 367192 6196 367244 6248
rect 303160 6128 303212 6180
rect 363328 6128 363380 6180
rect 326804 6060 326856 6112
rect 360752 6060 360804 6112
rect 323308 5992 323360 6044
rect 357716 5992 357768 6044
rect 330392 5924 330444 5976
rect 363144 5924 363196 5976
rect 44272 4088 44324 4140
rect 46204 4088 46256 4140
rect 213828 4088 213880 4140
rect 260656 4088 260708 4140
rect 332692 4088 332744 4140
rect 360476 4088 360528 4140
rect 467104 4088 467156 4140
rect 467656 4088 467708 4140
rect 219348 4020 219400 4072
rect 266544 4020 266596 4072
rect 328000 4020 328052 4072
rect 359188 4020 359240 4072
rect 177856 3952 177908 4004
rect 181444 3952 181496 4004
rect 216588 3952 216640 4004
rect 267740 3952 267792 4004
rect 324412 3952 324464 4004
rect 357532 3952 357584 4004
rect 215208 3884 215260 3936
rect 262956 3884 263008 3936
rect 329196 3884 329248 3936
rect 361856 3884 361908 3936
rect 4068 3816 4120 3868
rect 7564 3816 7616 3868
rect 213736 3816 213788 3868
rect 268844 3816 268896 3868
rect 325608 3816 325660 3868
rect 359004 3816 359056 3868
rect 69112 3748 69164 3800
rect 71044 3748 71096 3800
rect 135260 3748 135312 3800
rect 136456 3748 136508 3800
rect 170772 3748 170824 3800
rect 174544 3748 174596 3800
rect 212448 3748 212500 3800
rect 271236 3748 271288 3800
rect 309048 3748 309100 3800
rect 356704 3748 356756 3800
rect 357348 3748 357400 3800
rect 362040 3748 362092 3800
rect 25320 3680 25372 3732
rect 171876 3680 171928 3732
rect 217968 3680 218020 3732
rect 278320 3680 278372 3732
rect 294880 3680 294932 3732
rect 348516 3680 348568 3732
rect 349252 3680 349304 3732
rect 357624 3680 357676 3732
rect 1676 3544 1728 3596
rect 14464 3612 14516 3664
rect 14740 3612 14792 3664
rect 25596 3612 25648 3664
rect 33600 3612 33652 3664
rect 39396 3612 39448 3664
rect 52552 3612 52604 3664
rect 204904 3612 204956 3664
rect 212264 3612 212316 3664
rect 272432 3612 272484 3664
rect 291384 3612 291436 3664
rect 348424 3612 348476 3664
rect 350448 3612 350500 3664
rect 361948 3612 362000 3664
rect 12348 3544 12400 3596
rect 13084 3544 13136 3596
rect 15936 3544 15988 3596
rect 170404 3544 170456 3596
rect 193220 3544 193272 3596
rect 194416 3544 194468 3596
rect 215024 3544 215076 3596
rect 274824 3544 274876 3596
rect 292580 3544 292632 3596
rect 293316 3544 293368 3596
rect 296076 3544 296128 3596
rect 353944 3544 353996 3596
rect 357532 3544 357584 3596
rect 369308 3544 369360 3596
rect 413284 3544 413336 3596
rect 426164 3544 426216 3596
rect 475384 3544 475436 3596
rect 476948 3544 477000 3596
rect 496084 3544 496136 3596
rect 497096 3544 497148 3596
rect 498200 3544 498252 3596
rect 499028 3544 499080 3596
rect 504364 3544 504416 3596
rect 507676 3544 507728 3596
rect 511264 3544 511316 3596
rect 513564 3544 513616 3596
rect 514024 3544 514076 3596
rect 514760 3544 514812 3596
rect 538864 3544 538916 3596
rect 551468 3544 551520 3596
rect 564440 3544 564492 3596
rect 565268 3544 565320 3596
rect 6460 3476 6512 3528
rect 172060 3476 172112 3528
rect 217324 3476 217376 3528
rect 281908 3476 281960 3528
rect 299664 3476 299716 3528
rect 357348 3476 357400 3528
rect 357440 3476 357492 3528
rect 358728 3476 358780 3528
rect 374000 3476 374052 3528
rect 375288 3476 375340 3528
rect 390560 3476 390612 3528
rect 391848 3476 391900 3528
rect 415492 3476 415544 3528
rect 416688 3476 416740 3528
rect 422944 3476 422996 3528
rect 424968 3476 425020 3528
rect 428556 3476 428608 3528
rect 429660 3476 429712 3528
rect 431960 3476 432012 3528
rect 433248 3476 433300 3528
rect 440332 3476 440384 3528
rect 441528 3476 441580 3528
rect 448612 3476 448664 3528
rect 449808 3476 449860 3528
rect 465080 3476 465132 3528
rect 465908 3476 465960 3528
rect 471244 3476 471296 3528
rect 473452 3476 473504 3528
rect 480904 3476 480956 3528
rect 581000 3476 581052 3528
rect 572 3408 624 3460
rect 171784 3408 171836 3460
rect 173164 3408 173216 3460
rect 184204 3408 184256 3460
rect 219164 3408 219216 3460
rect 287796 3408 287848 3460
rect 288992 3408 289044 3460
rect 354128 3408 354180 3460
rect 356336 3408 356388 3460
rect 369860 3408 369912 3460
rect 378784 3408 378836 3460
rect 572720 3408 572772 3460
rect 38384 3340 38436 3392
rect 39304 3340 39356 3392
rect 93860 3340 93912 3392
rect 94780 3340 94832 3392
rect 110420 3340 110472 3392
rect 111616 3340 111668 3392
rect 213644 3340 213696 3392
rect 258264 3340 258316 3392
rect 331588 3340 331640 3392
rect 358912 3340 358964 3392
rect 171968 3272 172020 3324
rect 175924 3272 175976 3324
rect 212080 3272 212132 3324
rect 254676 3272 254728 3324
rect 336280 3272 336332 3324
rect 356152 3272 356204 3324
rect 212356 3204 212408 3256
rect 245200 3204 245252 3256
rect 335084 3204 335136 3256
rect 359280 3204 359332 3256
rect 567844 3204 567896 3256
rect 571524 3204 571576 3256
rect 354036 3136 354088 3188
rect 360936 3136 360988 3188
rect 356152 3068 356204 3120
rect 361672 3068 361724 3120
rect 476764 3068 476816 3120
rect 479340 3068 479392 3120
rect 30104 3000 30156 3052
rect 32404 3000 32456 3052
rect 355232 3000 355284 3052
rect 362224 3000 362276 3052
rect 467656 3000 467708 3052
rect 471060 3000 471112 3052
rect 571984 3000 572036 3052
rect 573916 3000 573968 3052
rect 20628 2864 20680 2916
rect 22744 2864 22796 2916
rect 398840 2184 398892 2236
rect 400128 2184 400180 2236
rect 407120 2184 407172 2236
rect 408408 2184 408460 2236
rect 456800 2184 456852 2236
rect 458088 2184 458140 2236
rect 382280 1912 382332 1964
rect 383568 1912 383620 1964
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 700398 8156 703520
rect 8116 700392 8168 700398
rect 8116 700334 8168 700340
rect 13084 700392 13136 700398
rect 13084 700334 13136 700340
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 10324 683188 10376 683194
rect 10324 683130 10376 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 8944 632120 8996 632126
rect 3476 632088 3478 632097
rect 8944 632062 8996 632068
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3422 606112 3478 606121
rect 3422 606047 3424 606056
rect 3476 606047 3478 606056
rect 7564 606076 7616 606082
rect 3424 606018 3476 606024
rect 7564 606018 7616 606024
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 553450 3464 553823
rect 3424 553444 3476 553450
rect 3424 553386 3476 553392
rect 2778 527912 2834 527921
rect 2778 527847 2834 527856
rect 2792 527202 2820 527847
rect 2780 527196 2832 527202
rect 2780 527138 2832 527144
rect 4804 527196 4856 527202
rect 4804 527138 4856 527144
rect 3422 514856 3478 514865
rect 3422 514791 3478 514800
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 3436 480254 3464 514791
rect 3436 480226 3556 480254
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3436 474774 3464 475623
rect 3424 474768 3476 474774
rect 3424 474710 3476 474716
rect 3528 471306 3556 480226
rect 3516 471300 3568 471306
rect 3516 471242 3568 471248
rect 3238 462632 3294 462641
rect 3238 462567 3294 462576
rect 3252 462398 3280 462567
rect 3240 462392 3292 462398
rect 3240 462334 3292 462340
rect 4816 461718 4844 527138
rect 4804 461712 4856 461718
rect 4804 461654 4856 461660
rect 7576 451926 7604 606018
rect 8956 458930 8984 632062
rect 8944 458924 8996 458930
rect 8944 458866 8996 458872
rect 10336 456074 10364 683130
rect 10324 456068 10376 456074
rect 10324 456010 10376 456016
rect 7564 451920 7616 451926
rect 7564 451862 7616 451868
rect 13096 450566 13124 700334
rect 24320 699718 24348 703520
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 25504 699712 25556 699718
rect 25504 699654 25556 699660
rect 14464 656940 14516 656946
rect 14464 656882 14516 656888
rect 13084 450560 13136 450566
rect 13084 450502 13136 450508
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 14476 440978 14504 656882
rect 21364 565888 21416 565894
rect 21364 565830 21416 565836
rect 17224 553444 17276 553450
rect 17224 553386 17276 553392
rect 17236 474026 17264 553386
rect 18604 501016 18656 501022
rect 18604 500958 18656 500964
rect 18616 478174 18644 500958
rect 18604 478168 18656 478174
rect 18604 478110 18656 478116
rect 17224 474020 17276 474026
rect 17224 473962 17276 473968
rect 21376 467226 21404 565830
rect 25516 469878 25544 699654
rect 32404 579692 32456 579698
rect 32404 579634 32456 579640
rect 25504 469872 25556 469878
rect 25504 469814 25556 469820
rect 21364 467220 21416 467226
rect 21364 467162 21416 467168
rect 32416 460222 32444 579634
rect 32404 460216 32456 460222
rect 32404 460158 32456 460164
rect 40052 454714 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 40040 454708 40092 454714
rect 40040 454650 40092 454656
rect 71792 447914 71820 702986
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 88352 465798 88380 702406
rect 105464 700330 105492 703520
rect 137848 700398 137876 703520
rect 154132 702434 154160 703520
rect 170324 702434 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 153212 702406 154160 702434
rect 169772 702406 170352 702434
rect 137836 700392 137888 700398
rect 137836 700334 137888 700340
rect 138664 700392 138716 700398
rect 138664 700334 138716 700340
rect 105452 700324 105504 700330
rect 105452 700266 105504 700272
rect 88340 465792 88392 465798
rect 88340 465734 88392 465740
rect 71780 447908 71832 447914
rect 71780 447850 71832 447856
rect 138676 446418 138704 700334
rect 153212 457502 153240 702406
rect 153200 457496 153252 457502
rect 153200 457438 153252 457444
rect 169772 453422 169800 702406
rect 180064 670744 180116 670750
rect 180064 670686 180116 670692
rect 180076 464438 180104 670686
rect 182824 618316 182876 618322
rect 182824 618258 182876 618264
rect 180064 464432 180116 464438
rect 180064 464374 180116 464380
rect 169760 453416 169812 453422
rect 169760 453358 169812 453364
rect 138664 446412 138716 446418
rect 138664 446354 138716 446360
rect 182836 442338 182864 618258
rect 201512 443834 201540 702986
rect 217968 700392 218020 700398
rect 217968 700334 218020 700340
rect 206284 700324 206336 700330
rect 206284 700266 206336 700272
rect 206296 445194 206324 700266
rect 217876 565140 217928 565146
rect 217876 565082 217928 565088
rect 217782 516896 217838 516905
rect 217782 516831 217838 516840
rect 217690 515944 217746 515953
rect 217690 515879 217746 515888
rect 217598 513768 217654 513777
rect 217598 513703 217654 513712
rect 217414 489968 217470 489977
rect 217414 489903 217470 489912
rect 217322 488064 217378 488073
rect 217322 487999 217378 488008
rect 217336 450702 217364 487999
rect 217428 478446 217456 489903
rect 217506 488336 217562 488345
rect 217506 488271 217562 488280
rect 217416 478440 217468 478446
rect 217416 478382 217468 478388
rect 217520 471374 217548 488271
rect 217612 475386 217640 513703
rect 217600 475380 217652 475386
rect 217600 475322 217652 475328
rect 217508 471368 217560 471374
rect 217508 471310 217560 471316
rect 217704 468586 217732 515879
rect 217692 468580 217744 468586
rect 217692 468522 217744 468528
rect 217796 465866 217824 516831
rect 217784 465860 217836 465866
rect 217784 465802 217836 465808
rect 217324 450696 217376 450702
rect 217324 450638 217376 450644
rect 206284 445188 206336 445194
rect 206284 445130 206336 445136
rect 201500 443828 201552 443834
rect 201500 443770 201552 443776
rect 182824 442332 182876 442338
rect 182824 442274 182876 442280
rect 14464 440972 14516 440978
rect 14464 440914 14516 440920
rect 210424 436620 210476 436626
rect 210424 436562 210476 436568
rect 203524 436552 203576 436558
rect 203524 436494 203576 436500
rect 198004 436484 198056 436490
rect 198004 436426 198056 436432
rect 88984 436280 89036 436286
rect 88984 436222 89036 436228
rect 14556 436212 14608 436218
rect 14556 436154 14608 436160
rect 8944 436144 8996 436150
rect 8944 436086 8996 436092
rect 7564 434920 7616 434926
rect 7564 434862 7616 434868
rect 3608 432744 3660 432750
rect 3608 432686 3660 432692
rect 3516 432676 3568 432682
rect 3516 432618 3568 432624
rect 3424 432608 3476 432614
rect 3424 432550 3476 432556
rect 3332 423632 3384 423638
rect 3330 423600 3332 423609
rect 3384 423600 3386 423609
rect 3330 423535 3386 423544
rect 3332 411256 3384 411262
rect 3332 411198 3384 411204
rect 3344 410553 3372 411198
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 3332 398812 3384 398818
rect 3332 398754 3384 398760
rect 3344 397497 3372 398754
rect 3330 397488 3386 397497
rect 3330 397423 3386 397432
rect 3332 372564 3384 372570
rect 3332 372506 3384 372512
rect 3344 371385 3372 372506
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 3332 320136 3384 320142
rect 3332 320078 3384 320084
rect 3344 319297 3372 320078
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3332 306332 3384 306338
rect 3332 306274 3384 306280
rect 3344 306241 3372 306274
rect 3330 306232 3386 306241
rect 3330 306167 3386 306176
rect 2780 272536 2832 272542
rect 2780 272478 2832 272484
rect 2792 16574 2820 272478
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3056 202836 3108 202842
rect 3056 202778 3108 202784
rect 3068 201929 3096 202778
rect 3054 201920 3110 201929
rect 3054 201855 3110 201864
rect 3436 45529 3464 432550
rect 3528 293185 3556 432618
rect 3620 345409 3648 432686
rect 7576 423638 7604 434862
rect 7564 423632 7616 423638
rect 7564 423574 7616 423580
rect 3700 376032 3752 376038
rect 3700 375974 3752 375980
rect 3712 358465 3740 375974
rect 3698 358456 3754 358465
rect 3698 358391 3754 358400
rect 3606 345400 3662 345409
rect 3606 345335 3662 345344
rect 3514 293176 3570 293185
rect 3514 293111 3570 293120
rect 3516 267708 3568 267714
rect 3516 267650 3568 267656
rect 3528 267209 3556 267650
rect 3514 267200 3570 267209
rect 3514 267135 3570 267144
rect 7564 260160 7616 260166
rect 7564 260102 7616 260108
rect 3516 255196 3568 255202
rect 3516 255138 3568 255144
rect 3528 254153 3556 255138
rect 3514 254144 3570 254153
rect 3514 254079 3570 254088
rect 4160 249076 4212 249082
rect 4160 249018 4212 249024
rect 3516 241460 3568 241466
rect 3516 241402 3568 241408
rect 3528 241097 3556 241402
rect 3514 241088 3570 241097
rect 3514 241023 3570 241032
rect 3516 189032 3568 189038
rect 3516 188974 3568 188980
rect 3528 188873 3556 188974
rect 3514 188864 3570 188873
rect 3514 188799 3570 188808
rect 3516 150408 3568 150414
rect 3516 150350 3568 150356
rect 3528 149841 3556 150350
rect 3514 149832 3570 149841
rect 3514 149767 3570 149776
rect 3516 137964 3568 137970
rect 3516 137906 3568 137912
rect 3528 136785 3556 137906
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 3516 97980 3568 97986
rect 3516 97922 3568 97928
rect 3528 97617 3556 97922
rect 3514 97608 3570 97617
rect 3514 97543 3570 97552
rect 3516 85536 3568 85542
rect 3516 85478 3568 85484
rect 3528 84697 3556 85478
rect 3514 84688 3570 84697
rect 3514 84623 3570 84632
rect 3516 71732 3568 71738
rect 3516 71674 3568 71680
rect 3528 71641 3556 71674
rect 3514 71632 3570 71641
rect 3514 71567 3570 71576
rect 3516 59356 3568 59362
rect 3516 59298 3568 59304
rect 3528 58585 3556 59298
rect 3514 58576 3570 58585
rect 3514 58511 3570 58520
rect 3422 45520 3478 45529
rect 3422 45455 3478 45464
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 4172 16574 4200 249018
rect 6920 246356 6972 246362
rect 6920 246298 6972 246304
rect 6932 16574 6960 246298
rect 2792 16546 2912 16574
rect 4172 16546 5304 16574
rect 6932 16546 7512 16574
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 1688 480 1716 3538
rect 2884 480 2912 16546
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 4068 3868 4120 3874
rect 4068 3810 4120 3816
rect 4080 480 4108 3810
rect 5276 480 5304 16546
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 7484 3482 7512 16546
rect 7576 3874 7604 260102
rect 8956 255202 8984 436086
rect 14464 373108 14516 373114
rect 14464 373050 14516 373056
rect 12440 286340 12492 286346
rect 12440 286282 12492 286288
rect 9680 260228 9732 260234
rect 9680 260170 9732 260176
rect 8944 255196 8996 255202
rect 8944 255138 8996 255144
rect 8300 251864 8352 251870
rect 8300 251806 8352 251812
rect 8312 16574 8340 251806
rect 8312 16546 8800 16574
rect 7564 3868 7616 3874
rect 7564 3810 7616 3816
rect 6472 480 6500 3470
rect 7484 3454 7696 3482
rect 7668 480 7696 3454
rect 8772 480 8800 16546
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 260170
rect 11060 250504 11112 250510
rect 11060 250446 11112 250452
rect 11072 16574 11100 250446
rect 12452 16574 12480 286282
rect 13084 279472 13136 279478
rect 13084 279414 13136 279420
rect 11072 16546 11192 16574
rect 12452 16546 13032 16574
rect 11164 480 11192 16546
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 12360 480 12388 3538
rect 13004 3482 13032 16546
rect 13096 3602 13124 279414
rect 14476 3670 14504 373050
rect 14568 241466 14596 436154
rect 25502 430808 25558 430817
rect 25502 430743 25558 430752
rect 22744 290488 22796 290494
rect 22744 290430 22796 290436
rect 17960 269816 18012 269822
rect 17960 269758 18012 269764
rect 16580 262880 16632 262886
rect 16580 262822 16632 262828
rect 14556 241460 14608 241466
rect 14556 241402 14608 241408
rect 16592 16574 16620 262822
rect 16592 16546 17080 16574
rect 14464 3664 14516 3670
rect 14464 3606 14516 3612
rect 14740 3664 14792 3670
rect 14740 3606 14792 3612
rect 13084 3596 13136 3602
rect 13084 3538 13136 3544
rect 13004 3454 13584 3482
rect 13556 480 13584 3454
rect 14752 480 14780 3606
rect 15936 3596 15988 3602
rect 15936 3538 15988 3544
rect 15948 480 15976 3538
rect 17052 480 17080 16546
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 269758
rect 22100 257372 22152 257378
rect 22100 257314 22152 257320
rect 19340 251932 19392 251938
rect 19340 251874 19392 251880
rect 19352 16574 19380 251874
rect 20720 247716 20772 247722
rect 20720 247658 20772 247664
rect 20732 16574 20760 247658
rect 22112 16574 22140 257314
rect 19352 16546 19472 16574
rect 20732 16546 21864 16574
rect 22112 16546 22600 16574
rect 19444 480 19472 16546
rect 20628 2916 20680 2922
rect 20628 2858 20680 2864
rect 20640 480 20668 2858
rect 21836 480 21864 16546
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 22756 2922 22784 290430
rect 23480 253224 23532 253230
rect 23480 253166 23532 253172
rect 23492 16574 23520 253166
rect 25516 59362 25544 430743
rect 32402 300112 32458 300121
rect 32402 300047 32458 300056
rect 31760 283620 31812 283626
rect 31760 283562 31812 283568
rect 25596 261520 25648 261526
rect 25596 261462 25648 261468
rect 25504 59356 25556 59362
rect 25504 59298 25556 59304
rect 23492 16546 24256 16574
rect 22744 2916 22796 2922
rect 22744 2858 22796 2864
rect 24228 480 24256 16546
rect 25320 3732 25372 3738
rect 25320 3674 25372 3680
rect 25332 480 25360 3674
rect 25608 3670 25636 261462
rect 27620 260296 27672 260302
rect 27620 260238 27672 260244
rect 26240 252000 26292 252006
rect 26240 251942 26292 251948
rect 25596 3664 25648 3670
rect 25596 3606 25648 3612
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 251942
rect 27632 6914 27660 260238
rect 30380 256080 30432 256086
rect 30380 256022 30432 256028
rect 27712 256012 27764 256018
rect 27712 255954 27764 255960
rect 27724 16574 27752 255954
rect 30392 16574 30420 256022
rect 31772 16574 31800 283562
rect 27724 16546 28488 16574
rect 30392 16546 30880 16574
rect 31772 16546 31984 16574
rect 27632 6886 27752 6914
rect 27724 480 27752 6886
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28460 354 28488 16546
rect 30104 3052 30156 3058
rect 30104 2994 30156 3000
rect 30116 480 30144 2994
rect 28878 354 28990 480
rect 28460 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 32416 3058 32444 300047
rect 64880 293276 64932 293282
rect 64880 293218 64932 293224
rect 39304 287700 39356 287706
rect 39304 287642 39356 287648
rect 38660 257508 38712 257514
rect 38660 257450 38712 257456
rect 35900 257440 35952 257446
rect 35900 257382 35952 257388
rect 34520 256148 34572 256154
rect 34520 256090 34572 256096
rect 33600 3664 33652 3670
rect 33600 3606 33652 3612
rect 32404 3052 32456 3058
rect 32404 2994 32456 3000
rect 33612 480 33640 3606
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 256090
rect 35912 6914 35940 257382
rect 35992 244928 36044 244934
rect 35992 244870 36044 244876
rect 36004 16574 36032 244870
rect 38672 16574 38700 257450
rect 36004 16546 36768 16574
rect 38672 16546 39160 16574
rect 35912 6886 36032 6914
rect 36004 480 36032 6886
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 38384 3392 38436 3398
rect 38384 3334 38436 3340
rect 38396 480 38424 3334
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 39316 3398 39344 287642
rect 44180 282192 44232 282198
rect 44180 282134 44232 282140
rect 39396 273964 39448 273970
rect 39396 273906 39448 273912
rect 39408 3670 39436 273906
rect 40040 265668 40092 265674
rect 40040 265610 40092 265616
rect 40052 16574 40080 265610
rect 42800 257576 42852 257582
rect 42800 257518 42852 257524
rect 41420 256216 41472 256222
rect 41420 256158 41472 256164
rect 41432 16574 41460 256158
rect 40052 16546 40264 16574
rect 41432 16546 41920 16574
rect 39396 3664 39448 3670
rect 39396 3606 39448 3612
rect 39304 3392 39356 3398
rect 39304 3334 39356 3340
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 41892 480 41920 16546
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 257518
rect 44192 16574 44220 282134
rect 45560 279540 45612 279546
rect 45560 279482 45612 279488
rect 45572 16574 45600 279482
rect 63500 267028 63552 267034
rect 63500 266970 63552 266976
rect 60740 265736 60792 265742
rect 60740 265678 60792 265684
rect 46204 264240 46256 264246
rect 46204 264182 46256 264188
rect 44192 16546 45048 16574
rect 45572 16546 46152 16574
rect 44272 4140 44324 4146
rect 44272 4082 44324 4088
rect 44284 480 44312 4082
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45020 354 45048 16546
rect 46124 3482 46152 16546
rect 46216 4146 46244 264182
rect 52460 262948 52512 262954
rect 52460 262890 52512 262896
rect 49700 261588 49752 261594
rect 49700 261530 49752 261536
rect 48320 249144 48372 249150
rect 48320 249086 48372 249092
rect 46940 244996 46992 245002
rect 46940 244938 46992 244944
rect 46952 16574 46980 244938
rect 48332 16574 48360 249086
rect 49712 16574 49740 261530
rect 51080 246424 51132 246430
rect 51080 246366 51132 246372
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 49712 16546 50200 16574
rect 46204 4140 46256 4146
rect 46204 4082 46256 4088
rect 46124 3454 46704 3482
rect 46676 480 46704 3454
rect 45438 354 45550 480
rect 45020 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50172 480 50200 16546
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51092 354 51120 246366
rect 52472 16574 52500 262890
rect 55220 250572 55272 250578
rect 55220 250514 55272 250520
rect 53840 246492 53892 246498
rect 53840 246434 53892 246440
rect 53852 16574 53880 246434
rect 55232 16574 55260 250514
rect 56600 249212 56652 249218
rect 56600 249154 56652 249160
rect 56612 16574 56640 249154
rect 57980 247784 58032 247790
rect 57980 247726 58032 247732
rect 57992 16574 58020 247726
rect 59360 246560 59412 246566
rect 59360 246502 59412 246508
rect 52472 16546 53328 16574
rect 53852 16546 54984 16574
rect 55232 16546 56088 16574
rect 56612 16546 56824 16574
rect 57992 16546 58480 16574
rect 52552 3664 52604 3670
rect 52552 3606 52604 3612
rect 52564 480 52592 3606
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53300 354 53328 16546
rect 54956 480 54984 16546
rect 56060 480 56088 16546
rect 53718 354 53830 480
rect 53300 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 58452 480 58480 16546
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 246502
rect 60752 6914 60780 265678
rect 62120 253292 62172 253298
rect 62120 253234 62172 253240
rect 60832 249280 60884 249286
rect 60832 249222 60884 249228
rect 60844 16574 60872 249222
rect 62132 16574 62160 253234
rect 63512 16574 63540 266970
rect 64892 16574 64920 293218
rect 71044 287768 71096 287774
rect 71044 287710 71096 287716
rect 66260 272604 66312 272610
rect 66260 272546 66312 272552
rect 66272 16574 66300 272546
rect 70400 265804 70452 265810
rect 70400 265746 70452 265752
rect 69020 253360 69072 253366
rect 69020 253302 69072 253308
rect 67640 247852 67692 247858
rect 67640 247794 67692 247800
rect 60844 16546 61608 16574
rect 62132 16546 63264 16574
rect 63512 16546 64368 16574
rect 64892 16546 65104 16574
rect 66272 16546 66760 16574
rect 60752 6886 60872 6914
rect 60844 480 60872 6886
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61580 354 61608 16546
rect 63236 480 63264 16546
rect 64340 480 64368 16546
rect 61998 354 62110 480
rect 61580 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66732 480 66760 16546
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 247794
rect 69032 16574 69060 253302
rect 70412 16574 70440 265746
rect 69032 16546 69888 16574
rect 70412 16546 70992 16574
rect 69112 3800 69164 3806
rect 69112 3742 69164 3748
rect 69124 480 69152 3742
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 16546
rect 70964 3482 70992 16546
rect 71056 3806 71084 287710
rect 84200 276752 84252 276758
rect 84200 276694 84252 276700
rect 71780 276684 71832 276690
rect 71780 276626 71832 276632
rect 71792 16574 71820 276626
rect 81440 271176 81492 271182
rect 81440 271118 81492 271124
rect 74540 264308 74592 264314
rect 74540 264250 74592 264256
rect 73160 254584 73212 254590
rect 73160 254526 73212 254532
rect 73172 16574 73200 254526
rect 74552 16574 74580 264250
rect 80060 256284 80112 256290
rect 80060 256226 80112 256232
rect 77300 254652 77352 254658
rect 77300 254594 77352 254600
rect 75920 250640 75972 250646
rect 75920 250582 75972 250588
rect 71792 16546 72648 16574
rect 73172 16546 73384 16574
rect 74552 16546 75040 16574
rect 71044 3800 71096 3806
rect 71044 3742 71096 3748
rect 70964 3454 71544 3482
rect 71516 480 71544 3454
rect 72620 480 72648 16546
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 16546
rect 75012 480 75040 16546
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 250582
rect 77312 6914 77340 254594
rect 78680 252068 78732 252074
rect 78680 252010 78732 252016
rect 77392 250708 77444 250714
rect 77392 250650 77444 250656
rect 77404 16574 77432 250650
rect 78692 16574 78720 252010
rect 80072 16574 80100 256226
rect 81452 16574 81480 271118
rect 82820 253428 82872 253434
rect 82820 253370 82872 253376
rect 82832 16574 82860 253370
rect 77404 16546 78168 16574
rect 78692 16546 79272 16574
rect 80072 16546 80928 16574
rect 81452 16546 81664 16574
rect 82832 16546 83320 16574
rect 77312 6886 77432 6914
rect 77404 480 77432 6886
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78140 354 78168 16546
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 79244 354 79272 16546
rect 80900 480 80928 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83292 480 83320 16546
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 276694
rect 85580 274032 85632 274038
rect 85580 273974 85632 273980
rect 85592 6914 85620 273974
rect 88340 272672 88392 272678
rect 88340 272614 88392 272620
rect 85672 261656 85724 261662
rect 85672 261598 85724 261604
rect 85684 16574 85712 261598
rect 86960 252136 87012 252142
rect 86960 252078 87012 252084
rect 86972 16574 87000 252078
rect 88352 16574 88380 272614
rect 85684 16546 86448 16574
rect 86972 16546 87552 16574
rect 88352 16546 88932 16574
rect 85592 6886 85712 6914
rect 85684 480 85712 6886
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86420 354 86448 16546
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 87524 354 87552 16546
rect 88904 3482 88932 16546
rect 88996 6866 89024 436222
rect 98644 435260 98696 435266
rect 98644 435202 98696 435208
rect 94504 434240 94556 434246
rect 94504 434182 94556 434188
rect 94516 306338 94544 434182
rect 97908 432540 97960 432546
rect 97908 432482 97960 432488
rect 97724 371544 97776 371550
rect 97724 371486 97776 371492
rect 97736 362001 97764 371486
rect 97816 371476 97868 371482
rect 97816 371418 97868 371424
rect 97828 364721 97856 371418
rect 97814 364712 97870 364721
rect 97814 364647 97870 364656
rect 97722 361992 97778 362001
rect 97722 361927 97778 361936
rect 97814 356552 97870 356561
rect 97814 356487 97870 356496
rect 97722 345672 97778 345681
rect 97722 345607 97778 345616
rect 97630 340232 97686 340241
rect 97630 340167 97686 340176
rect 97538 332072 97594 332081
rect 97538 332007 97594 332016
rect 97446 326632 97502 326641
rect 97446 326567 97502 326576
rect 97354 315752 97410 315761
rect 97354 315687 97410 315696
rect 97262 310312 97318 310321
rect 97262 310247 97318 310256
rect 94504 306332 94556 306338
rect 94504 306274 94556 306280
rect 97172 305244 97224 305250
rect 97172 305186 97224 305192
rect 97184 299441 97212 305186
rect 97276 300762 97304 310247
rect 97264 300756 97316 300762
rect 97264 300698 97316 300704
rect 97368 300286 97396 315687
rect 97460 300830 97488 326567
rect 97552 305250 97580 332007
rect 97540 305244 97592 305250
rect 97540 305186 97592 305192
rect 97540 305108 97592 305114
rect 97540 305050 97592 305056
rect 97448 300824 97500 300830
rect 97448 300766 97500 300772
rect 97356 300280 97408 300286
rect 97356 300222 97408 300228
rect 97170 299432 97226 299441
rect 97170 299367 97226 299376
rect 97552 299305 97580 305050
rect 97644 300422 97672 340167
rect 97736 300626 97764 345607
rect 97828 305114 97856 356487
rect 97920 351121 97948 432482
rect 97906 351112 97962 351121
rect 97906 351047 97962 351056
rect 97906 348392 97962 348401
rect 97906 348327 97962 348336
rect 97816 305108 97868 305114
rect 97816 305050 97868 305056
rect 97920 304994 97948 348327
rect 98550 321192 98606 321201
rect 98550 321127 98606 321136
rect 97828 304966 97948 304994
rect 97724 300620 97776 300626
rect 97724 300562 97776 300568
rect 97828 300558 97856 304966
rect 97906 304872 97962 304881
rect 97906 304807 97962 304816
rect 97816 300552 97868 300558
rect 97816 300494 97868 300500
rect 97632 300416 97684 300422
rect 97632 300358 97684 300364
rect 97920 299470 97948 304807
rect 97908 299464 97960 299470
rect 97908 299406 97960 299412
rect 97538 299296 97594 299305
rect 98564 299266 98592 321127
rect 98656 320142 98684 435202
rect 100024 434988 100076 434994
rect 100024 434930 100076 434936
rect 100036 372570 100064 434930
rect 196624 432336 196676 432342
rect 196624 432278 196676 432284
rect 140780 432268 140832 432274
rect 140780 432210 140832 432216
rect 140792 383654 140820 432210
rect 140792 383626 141464 383654
rect 121276 374876 121328 374882
rect 121276 374818 121328 374824
rect 108396 374808 108448 374814
rect 108396 374750 108448 374756
rect 100668 372836 100720 372842
rect 100668 372778 100720 372784
rect 100024 372564 100076 372570
rect 100024 372506 100076 372512
rect 100680 372028 100708 372778
rect 103244 372700 103296 372706
rect 103244 372642 103296 372648
rect 103256 372028 103284 372642
rect 108408 372028 108436 374750
rect 116124 374536 116176 374542
rect 116124 374478 116176 374484
rect 110972 374468 111024 374474
rect 110972 374410 111024 374416
rect 110984 372028 111012 374410
rect 113548 374128 113600 374134
rect 113548 374070 113600 374076
rect 113560 372028 113588 374070
rect 116136 372028 116164 374478
rect 121288 372028 121316 374818
rect 131580 374740 131632 374746
rect 131580 374682 131632 374688
rect 129004 374196 129056 374202
rect 129004 374138 129056 374144
rect 126428 372904 126480 372910
rect 126428 372846 126480 372852
rect 126440 372028 126468 372846
rect 129016 372028 129044 374138
rect 131592 372028 131620 374682
rect 139308 374604 139360 374610
rect 139308 374546 139360 374552
rect 136732 373040 136784 373046
rect 136732 372982 136784 372988
rect 134154 372736 134210 372745
rect 134154 372671 134210 372680
rect 134168 372028 134196 372671
rect 136744 372028 136772 372982
rect 139320 372028 139348 374546
rect 141436 372042 141464 383626
rect 167644 374944 167696 374950
rect 167644 374886 167696 374892
rect 174636 374944 174688 374950
rect 174636 374886 174688 374892
rect 147036 374672 147088 374678
rect 147036 374614 147088 374620
rect 144460 372972 144512 372978
rect 144460 372914 144512 372920
rect 141436 372014 141910 372042
rect 144472 372028 144500 372914
rect 147048 372028 147076 374614
rect 165528 374400 165580 374406
rect 165528 374342 165580 374348
rect 162492 374332 162544 374338
rect 162492 374274 162544 374280
rect 157340 374264 157392 374270
rect 157340 374206 157392 374212
rect 152188 372768 152240 372774
rect 152188 372710 152240 372716
rect 149612 372632 149664 372638
rect 149612 372574 149664 372580
rect 149624 372028 149652 372574
rect 152200 372028 152228 372710
rect 157352 372028 157380 374206
rect 159914 374096 159970 374105
rect 159914 374031 159970 374040
rect 159928 372028 159956 374031
rect 162504 372028 162532 374274
rect 165540 373114 165568 374342
rect 165068 373108 165120 373114
rect 165068 373050 165120 373056
rect 165528 373108 165580 373114
rect 165528 373050 165580 373056
rect 165080 372028 165108 373050
rect 167656 372028 167684 374886
rect 170772 374876 170824 374882
rect 170772 374818 170824 374824
rect 170404 374672 170456 374678
rect 170404 374614 170456 374620
rect 99840 371816 99892 371822
rect 99840 371758 99892 371764
rect 99852 367985 99880 371758
rect 154790 371754 155080 371770
rect 154790 371748 155092 371754
rect 154790 371742 155040 371748
rect 155040 371690 155092 371696
rect 170036 371748 170088 371754
rect 170036 371690 170088 371696
rect 118330 371648 118386 371657
rect 105846 371618 106136 371634
rect 105846 371612 106148 371618
rect 105846 371606 106096 371612
rect 119066 371648 119122 371657
rect 118726 371618 119016 371634
rect 118726 371612 119028 371618
rect 118726 371606 118976 371612
rect 118330 371583 118332 371592
rect 106096 371554 106148 371560
rect 118384 371583 118386 371592
rect 118332 371554 118384 371560
rect 123878 371618 124168 371634
rect 123878 371612 124180 371618
rect 123878 371606 124128 371612
rect 119066 371583 119068 371592
rect 118976 371554 119028 371560
rect 119120 371583 119122 371592
rect 119068 371554 119120 371560
rect 124128 371554 124180 371560
rect 169602 371470 169984 371498
rect 99838 367976 99894 367985
rect 169956 367946 169984 371470
rect 170048 371346 170076 371690
rect 170036 371340 170088 371346
rect 170036 371282 170088 371288
rect 99838 367911 99894 367920
rect 169944 367940 169996 367946
rect 169944 367882 169996 367888
rect 99286 359272 99342 359281
rect 99286 359207 99342 359216
rect 99194 353832 99250 353841
rect 99194 353767 99250 353776
rect 99102 342952 99158 342961
rect 99102 342887 99158 342896
rect 99010 337512 99066 337521
rect 99010 337447 99066 337456
rect 98918 329352 98974 329361
rect 98918 329287 98974 329296
rect 98826 323912 98882 323921
rect 98826 323847 98882 323856
rect 98644 320136 98696 320142
rect 98644 320078 98696 320084
rect 98734 318472 98790 318481
rect 98734 318407 98790 318416
rect 98642 307592 98698 307601
rect 98642 307527 98698 307536
rect 98656 299402 98684 307527
rect 98644 299396 98696 299402
rect 98644 299338 98696 299344
rect 97538 299231 97594 299240
rect 98552 299260 98604 299266
rect 98552 299202 98604 299208
rect 98748 297158 98776 318407
rect 98840 299334 98868 323847
rect 98932 300082 98960 329287
rect 99024 300490 99052 337447
rect 99012 300484 99064 300490
rect 99012 300426 99064 300432
rect 98920 300076 98972 300082
rect 98920 300018 98972 300024
rect 98828 299328 98880 299334
rect 98828 299270 98880 299276
rect 98736 297152 98788 297158
rect 98736 297094 98788 297100
rect 99116 296682 99144 342887
rect 99208 300150 99236 353767
rect 99300 300801 99328 359207
rect 99378 334792 99434 334801
rect 99378 334727 99434 334736
rect 99286 300792 99342 300801
rect 99286 300727 99342 300736
rect 99392 300694 99420 334727
rect 99470 313032 99526 313041
rect 99470 312967 99526 312976
rect 99380 300688 99432 300694
rect 99380 300630 99432 300636
rect 99484 300354 99512 312967
rect 170416 307358 170444 374614
rect 170680 373040 170732 373046
rect 170680 372982 170732 372988
rect 170588 372632 170640 372638
rect 170588 372574 170640 372580
rect 170496 367940 170548 367946
rect 170496 367882 170548 367888
rect 170508 309194 170536 367882
rect 170496 309188 170548 309194
rect 170496 309130 170548 309136
rect 170600 308650 170628 372574
rect 170588 308644 170640 308650
rect 170588 308586 170640 308592
rect 170692 308446 170720 372982
rect 170784 309777 170812 374818
rect 171876 374740 171928 374746
rect 171876 374682 171928 374688
rect 170864 374604 170916 374610
rect 170864 374546 170916 374552
rect 170876 311166 170904 374546
rect 170956 374468 171008 374474
rect 170956 374410 171008 374416
rect 170864 311160 170916 311166
rect 170864 311102 170916 311108
rect 170770 309768 170826 309777
rect 170770 309703 170826 309712
rect 170968 309369 170996 374410
rect 171782 350432 171838 350441
rect 171782 350367 171838 350376
rect 171322 323232 171378 323241
rect 171322 323167 171378 323176
rect 171336 322998 171364 323167
rect 171324 322992 171376 322998
rect 171324 322934 171376 322940
rect 171506 320512 171562 320521
rect 171506 320447 171562 320456
rect 171520 320210 171548 320447
rect 171508 320204 171560 320210
rect 171508 320146 171560 320152
rect 171506 317792 171562 317801
rect 171506 317727 171562 317736
rect 171520 317490 171548 317727
rect 171508 317484 171560 317490
rect 171508 317426 171560 317432
rect 170954 309360 171010 309369
rect 170954 309295 171010 309304
rect 171796 309126 171824 350367
rect 171784 309120 171836 309126
rect 171784 309062 171836 309068
rect 170680 308440 170732 308446
rect 170680 308382 170732 308388
rect 170404 307352 170456 307358
rect 170404 307294 170456 307300
rect 170496 307284 170548 307290
rect 170496 307226 170548 307232
rect 169944 306196 169996 306202
rect 169944 306138 169996 306144
rect 169852 304496 169904 304502
rect 169852 304438 169904 304444
rect 99838 302152 99894 302161
rect 99838 302087 99894 302096
rect 99472 300348 99524 300354
rect 99472 300290 99524 300296
rect 99852 300218 99880 302087
rect 169758 301744 169814 301753
rect 169680 301702 169758 301730
rect 166630 300656 166686 300665
rect 166382 300614 166630 300642
rect 169680 300642 169708 301702
rect 169758 301679 169814 301688
rect 169864 300665 169892 304438
rect 168958 300614 169708 300642
rect 169850 300656 169906 300665
rect 166630 300591 166686 300600
rect 169850 300591 169906 300600
rect 168378 300384 168434 300393
rect 168378 300319 168434 300328
rect 160098 300248 160154 300257
rect 99840 300212 99892 300218
rect 160098 300183 160154 300192
rect 99840 300154 99892 300160
rect 99196 300144 99248 300150
rect 99196 300086 99248 300092
rect 100036 297702 100064 300084
rect 100024 297696 100076 297702
rect 100024 297638 100076 297644
rect 101968 297090 101996 300084
rect 104544 299198 104572 300084
rect 104532 299192 104584 299198
rect 104532 299134 104584 299140
rect 107120 297634 107148 300084
rect 107108 297628 107160 297634
rect 107108 297570 107160 297576
rect 109696 297566 109724 300084
rect 109684 297560 109736 297566
rect 109684 297502 109736 297508
rect 112272 297498 112300 300084
rect 114848 299130 114876 300084
rect 117332 300070 117438 300098
rect 114836 299124 114888 299130
rect 114836 299066 114888 299072
rect 112260 297492 112312 297498
rect 112260 297434 112312 297440
rect 101956 297084 102008 297090
rect 101956 297026 102008 297032
rect 99104 296676 99156 296682
rect 99104 296618 99156 296624
rect 117332 296614 117360 300070
rect 120000 299062 120028 300084
rect 119988 299056 120040 299062
rect 119988 298998 120040 299004
rect 122576 297906 122604 300084
rect 125152 298994 125180 300084
rect 126992 300070 127742 300098
rect 125140 298988 125192 298994
rect 125140 298930 125192 298936
rect 122564 297900 122616 297906
rect 122564 297842 122616 297848
rect 117320 296608 117372 296614
rect 117320 296550 117372 296556
rect 126992 296546 127020 300070
rect 130304 297770 130332 300084
rect 132880 297974 132908 300084
rect 132868 297968 132920 297974
rect 132868 297910 132920 297916
rect 130292 297764 130344 297770
rect 130292 297706 130344 297712
rect 135456 297430 135484 300084
rect 138032 297838 138060 300084
rect 140608 298926 140636 300084
rect 140596 298920 140648 298926
rect 140596 298862 140648 298868
rect 138020 297832 138072 297838
rect 138020 297774 138072 297780
rect 135444 297424 135496 297430
rect 135444 297366 135496 297372
rect 143184 297362 143212 300084
rect 145760 298722 145788 300084
rect 146944 298784 146996 298790
rect 146944 298726 146996 298732
rect 145748 298716 145800 298722
rect 145748 298658 145800 298664
rect 146956 297770 146984 298726
rect 148336 297770 148364 300084
rect 150912 297945 150940 300084
rect 153212 300070 153502 300098
rect 150898 297936 150954 297945
rect 150898 297871 150954 297880
rect 146944 297764 146996 297770
rect 146944 297706 146996 297712
rect 148324 297764 148376 297770
rect 148324 297706 148376 297712
rect 143172 297356 143224 297362
rect 143172 297298 143224 297304
rect 126980 296540 127032 296546
rect 126980 296482 127032 296488
rect 153212 296478 153240 300070
rect 156064 298858 156092 300084
rect 156052 298852 156104 298858
rect 156052 298794 156104 298800
rect 158640 298110 158668 300084
rect 158628 298104 158680 298110
rect 158628 298046 158680 298052
rect 153200 296472 153252 296478
rect 153200 296414 153252 296420
rect 149060 296132 149112 296138
rect 149060 296074 149112 296080
rect 143540 296064 143592 296070
rect 143540 296006 143592 296012
rect 125600 295996 125652 296002
rect 125600 295938 125652 295944
rect 103520 284980 103572 284986
rect 103520 284922 103572 284928
rect 102140 279608 102192 279614
rect 102140 279550 102192 279556
rect 99380 269884 99432 269890
rect 99380 269826 99432 269832
rect 95240 268456 95292 268462
rect 95240 268398 95292 268404
rect 92480 268388 92532 268394
rect 92480 268330 92532 268336
rect 91100 254720 91152 254726
rect 91100 254662 91152 254668
rect 89720 249348 89772 249354
rect 89720 249290 89772 249296
rect 89732 16574 89760 249290
rect 91112 16574 91140 254662
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 88984 6860 89036 6866
rect 88984 6802 89036 6808
rect 88904 3454 89208 3482
rect 89180 480 89208 3454
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 268330
rect 93860 258732 93912 258738
rect 93860 258674 93912 258680
rect 93872 3398 93900 258674
rect 93952 254788 94004 254794
rect 93952 254730 94004 254736
rect 93860 3392 93912 3398
rect 93860 3334 93912 3340
rect 93964 480 93992 254730
rect 95252 16574 95280 268398
rect 98000 261724 98052 261730
rect 98000 261666 98052 261672
rect 96620 257644 96672 257650
rect 96620 257586 96672 257592
rect 96632 16574 96660 257586
rect 98012 16574 98040 261666
rect 99392 16574 99420 269826
rect 100760 264376 100812 264382
rect 100760 264318 100812 264324
rect 95252 16546 95832 16574
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 94780 3392 94832 3398
rect 94780 3334 94832 3340
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94792 354 94820 3334
rect 95118 354 95230 480
rect 94792 326 95230 354
rect 95804 354 95832 16546
rect 97460 480 97488 16546
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 264318
rect 102152 6914 102180 279550
rect 102232 254856 102284 254862
rect 102232 254798 102284 254804
rect 102244 16574 102272 254798
rect 103532 16574 103560 284922
rect 111800 283688 111852 283694
rect 111800 283630 111852 283636
rect 110420 280832 110472 280838
rect 110420 280774 110472 280780
rect 106280 276820 106332 276826
rect 106280 276762 106332 276768
rect 104900 263016 104952 263022
rect 104900 262958 104952 262964
rect 104912 16574 104940 262958
rect 106292 16574 106320 276762
rect 107660 269952 107712 269958
rect 107660 269894 107712 269900
rect 107672 16574 107700 269894
rect 109040 245064 109092 245070
rect 109040 245006 109092 245012
rect 102244 16546 103376 16574
rect 103532 16546 104112 16574
rect 104912 16546 105768 16574
rect 106292 16546 106504 16574
rect 107672 16546 108160 16574
rect 102152 6886 102272 6914
rect 102244 480 102272 6886
rect 103348 480 103376 16546
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105740 480 105768 16546
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108132 480 108160 16546
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109052 354 109080 245006
rect 110432 3398 110460 280774
rect 110512 260364 110564 260370
rect 110512 260306 110564 260312
rect 110420 3392 110472 3398
rect 110420 3334 110472 3340
rect 110524 480 110552 260306
rect 111812 16574 111840 283630
rect 117320 278044 117372 278050
rect 117320 277986 117372 277992
rect 115940 268524 115992 268530
rect 115940 268466 115992 268472
rect 114560 267096 114612 267102
rect 114560 267038 114612 267044
rect 113180 263084 113232 263090
rect 113180 263026 113232 263032
rect 113192 16574 113220 263026
rect 114572 16574 114600 267038
rect 115952 16574 115980 268466
rect 111812 16546 112392 16574
rect 113192 16546 114048 16574
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 111616 3392 111668 3398
rect 111616 3334 111668 3340
rect 111628 480 111656 3334
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114020 480 114048 16546
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 277986
rect 124220 270020 124272 270026
rect 124220 269962 124272 269968
rect 122840 267164 122892 267170
rect 122840 267106 122892 267112
rect 121460 253564 121512 253570
rect 121460 253506 121512 253512
rect 118700 253496 118752 253502
rect 118700 253438 118752 253444
rect 118712 6914 118740 253438
rect 118792 246628 118844 246634
rect 118792 246570 118844 246576
rect 118804 16574 118832 246570
rect 120080 245132 120132 245138
rect 120080 245074 120132 245080
rect 120092 16574 120120 245074
rect 121472 16574 121500 253506
rect 122852 16574 122880 267106
rect 124232 16574 124260 269962
rect 118804 16546 119936 16574
rect 120092 16546 120672 16574
rect 121472 16546 122328 16574
rect 122852 16546 123064 16574
rect 124232 16546 124720 16574
rect 118712 6886 118832 6914
rect 118804 480 118832 6886
rect 119908 480 119936 16546
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 122300 480 122328 16546
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124692 480 124720 16546
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125612 354 125640 295938
rect 139400 294636 139452 294642
rect 139400 294578 139452 294584
rect 128360 291848 128412 291854
rect 128360 291790 128412 291796
rect 126980 283756 127032 283762
rect 126980 283698 127032 283704
rect 126992 480 127020 283698
rect 127072 274100 127124 274106
rect 127072 274042 127124 274048
rect 127084 16574 127112 274042
rect 128372 16574 128400 291790
rect 132500 290556 132552 290562
rect 132500 290498 132552 290504
rect 131120 282260 131172 282266
rect 131120 282202 131172 282208
rect 129740 275324 129792 275330
rect 129740 275266 129792 275272
rect 129752 16574 129780 275266
rect 131132 16574 131160 282202
rect 132512 16574 132540 290498
rect 135260 289128 135312 289134
rect 135260 289070 135312 289076
rect 133880 270088 133932 270094
rect 133880 270030 133932 270036
rect 127084 16546 128216 16574
rect 128372 16546 128952 16574
rect 129752 16546 130608 16574
rect 131132 16546 131344 16574
rect 132512 16546 133000 16574
rect 128188 480 128216 16546
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 16546
rect 130580 480 130608 16546
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 132972 480 133000 16546
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 133892 354 133920 270030
rect 135272 3806 135300 289070
rect 135352 285048 135404 285054
rect 135352 284990 135404 284996
rect 135260 3800 135312 3806
rect 135260 3742 135312 3748
rect 135364 3482 135392 284990
rect 136640 268592 136692 268598
rect 136640 268534 136692 268540
rect 136652 16574 136680 268534
rect 138020 265872 138072 265878
rect 138020 265814 138072 265820
rect 138032 16574 138060 265814
rect 139412 16574 139440 294578
rect 140780 280900 140832 280906
rect 140780 280842 140832 280848
rect 140792 16574 140820 280842
rect 142160 250776 142212 250782
rect 142160 250718 142212 250724
rect 136652 16546 137232 16574
rect 138032 16546 138888 16574
rect 139412 16546 139624 16574
rect 140792 16546 141280 16574
rect 136456 3800 136508 3806
rect 136456 3742 136508 3748
rect 135272 3454 135392 3482
rect 135272 480 135300 3454
rect 136468 480 136496 3742
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 16546
rect 138860 480 138888 16546
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 139596 354 139624 16546
rect 141252 480 141280 16546
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142172 354 142200 250718
rect 143552 480 143580 296006
rect 146300 287836 146352 287842
rect 146300 287778 146352 287784
rect 143632 271244 143684 271250
rect 143632 271186 143684 271192
rect 143644 16574 143672 271186
rect 144920 264444 144972 264450
rect 144920 264386 144972 264392
rect 144932 16574 144960 264386
rect 146312 16574 146340 287778
rect 147680 278112 147732 278118
rect 147680 278054 147732 278060
rect 147692 16574 147720 278054
rect 149072 16574 149100 296074
rect 150440 293344 150492 293350
rect 150440 293286 150492 293292
rect 150452 16574 150480 293286
rect 153200 286408 153252 286414
rect 153200 286350 153252 286356
rect 151820 276888 151872 276894
rect 151820 276830 151872 276836
rect 143644 16546 144776 16574
rect 144932 16546 145512 16574
rect 146312 16546 147168 16574
rect 147692 16546 147904 16574
rect 149072 16546 149560 16574
rect 150452 16546 150664 16574
rect 144748 480 144776 16546
rect 142406 354 142518 480
rect 142172 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 147140 480 147168 16546
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 149532 480 149560 16546
rect 150636 480 150664 16546
rect 151832 480 151860 276830
rect 151912 271312 151964 271318
rect 151912 271254 151964 271260
rect 151924 16574 151952 271254
rect 153212 16574 153240 286350
rect 157340 285116 157392 285122
rect 157340 285058 157392 285064
rect 154580 263152 154632 263158
rect 154580 263094 154632 263100
rect 154592 16574 154620 263094
rect 155960 247920 156012 247926
rect 155960 247862 156012 247868
rect 155972 16574 156000 247862
rect 157352 16574 157380 285058
rect 158720 245268 158772 245274
rect 158720 245210 158772 245216
rect 158732 16574 158760 245210
rect 151924 16546 153056 16574
rect 153212 16546 153792 16574
rect 154592 16546 155448 16574
rect 155972 16546 156184 16574
rect 157352 16546 157840 16574
rect 158732 16546 158944 16574
rect 153028 480 153056 16546
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 16546
rect 155420 480 155448 16546
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156156 354 156184 16546
rect 157812 480 157840 16546
rect 158916 480 158944 16546
rect 160112 11762 160140 300183
rect 161216 298654 161244 300084
rect 161204 298648 161256 298654
rect 161204 298590 161256 298596
rect 163792 298586 163820 300084
rect 163780 298580 163832 298586
rect 163780 298522 163832 298528
rect 164240 294704 164292 294710
rect 164240 294646 164292 294652
rect 161480 282328 161532 282334
rect 161480 282270 161532 282276
rect 160192 245336 160244 245342
rect 160192 245278 160244 245284
rect 160100 11756 160152 11762
rect 160100 11698 160152 11704
rect 160204 6914 160232 245278
rect 161492 16574 161520 282270
rect 162860 265940 162912 265946
rect 162860 265882 162912 265888
rect 162872 16574 162900 265882
rect 164252 16574 164280 294646
rect 165620 281036 165672 281042
rect 165620 280978 165672 280984
rect 165632 16574 165660 280978
rect 167000 272740 167052 272746
rect 167000 272682 167052 272688
rect 167012 16574 167040 272682
rect 161492 16546 162072 16574
rect 162872 16546 163728 16574
rect 164252 16546 164464 16574
rect 165632 16546 166120 16574
rect 167012 16546 167224 16574
rect 161296 11756 161348 11762
rect 161296 11698 161348 11704
rect 160112 6886 160232 6914
rect 160112 480 160140 6886
rect 161308 480 161336 11698
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 354 162072 16546
rect 163700 480 163728 16546
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164436 354 164464 16546
rect 166092 480 166120 16546
rect 167196 480 167224 16546
rect 168392 480 168420 300319
rect 169956 298110 169984 306138
rect 170402 305688 170458 305697
rect 170402 305623 170458 305632
rect 170036 304360 170088 304366
rect 170036 304302 170088 304308
rect 169944 298104 169996 298110
rect 169944 298046 169996 298052
rect 170048 297566 170076 304302
rect 170036 297560 170088 297566
rect 170036 297502 170088 297508
rect 168472 279676 168524 279682
rect 168472 279618 168524 279624
rect 168484 16574 168512 279618
rect 168484 16546 169616 16574
rect 169588 480 169616 16546
rect 170416 3602 170444 305623
rect 170508 297634 170536 307226
rect 171692 304428 171744 304434
rect 171692 304370 171744 304376
rect 170496 297628 170548 297634
rect 170496 297570 170548 297576
rect 171704 297430 171732 304370
rect 171692 297424 171744 297430
rect 171692 297366 171744 297372
rect 170772 3800 170824 3806
rect 170772 3742 170824 3748
rect 170404 3596 170456 3602
rect 170404 3538 170456 3544
rect 170784 480 170812 3742
rect 171796 3466 171824 309062
rect 171888 307018 171916 374682
rect 173256 374536 173308 374542
rect 173256 374478 173308 374484
rect 173164 372904 173216 372910
rect 173164 372846 173216 372852
rect 172334 369472 172390 369481
rect 172334 369407 172390 369416
rect 172348 368558 172376 369407
rect 172336 368552 172388 368558
rect 172336 368494 172388 368500
rect 171966 366752 172022 366761
rect 171966 366687 172022 366696
rect 171980 310690 172008 366687
rect 172334 364032 172390 364041
rect 172334 363967 172390 363976
rect 172348 362982 172376 363967
rect 172336 362976 172388 362982
rect 172336 362918 172388 362924
rect 172058 361312 172114 361321
rect 172058 361247 172114 361256
rect 171968 310684 172020 310690
rect 171968 310626 172020 310632
rect 172072 310622 172100 361247
rect 172426 358592 172482 358601
rect 172426 358527 172482 358536
rect 172440 357474 172468 358527
rect 172428 357468 172480 357474
rect 172428 357410 172480 357416
rect 172426 355872 172482 355881
rect 172426 355807 172482 355816
rect 172440 354754 172468 355807
rect 172428 354748 172480 354754
rect 172428 354690 172480 354696
rect 172426 353152 172482 353161
rect 172426 353087 172482 353096
rect 172440 351966 172468 353087
rect 172428 351960 172480 351966
rect 172428 351902 172480 351908
rect 172426 347712 172482 347721
rect 172426 347647 172482 347656
rect 172440 346458 172468 347647
rect 172428 346452 172480 346458
rect 172428 346394 172480 346400
rect 172150 344992 172206 345001
rect 172150 344927 172206 344936
rect 172164 310758 172192 344927
rect 172428 342304 172480 342310
rect 172426 342272 172428 342281
rect 172480 342272 172482 342281
rect 172426 342207 172482 342216
rect 172426 339552 172482 339561
rect 172426 339487 172428 339496
rect 172480 339487 172482 339496
rect 172428 339458 172480 339464
rect 172426 336832 172482 336841
rect 172426 336767 172428 336776
rect 172480 336767 172482 336776
rect 172428 336738 172480 336744
rect 172242 334112 172298 334121
rect 172242 334047 172298 334056
rect 172256 311234 172284 334047
rect 172426 331392 172482 331401
rect 172426 331327 172482 331336
rect 172440 331294 172468 331327
rect 172428 331288 172480 331294
rect 172428 331230 172480 331236
rect 172426 328672 172482 328681
rect 172426 328607 172482 328616
rect 172440 328506 172468 328607
rect 172428 328500 172480 328506
rect 172428 328442 172480 328448
rect 172334 325952 172390 325961
rect 172334 325887 172390 325896
rect 172348 311302 172376 325887
rect 172426 315072 172482 315081
rect 172426 315007 172482 315016
rect 172440 314702 172468 315007
rect 172428 314696 172480 314702
rect 172428 314638 172480 314644
rect 172426 312352 172482 312361
rect 172426 312287 172482 312296
rect 172440 311914 172468 312287
rect 172428 311908 172480 311914
rect 172428 311850 172480 311856
rect 172336 311296 172388 311302
rect 172336 311238 172388 311244
rect 172244 311228 172296 311234
rect 172244 311170 172296 311176
rect 172152 310752 172204 310758
rect 172152 310694 172204 310700
rect 172060 310616 172112 310622
rect 172060 310558 172112 310564
rect 172428 310004 172480 310010
rect 172428 309946 172480 309952
rect 172440 309641 172468 309946
rect 172426 309632 172482 309641
rect 172426 309567 172482 309576
rect 173176 308582 173204 372846
rect 173268 309505 173296 374478
rect 174544 372836 174596 372842
rect 174544 372778 174596 372784
rect 173440 371680 173492 371686
rect 173440 371622 173492 371628
rect 173348 371612 173400 371618
rect 173348 371554 173400 371560
rect 173254 309496 173310 309505
rect 173254 309431 173310 309440
rect 173164 308576 173216 308582
rect 173164 308518 173216 308524
rect 173360 308378 173388 371554
rect 173452 308961 173480 371622
rect 173624 371408 173676 371414
rect 173624 371350 173676 371356
rect 173438 308952 173494 308961
rect 173438 308887 173494 308896
rect 173636 308825 173664 371350
rect 173622 308816 173678 308825
rect 173622 308751 173678 308760
rect 174556 308553 174584 372778
rect 174648 309233 174676 374886
rect 188344 372972 188396 372978
rect 188344 372914 188396 372920
rect 182824 336796 182876 336802
rect 182824 336738 182876 336744
rect 182836 309262 182864 336738
rect 182824 309256 182876 309262
rect 174634 309224 174690 309233
rect 182824 309198 182876 309204
rect 174634 309159 174690 309168
rect 188356 308786 188384 372914
rect 188344 308780 188396 308786
rect 188344 308722 188396 308728
rect 174542 308544 174598 308553
rect 174542 308479 174598 308488
rect 173348 308372 173400 308378
rect 173348 308314 173400 308320
rect 172428 307624 172480 307630
rect 172428 307566 172480 307572
rect 171876 307012 171928 307018
rect 171876 306954 171928 306960
rect 172440 306921 172468 307566
rect 195980 307080 196032 307086
rect 195980 307022 196032 307028
rect 172426 306912 172482 306921
rect 172426 306847 172482 306856
rect 172244 305992 172296 305998
rect 172244 305934 172296 305940
rect 171876 304292 171928 304298
rect 171876 304234 171928 304240
rect 171888 3738 171916 304234
rect 171968 303000 172020 303006
rect 171968 302942 172020 302948
rect 171980 16574 172008 302942
rect 172256 297702 172284 305934
rect 175924 305652 175976 305658
rect 175924 305594 175976 305600
rect 172612 305448 172664 305454
rect 172612 305390 172664 305396
rect 172336 304972 172388 304978
rect 172336 304914 172388 304920
rect 172348 304201 172376 304914
rect 172334 304192 172390 304201
rect 172334 304127 172390 304136
rect 172336 302728 172388 302734
rect 172336 302670 172388 302676
rect 172244 297696 172296 297702
rect 172244 297638 172296 297644
rect 172348 297362 172376 302670
rect 172428 302184 172480 302190
rect 172428 302126 172480 302132
rect 172440 301481 172468 302126
rect 172426 301472 172482 301481
rect 172426 301407 172482 301416
rect 172624 297498 172652 305390
rect 175280 302932 175332 302938
rect 175280 302874 175332 302880
rect 172612 297492 172664 297498
rect 172612 297434 172664 297440
rect 172336 297356 172388 297362
rect 172336 297298 172388 297304
rect 174544 264512 174596 264518
rect 174544 264454 174596 264460
rect 173900 247988 173952 247994
rect 173900 247930 173952 247936
rect 171980 16546 172100 16574
rect 171876 3732 171928 3738
rect 171876 3674 171928 3680
rect 172072 3534 172100 16546
rect 172060 3528 172112 3534
rect 172060 3470 172112 3476
rect 171784 3460 171836 3466
rect 171784 3402 171836 3408
rect 173164 3460 173216 3466
rect 173164 3402 173216 3408
rect 171968 3324 172020 3330
rect 171968 3266 172020 3272
rect 171980 480 172008 3266
rect 173176 480 173204 3402
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 173912 354 173940 247930
rect 174556 3806 174584 264454
rect 175292 16574 175320 302874
rect 175292 16546 175504 16574
rect 174544 3800 174596 3806
rect 174544 3742 174596 3748
rect 175476 480 175504 16546
rect 175936 3330 175964 305594
rect 184204 291916 184256 291922
rect 184204 291858 184256 291864
rect 181444 279744 181496 279750
rect 181444 279686 181496 279692
rect 180800 261792 180852 261798
rect 180800 261734 180852 261740
rect 179420 258868 179472 258874
rect 179420 258810 179472 258816
rect 176660 258800 176712 258806
rect 176660 258742 176712 258748
rect 175924 3324 175976 3330
rect 175924 3266 175976 3272
rect 176672 480 176700 258742
rect 178040 246696 178092 246702
rect 178040 246638 178092 246644
rect 178052 16574 178080 246638
rect 179432 16574 179460 258810
rect 180812 16574 180840 261734
rect 178052 16546 178632 16574
rect 179432 16546 180288 16574
rect 180812 16546 181024 16574
rect 177856 4004 177908 4010
rect 177856 3946 177908 3952
rect 177868 480 177896 3946
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 180260 480 180288 16546
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 181456 4010 181484 279686
rect 183560 258936 183612 258942
rect 183560 258878 183612 258884
rect 182180 248056 182232 248062
rect 182180 247998 182232 248004
rect 181444 4004 181496 4010
rect 181444 3946 181496 3952
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 182192 354 182220 247998
rect 183572 16574 183600 258878
rect 183572 16546 183784 16574
rect 183756 480 183784 16546
rect 184216 3466 184244 291858
rect 184940 275392 184992 275398
rect 184940 275334 184992 275340
rect 184204 3460 184256 3466
rect 184204 3402 184256 3408
rect 184952 480 184980 275334
rect 194600 270156 194652 270162
rect 194600 270098 194652 270104
rect 191840 268660 191892 268666
rect 191840 268602 191892 268608
rect 187700 267232 187752 267238
rect 187700 267174 187752 267180
rect 186320 260500 186372 260506
rect 186320 260442 186372 260448
rect 185032 248124 185084 248130
rect 185032 248066 185084 248072
rect 185044 16574 185072 248066
rect 186332 16574 186360 260442
rect 187712 16574 187740 267174
rect 190460 260568 190512 260574
rect 190460 260510 190512 260516
rect 189080 249416 189132 249422
rect 189080 249358 189132 249364
rect 189092 16574 189120 249358
rect 185044 16546 186176 16574
rect 186332 16546 186912 16574
rect 187712 16546 188568 16574
rect 189092 16546 189304 16574
rect 186148 480 186176 16546
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 188540 480 188568 16546
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189276 354 189304 16546
rect 189694 354 189806 480
rect 189276 326 189806 354
rect 190472 354 190500 260510
rect 191852 16574 191880 268602
rect 193220 261860 193272 261866
rect 193220 261802 193272 261808
rect 191852 16546 192064 16574
rect 192036 480 192064 16546
rect 193232 3602 193260 261802
rect 193312 253700 193364 253706
rect 193312 253642 193364 253648
rect 193220 3596 193272 3602
rect 193220 3538 193272 3544
rect 193324 3482 193352 253642
rect 194612 16574 194640 270098
rect 195992 16574 196020 307022
rect 196636 20670 196664 432278
rect 197360 261928 197412 261934
rect 197360 261870 197412 261876
rect 196624 20664 196676 20670
rect 196624 20606 196676 20612
rect 197372 16574 197400 261870
rect 198016 97986 198044 436426
rect 199384 433492 199436 433498
rect 199384 433434 199436 433440
rect 198740 270224 198792 270230
rect 198740 270166 198792 270172
rect 198004 97980 198056 97986
rect 198004 97922 198056 97928
rect 194612 16546 195192 16574
rect 195992 16546 196848 16574
rect 197372 16546 197952 16574
rect 194416 3596 194468 3602
rect 194416 3538 194468 3544
rect 193232 3454 193352 3482
rect 193232 480 193260 3454
rect 194428 480 194456 3538
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 189694 -960 189806 326
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 196820 480 196848 16546
rect 197924 480 197952 16546
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 270166
rect 199396 202842 199424 433434
rect 200764 432404 200816 432410
rect 200764 432346 200816 432352
rect 200120 254924 200172 254930
rect 200120 254866 200172 254872
rect 199384 202836 199436 202842
rect 199384 202778 199436 202784
rect 200132 16574 200160 254866
rect 200776 85542 200804 432346
rect 201500 268728 201552 268734
rect 201500 268670 201552 268676
rect 200764 85536 200816 85542
rect 200764 85478 200816 85484
rect 200132 16546 200344 16574
rect 200316 480 200344 16546
rect 201512 11762 201540 268670
rect 201592 263220 201644 263226
rect 201592 263162 201644 263168
rect 201500 11756 201552 11762
rect 201500 11698 201552 11704
rect 201604 6914 201632 263162
rect 202880 254992 202932 254998
rect 202880 254934 202932 254940
rect 202892 16574 202920 254934
rect 203536 137970 203564 436494
rect 207664 435124 207716 435130
rect 207664 435066 207716 435072
rect 206284 432472 206336 432478
rect 206284 432414 206336 432420
rect 205640 271380 205692 271386
rect 205640 271322 205692 271328
rect 204260 264580 204312 264586
rect 204260 264522 204312 264528
rect 203524 137964 203576 137970
rect 203524 137906 203576 137912
rect 204272 16574 204300 264522
rect 204904 248192 204956 248198
rect 204904 248134 204956 248140
rect 202892 16546 203472 16574
rect 204272 16546 204852 16574
rect 202696 11756 202748 11762
rect 202696 11698 202748 11704
rect 201512 6886 201632 6914
rect 201512 480 201540 6886
rect 202708 480 202736 11698
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203444 354 203472 16546
rect 204824 3482 204852 16546
rect 204916 3670 204944 248134
rect 205652 16574 205680 271322
rect 206296 189038 206324 432414
rect 207020 256420 207072 256426
rect 207020 256362 207072 256368
rect 206284 189032 206336 189038
rect 206284 188974 206336 188980
rect 205652 16546 206232 16574
rect 204904 3664 204956 3670
rect 204904 3606 204956 3612
rect 204824 3454 205128 3482
rect 205100 480 205128 3454
rect 206204 480 206232 16546
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 256362
rect 207676 71738 207704 435066
rect 209044 433560 209096 433566
rect 209044 433502 209096 433508
rect 208400 264648 208452 264654
rect 208400 264590 208452 264596
rect 207664 71732 207716 71738
rect 207664 71674 207716 71680
rect 208412 16574 208440 264590
rect 209056 215286 209084 433502
rect 209780 271448 209832 271454
rect 209780 271390 209832 271396
rect 209044 215280 209096 215286
rect 209044 215222 209096 215228
rect 208412 16546 208624 16574
rect 208596 480 208624 16546
rect 209792 480 209820 271390
rect 209872 257712 209924 257718
rect 209872 257654 209924 257660
rect 209884 16574 209912 257654
rect 210436 150414 210464 436562
rect 217888 434042 217916 565082
rect 217980 478514 218008 700334
rect 217968 478508 218020 478514
rect 217968 478450 218020 478456
rect 218072 468654 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 219348 700460 219400 700466
rect 219348 700402 219400 700408
rect 219256 700324 219308 700330
rect 219256 700266 219308 700272
rect 219162 512816 219218 512825
rect 219162 512751 219218 512760
rect 219070 511048 219126 511057
rect 219070 510983 219126 510992
rect 218886 509960 218942 509969
rect 218886 509895 218942 509904
rect 218900 478310 218928 509895
rect 218978 508192 219034 508201
rect 218978 508127 219034 508136
rect 218888 478304 218940 478310
rect 218888 478246 218940 478252
rect 218992 472734 219020 508127
rect 218980 472728 219032 472734
rect 218980 472670 219032 472676
rect 219084 469946 219112 510983
rect 219072 469940 219124 469946
rect 219072 469882 219124 469888
rect 218060 468648 218112 468654
rect 218060 468590 218112 468596
rect 219176 443766 219204 512751
rect 219268 478582 219296 700266
rect 219256 478576 219308 478582
rect 219256 478518 219308 478524
rect 219164 443760 219216 443766
rect 219164 443702 219216 443708
rect 219360 436966 219388 700402
rect 234632 565146 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 700466 267688 703520
rect 267648 700460 267700 700466
rect 267648 700402 267700 700408
rect 283852 700398 283880 703520
rect 283840 700392 283892 700398
rect 283840 700334 283892 700340
rect 300136 700330 300164 703520
rect 332520 700330 332548 703520
rect 348804 700398 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 348792 700392 348844 700398
rect 348792 700334 348844 700340
rect 357440 700392 357492 700398
rect 357440 700334 357492 700340
rect 300124 700324 300176 700330
rect 300124 700266 300176 700272
rect 332508 700324 332560 700330
rect 332508 700266 332560 700272
rect 234620 565140 234672 565146
rect 234620 565082 234672 565088
rect 266452 478576 266504 478582
rect 266452 478518 266504 478524
rect 266360 478372 266412 478378
rect 266360 478314 266412 478320
rect 264980 478236 265032 478242
rect 264980 478178 265032 478184
rect 238482 477320 238538 477329
rect 238482 477255 238538 477264
rect 238496 476678 238524 477255
rect 242806 477184 242862 477193
rect 242806 477119 242862 477128
rect 240046 476912 240102 476921
rect 240046 476847 240102 476856
rect 241426 476912 241482 476921
rect 241426 476847 241482 476856
rect 238484 476672 238536 476678
rect 238484 476614 238536 476620
rect 237378 476368 237434 476377
rect 237378 476303 237434 476312
rect 237286 476232 237342 476241
rect 237286 476167 237342 476176
rect 237300 475454 237328 476167
rect 237288 475448 237340 475454
rect 237288 475390 237340 475396
rect 237392 474162 237420 476303
rect 240060 476202 240088 476847
rect 241440 476814 241468 476847
rect 241428 476808 241480 476814
rect 241428 476750 241480 476756
rect 242820 476746 242848 477119
rect 242808 476740 242860 476746
rect 242808 476682 242860 476688
rect 249062 476640 249118 476649
rect 249062 476575 249118 476584
rect 259274 476640 259330 476649
rect 259274 476575 259330 476584
rect 264886 476640 264942 476649
rect 264886 476575 264888 476584
rect 245474 476368 245530 476377
rect 245474 476303 245530 476312
rect 247682 476368 247738 476377
rect 247682 476303 247738 476312
rect 244186 476232 244242 476241
rect 240048 476196 240100 476202
rect 244186 476167 244242 476176
rect 240048 476138 240100 476144
rect 237380 474156 237432 474162
rect 237380 474098 237432 474104
rect 244200 438326 244228 476167
rect 245488 439890 245516 476303
rect 246302 476232 246358 476241
rect 246302 476167 246358 476176
rect 246316 452062 246344 476167
rect 246304 452056 246356 452062
rect 246304 451998 246356 452004
rect 247696 449274 247724 476303
rect 248234 476232 248290 476241
rect 248234 476167 248290 476176
rect 247684 449268 247736 449274
rect 247684 449210 247736 449216
rect 248248 441046 248276 476167
rect 249076 453490 249104 476575
rect 253846 476504 253902 476513
rect 253846 476439 253902 476448
rect 253860 476406 253888 476439
rect 253848 476400 253900 476406
rect 251086 476368 251142 476377
rect 251086 476303 251142 476312
rect 252374 476368 252430 476377
rect 253848 476342 253900 476348
rect 256606 476368 256662 476377
rect 252374 476303 252430 476312
rect 256606 476303 256662 476312
rect 249706 476232 249762 476241
rect 249706 476167 249762 476176
rect 250994 476232 251050 476241
rect 250994 476167 251050 476176
rect 249064 453484 249116 453490
rect 249064 453426 249116 453432
rect 249720 442406 249748 476167
rect 251008 460426 251036 476167
rect 250996 460420 251048 460426
rect 250996 460362 251048 460368
rect 249800 456816 249852 456822
rect 249800 456758 249852 456764
rect 249708 442400 249760 442406
rect 249708 442342 249760 442348
rect 249812 441614 249840 456758
rect 251100 456210 251128 476303
rect 252388 472802 252416 476303
rect 252466 476232 252522 476241
rect 252466 476167 252522 476176
rect 253754 476232 253810 476241
rect 253754 476167 253810 476176
rect 255226 476232 255282 476241
rect 255226 476167 255282 476176
rect 256514 476232 256570 476241
rect 256514 476167 256570 476176
rect 252376 472796 252428 472802
rect 252376 472738 252428 472744
rect 251824 470620 251876 470626
rect 251824 470562 251876 470568
rect 251180 464364 251232 464370
rect 251180 464306 251232 464312
rect 251088 456204 251140 456210
rect 251088 456146 251140 456152
rect 249812 441586 250576 441614
rect 248236 441040 248288 441046
rect 248236 440982 248288 440988
rect 245476 439884 245528 439890
rect 245476 439826 245528 439832
rect 244188 438320 244240 438326
rect 244188 438262 244240 438268
rect 219348 436960 219400 436966
rect 219348 436902 219400 436908
rect 231216 436688 231268 436694
rect 231216 436630 231268 436636
rect 225604 435192 225656 435198
rect 225604 435134 225656 435140
rect 217876 434036 217928 434042
rect 217876 433978 217928 433984
rect 220084 351960 220136 351966
rect 220084 351902 220136 351908
rect 220096 307562 220124 351902
rect 224224 346452 224276 346458
rect 224224 346394 224276 346400
rect 222292 310684 222344 310690
rect 222292 310626 222344 310632
rect 222304 310350 222332 310626
rect 222292 310344 222344 310350
rect 222292 310286 222344 310292
rect 220084 307556 220136 307562
rect 220084 307498 220136 307504
rect 224236 307426 224264 346394
rect 224224 307420 224276 307426
rect 224224 307362 224276 307368
rect 215208 307216 215260 307222
rect 215208 307158 215260 307164
rect 210976 307148 211028 307154
rect 210976 307090 211028 307096
rect 210884 295248 210936 295254
rect 210884 295190 210936 295196
rect 210896 193186 210924 295190
rect 210884 193180 210936 193186
rect 210884 193122 210936 193128
rect 210988 189038 211016 307090
rect 214932 306060 214984 306066
rect 214932 306002 214984 306008
rect 213828 305788 213880 305794
rect 213828 305730 213880 305736
rect 212080 305720 212132 305726
rect 212080 305662 212132 305668
rect 211988 301572 212040 301578
rect 211988 301514 212040 301520
rect 211894 300520 211950 300529
rect 211894 300455 211950 300464
rect 211802 297664 211858 297673
rect 211712 297628 211764 297634
rect 211802 297599 211858 297608
rect 211712 297570 211764 297576
rect 211066 297392 211122 297401
rect 211066 297327 211122 297336
rect 210976 189032 211028 189038
rect 210976 188974 211028 188980
rect 211080 155582 211108 297327
rect 211620 294840 211672 294846
rect 211620 294782 211672 294788
rect 211632 158030 211660 294782
rect 211620 158024 211672 158030
rect 211620 157966 211672 157972
rect 211068 155576 211120 155582
rect 211068 155518 211120 155524
rect 211724 155514 211752 297570
rect 211816 155718 211844 297599
rect 211908 158506 211936 300455
rect 212000 158778 212028 301514
rect 212092 159934 212120 305662
rect 213460 303136 213512 303142
rect 213460 303078 213512 303084
rect 212448 303068 212500 303074
rect 212448 303010 212500 303016
rect 212354 297800 212410 297809
rect 212354 297735 212410 297744
rect 212170 297528 212226 297537
rect 212170 297463 212226 297472
rect 212080 159928 212132 159934
rect 212080 159870 212132 159876
rect 211988 158772 212040 158778
rect 211988 158714 212040 158720
rect 211896 158500 211948 158506
rect 211896 158442 211948 158448
rect 211804 155712 211856 155718
rect 211804 155654 211856 155660
rect 211712 155508 211764 155514
rect 211712 155450 211764 155456
rect 210424 150408 210476 150414
rect 210424 150350 210476 150356
rect 209884 16546 211016 16574
rect 210988 480 211016 16546
rect 212184 6914 212212 297463
rect 212264 297424 212316 297430
rect 212264 297366 212316 297372
rect 212092 6886 212212 6914
rect 212092 3330 212120 6886
rect 212276 3670 212304 297366
rect 212264 3664 212316 3670
rect 212264 3606 212316 3612
rect 212170 3496 212226 3505
rect 212170 3431 212226 3440
rect 212080 3324 212132 3330
rect 212080 3266 212132 3272
rect 212184 480 212212 3431
rect 212368 3262 212396 297735
rect 212460 3806 212488 303010
rect 213368 301504 213420 301510
rect 213368 301446 213420 301452
rect 213276 297560 213328 297566
rect 213276 297502 213328 297508
rect 213184 297492 213236 297498
rect 213184 297434 213236 297440
rect 213092 294976 213144 294982
rect 213092 294918 213144 294924
rect 213000 294772 213052 294778
rect 213000 294714 213052 294720
rect 213012 195294 213040 294714
rect 213000 195288 213052 195294
rect 213000 195230 213052 195236
rect 213104 159662 213132 294918
rect 213092 159656 213144 159662
rect 213092 159598 213144 159604
rect 213196 158914 213224 297434
rect 213288 158982 213316 297502
rect 213276 158976 213328 158982
rect 213276 158918 213328 158924
rect 213184 158908 213236 158914
rect 213184 158850 213236 158856
rect 213380 158846 213408 301446
rect 213472 159730 213500 303078
rect 213552 299940 213604 299946
rect 213552 299882 213604 299888
rect 213460 159724 213512 159730
rect 213460 159666 213512 159672
rect 213368 158840 213420 158846
rect 213368 158782 213420 158788
rect 213564 155786 213592 299882
rect 213736 297696 213788 297702
rect 213736 297638 213788 297644
rect 213644 297356 213696 297362
rect 213644 297298 213696 297304
rect 213552 155780 213604 155786
rect 213552 155722 213604 155728
rect 212448 3800 212500 3806
rect 212448 3742 212500 3748
rect 213366 3496 213422 3505
rect 213366 3431 213422 3440
rect 212356 3256 212408 3262
rect 212356 3198 212408 3204
rect 213380 480 213408 3431
rect 213656 3398 213684 297298
rect 213748 3874 213776 297638
rect 213840 4146 213868 305730
rect 214748 303544 214800 303550
rect 214748 303486 214800 303492
rect 214656 303272 214708 303278
rect 214656 303214 214708 303220
rect 214562 297936 214618 297945
rect 214562 297871 214618 297880
rect 214380 295044 214432 295050
rect 214380 294986 214432 294992
rect 214392 195566 214420 294986
rect 214472 294908 214524 294914
rect 214472 294850 214524 294856
rect 214380 195560 214432 195566
rect 214380 195502 214432 195508
rect 214484 159390 214512 294850
rect 214472 159384 214524 159390
rect 214472 159326 214524 159332
rect 214576 155650 214604 297871
rect 214668 158370 214696 303214
rect 214656 158364 214708 158370
rect 214656 158306 214708 158312
rect 214760 157894 214788 303486
rect 214840 303340 214892 303346
rect 214840 303282 214892 303288
rect 214852 158574 214880 303282
rect 214840 158568 214892 158574
rect 214840 158510 214892 158516
rect 214944 158302 214972 306002
rect 215024 303204 215076 303210
rect 215024 303146 215076 303152
rect 214932 158296 214984 158302
rect 214932 158238 214984 158244
rect 214748 157888 214800 157894
rect 214748 157830 214800 157836
rect 214564 155644 214616 155650
rect 214564 155586 214616 155592
rect 213828 4140 213880 4146
rect 213828 4082 213880 4088
rect 213736 3868 213788 3874
rect 213736 3810 213788 3816
rect 215036 3602 215064 303146
rect 215116 302796 215168 302802
rect 215116 302738 215168 302744
rect 215024 3596 215076 3602
rect 215024 3538 215076 3544
rect 214470 3496 214526 3505
rect 214470 3431 214526 3440
rect 213644 3392 213696 3398
rect 213644 3334 213696 3340
rect 214484 480 214512 3431
rect 215128 3233 215156 302738
rect 215220 3942 215248 307158
rect 218980 306332 219032 306338
rect 218980 306274 219032 306280
rect 218888 306264 218940 306270
rect 218888 306206 218940 306212
rect 216404 306128 216456 306134
rect 216404 306070 216456 306076
rect 216312 305924 216364 305930
rect 216312 305866 216364 305872
rect 216128 303612 216180 303618
rect 216128 303554 216180 303560
rect 216036 302864 216088 302870
rect 216036 302806 216088 302812
rect 215944 297288 215996 297294
rect 215944 297230 215996 297236
rect 215852 295112 215904 295118
rect 215852 295054 215904 295060
rect 215760 243568 215812 243574
rect 215760 243510 215812 243516
rect 215772 155242 215800 243510
rect 215864 189446 215892 295054
rect 215852 189440 215904 189446
rect 215852 189382 215904 189388
rect 215956 159526 215984 297230
rect 215944 159520 215996 159526
rect 215944 159462 215996 159468
rect 216048 157962 216076 302806
rect 216140 158642 216168 303554
rect 216220 303408 216272 303414
rect 216220 303350 216272 303356
rect 216128 158636 216180 158642
rect 216128 158578 216180 158584
rect 216232 158234 216260 303350
rect 216324 159798 216352 305866
rect 216312 159792 216364 159798
rect 216312 159734 216364 159740
rect 216220 158228 216272 158234
rect 216220 158170 216272 158176
rect 216416 158166 216444 306070
rect 216588 305856 216640 305862
rect 216588 305798 216640 305804
rect 216496 303476 216548 303482
rect 216496 303418 216548 303424
rect 216404 158160 216456 158166
rect 216404 158102 216456 158108
rect 216036 157956 216088 157962
rect 216036 157898 216088 157904
rect 215760 155236 215812 155242
rect 215760 155178 215812 155184
rect 215208 3936 215260 3942
rect 215208 3878 215260 3884
rect 215666 3496 215722 3505
rect 215666 3431 215722 3440
rect 215114 3224 215170 3233
rect 215114 3159 215170 3168
rect 215680 480 215708 3431
rect 216508 3369 216536 303418
rect 216600 4010 216628 305798
rect 217968 300008 218020 300014
rect 217968 299950 218020 299956
rect 217876 295180 217928 295186
rect 217876 295122 217928 295128
rect 217692 293412 217744 293418
rect 217692 293354 217744 293360
rect 217416 282396 217468 282402
rect 217416 282338 217468 282344
rect 217140 256352 217192 256358
rect 217140 256294 217192 256300
rect 217048 253632 217100 253638
rect 217048 253574 217100 253580
rect 216772 193180 216824 193186
rect 216772 193122 216824 193128
rect 216680 189032 216732 189038
rect 216680 188974 216732 188980
rect 216692 188193 216720 188974
rect 216678 188184 216734 188193
rect 216678 188119 216734 188128
rect 216784 180794 216812 193122
rect 217060 192817 217088 253574
rect 217152 196897 217180 256294
rect 217232 245200 217284 245206
rect 217232 245142 217284 245148
rect 217138 196888 217194 196897
rect 217138 196823 217194 196832
rect 217140 195560 217192 195566
rect 217140 195502 217192 195508
rect 217046 192808 217102 192817
rect 217046 192743 217102 192752
rect 216692 180766 216812 180794
rect 216692 16574 216720 180766
rect 217152 159594 217180 195502
rect 217244 168337 217272 245142
rect 217428 195945 217456 282338
rect 217600 260432 217652 260438
rect 217600 260374 217652 260380
rect 217508 243636 217560 243642
rect 217508 243578 217560 243584
rect 217414 195936 217470 195945
rect 217414 195871 217470 195880
rect 217324 195288 217376 195294
rect 217324 195230 217376 195236
rect 217230 168328 217286 168337
rect 217230 168263 217286 168272
rect 217140 159588 217192 159594
rect 217140 159530 217192 159536
rect 216692 16546 216904 16574
rect 216588 4004 216640 4010
rect 216588 3946 216640 3952
rect 216494 3360 216550 3369
rect 216494 3295 216550 3304
rect 216876 480 216904 16546
rect 217336 3534 217364 195230
rect 217520 155310 217548 243578
rect 217612 169969 217640 260374
rect 217704 193769 217732 293354
rect 217784 286476 217836 286482
rect 217784 286418 217836 286424
rect 217690 193760 217746 193769
rect 217690 193695 217746 193704
rect 217598 169960 217654 169969
rect 217598 169895 217654 169904
rect 217796 168065 217824 286418
rect 217782 168056 217838 168065
rect 217782 167991 217838 168000
rect 217888 159458 217916 295122
rect 217876 159452 217928 159458
rect 217876 159394 217928 159400
rect 217508 155304 217560 155310
rect 217508 155246 217560 155252
rect 217980 3738 218008 299950
rect 218796 297220 218848 297226
rect 218796 297162 218848 297168
rect 218428 283824 218480 283830
rect 218428 283766 218480 283772
rect 218440 243545 218468 283766
rect 218704 280968 218756 280974
rect 218704 280910 218756 280916
rect 218520 252204 218572 252210
rect 218520 252146 218572 252152
rect 218426 243536 218482 243545
rect 218426 243471 218482 243480
rect 218532 191049 218560 252146
rect 218612 243772 218664 243778
rect 218612 243714 218664 243720
rect 218518 191040 218574 191049
rect 218518 190975 218574 190984
rect 218520 189440 218572 189446
rect 218520 189382 218572 189388
rect 218532 155378 218560 189382
rect 218624 155446 218652 243714
rect 218716 189961 218744 280910
rect 218702 189952 218758 189961
rect 218702 189887 218758 189896
rect 218808 159866 218836 297162
rect 218796 159860 218848 159866
rect 218796 159802 218848 159808
rect 218900 158098 218928 306206
rect 218992 158438 219020 306274
rect 219072 305584 219124 305590
rect 219072 305526 219124 305532
rect 219084 158710 219112 305526
rect 219164 305516 219216 305522
rect 219164 305458 219216 305464
rect 219072 158704 219124 158710
rect 219072 158646 219124 158652
rect 218980 158432 219032 158438
rect 218980 158374 219032 158380
rect 218888 158092 218940 158098
rect 218888 158034 218940 158040
rect 219176 157826 219204 305458
rect 219348 301640 219400 301646
rect 219348 301582 219400 301588
rect 219256 243704 219308 243710
rect 219256 243646 219308 243652
rect 219164 157820 219216 157826
rect 219164 157762 219216 157768
rect 218612 155440 218664 155446
rect 218612 155382 218664 155388
rect 218520 155372 218572 155378
rect 218520 155314 218572 155320
rect 219268 6914 219296 243646
rect 219176 6886 219296 6914
rect 217968 3732 218020 3738
rect 217968 3674 218020 3680
rect 218058 3632 218114 3641
rect 218058 3567 218114 3576
rect 217324 3528 217376 3534
rect 217324 3470 217376 3476
rect 218072 480 218100 3567
rect 219176 3466 219204 6886
rect 219360 4078 219388 301582
rect 225616 267714 225644 435134
rect 229744 433696 229796 433702
rect 229744 433638 229796 433644
rect 229756 411262 229784 433638
rect 231124 433628 231176 433634
rect 231124 433570 231176 433576
rect 229744 411256 229796 411262
rect 229744 411198 229796 411204
rect 231136 376038 231164 433570
rect 231228 398818 231256 436630
rect 244832 436416 244884 436422
rect 244832 436358 244884 436364
rect 244188 436348 244240 436354
rect 244188 436290 244240 436296
rect 237470 436248 237526 436257
rect 237470 436183 237526 436192
rect 235722 436112 235778 436121
rect 235722 436047 235778 436056
rect 234434 434752 234490 434761
rect 234434 434687 234490 434696
rect 233882 433800 233938 433809
rect 233882 433735 233938 433744
rect 232686 433392 232742 433401
rect 232686 433327 232742 433336
rect 232700 432276 232728 433327
rect 233896 432276 233924 433735
rect 234448 432276 234476 434687
rect 235736 432276 235764 436047
rect 236274 434888 236330 434897
rect 236274 434823 236330 434832
rect 236288 432276 236316 434823
rect 237484 432276 237512 436183
rect 241152 434784 241204 434790
rect 241152 434726 241204 434732
rect 238760 434104 238812 434110
rect 238760 434046 238812 434052
rect 238114 433528 238170 433537
rect 238114 433463 238170 433472
rect 238128 432276 238156 433463
rect 238772 432276 238800 434046
rect 240508 433900 240560 433906
rect 240508 433842 240560 433848
rect 239310 433664 239366 433673
rect 239310 433599 239366 433608
rect 239324 432276 239352 433599
rect 240046 432304 240102 432313
rect 239982 432262 240046 432290
rect 240520 432276 240548 433842
rect 241164 432276 241192 434726
rect 243544 434512 243596 434518
rect 243544 434454 243596 434460
rect 242348 433764 242400 433770
rect 242348 433706 242400 433712
rect 242360 432276 242388 433706
rect 243556 432276 243584 434454
rect 244200 432276 244228 436290
rect 244844 432276 244872 436358
rect 246028 435056 246080 435062
rect 246028 434998 246080 435004
rect 246040 432276 246068 434998
rect 246672 434172 246724 434178
rect 246672 434114 246724 434120
rect 246684 432276 246712 434114
rect 248420 433832 248472 433838
rect 248420 433774 248472 433780
rect 247868 433424 247920 433430
rect 247868 433366 247920 433372
rect 247880 432276 247908 433366
rect 248432 432276 248460 433774
rect 249708 433356 249760 433362
rect 249708 433298 249760 433304
rect 249090 432274 249472 432290
rect 249720 432276 249748 433298
rect 250548 432290 250576 441586
rect 251192 432290 251220 464306
rect 251836 432546 251864 470562
rect 252480 454850 252508 476167
rect 252560 467152 252612 467158
rect 252560 467094 252612 467100
rect 252468 454844 252520 454850
rect 252468 454786 252520 454792
rect 252572 441614 252600 467094
rect 253768 450770 253796 476167
rect 255240 474094 255268 476167
rect 255228 474088 255280 474094
rect 255228 474030 255280 474036
rect 255320 472660 255372 472666
rect 255320 472602 255372 472608
rect 253940 458856 253992 458862
rect 253940 458798 253992 458804
rect 253756 450764 253808 450770
rect 253756 450706 253808 450712
rect 252572 441586 252968 441614
rect 252744 440904 252796 440910
rect 252744 440846 252796 440852
rect 251824 432540 251876 432546
rect 251824 432482 251876 432488
rect 251836 432290 251864 432482
rect 249090 432268 249484 432274
rect 249090 432262 249432 432268
rect 240046 432239 240102 432248
rect 250548 432262 250930 432290
rect 251192 432262 251482 432290
rect 251836 432262 252126 432290
rect 252756 432276 252784 440846
rect 252940 432290 252968 441586
rect 253202 433936 253258 433945
rect 253202 433871 253258 433880
rect 253216 432614 253244 433871
rect 253204 432608 253256 432614
rect 253204 432550 253256 432556
rect 252940 432262 253322 432290
rect 253952 432276 253980 458798
rect 254032 453348 254084 453354
rect 254032 453290 254084 453296
rect 254044 436830 254072 453290
rect 254124 442264 254176 442270
rect 254124 442206 254176 442212
rect 254032 436824 254084 436830
rect 254032 436766 254084 436772
rect 254136 432290 254164 442206
rect 254860 436824 254912 436830
rect 254860 436766 254912 436772
rect 254872 432290 254900 436766
rect 255332 432290 255360 472602
rect 256528 461854 256556 476167
rect 256516 461848 256568 461854
rect 256516 461790 256568 461796
rect 256620 447982 256648 476303
rect 257986 476232 258042 476241
rect 257986 476167 258042 476176
rect 256700 460284 256752 460290
rect 256700 460226 256752 460232
rect 256608 447976 256660 447982
rect 256608 447918 256660 447924
rect 255412 443692 255464 443698
rect 255412 443634 255464 443640
rect 255424 441614 255452 443634
rect 255424 441586 255912 441614
rect 255884 432290 255912 441586
rect 256712 436830 256740 460226
rect 256792 454776 256844 454782
rect 256792 454718 256844 454724
rect 256700 436824 256752 436830
rect 256700 436766 256752 436772
rect 256804 432290 256832 454718
rect 258000 445126 258028 476167
rect 259288 463010 259316 476575
rect 264940 476575 264942 476584
rect 264888 476546 264940 476552
rect 259366 476504 259422 476513
rect 259366 476439 259368 476448
rect 259420 476439 259422 476448
rect 259368 476410 259420 476416
rect 260654 476368 260710 476377
rect 260654 476303 260710 476312
rect 262034 476368 262090 476377
rect 262034 476303 262090 476312
rect 259460 465724 259512 465730
rect 259460 465666 259512 465672
rect 259276 463004 259328 463010
rect 259276 462946 259328 462952
rect 258080 461644 258132 461650
rect 258080 461586 258132 461592
rect 257988 445120 258040 445126
rect 257988 445062 258040 445068
rect 258092 436830 258120 461586
rect 258172 449200 258224 449206
rect 258172 449142 258224 449148
rect 258184 436898 258212 449142
rect 258264 445052 258316 445058
rect 258264 444994 258316 445000
rect 258276 441614 258304 444994
rect 258276 441586 258396 441614
rect 258172 436892 258224 436898
rect 258172 436834 258224 436840
rect 257252 436824 257304 436830
rect 257252 436766 257304 436772
rect 258080 436824 258132 436830
rect 258080 436766 258132 436772
rect 257264 432290 257292 436766
rect 258368 432290 258396 441586
rect 258540 436892 258592 436898
rect 258540 436834 258592 436840
rect 254136 432262 254518 432290
rect 254872 432262 255162 432290
rect 255332 432262 255806 432290
rect 255884 432262 256358 432290
rect 256804 432262 257002 432290
rect 257264 432262 257554 432290
rect 258198 432262 258396 432290
rect 258552 432290 258580 436834
rect 259472 436830 259500 465666
rect 260668 457570 260696 476303
rect 260746 476232 260802 476241
rect 260746 476167 260802 476176
rect 260656 457564 260708 457570
rect 260656 457506 260708 457512
rect 260760 446554 260788 476167
rect 262048 459066 262076 476303
rect 262126 476232 262182 476241
rect 262126 476167 262182 476176
rect 263506 476232 263562 476241
rect 263506 476167 263562 476176
rect 264794 476232 264850 476241
rect 264794 476167 264850 476176
rect 262036 459060 262088 459066
rect 262036 459002 262088 459008
rect 260840 447840 260892 447846
rect 260840 447782 260892 447788
rect 260748 446548 260800 446554
rect 260748 446490 260800 446496
rect 259552 446480 259604 446486
rect 259552 446422 259604 446428
rect 259092 436824 259144 436830
rect 259092 436766 259144 436772
rect 259460 436824 259512 436830
rect 259460 436766 259512 436772
rect 259104 432290 259132 436766
rect 259564 432290 259592 446422
rect 260852 441614 260880 447782
rect 260852 441586 261432 441614
rect 260380 436824 260432 436830
rect 260380 436766 260432 436772
rect 260392 432290 260420 436766
rect 261208 435736 261260 435742
rect 261208 435678 261260 435684
rect 258552 432262 258842 432290
rect 259104 432262 259394 432290
rect 259564 432262 260038 432290
rect 260392 432262 260682 432290
rect 261220 432276 261248 435678
rect 261404 432290 261432 441586
rect 262140 438258 262168 476167
rect 262220 456136 262272 456142
rect 262220 456078 262272 456084
rect 262128 438252 262180 438258
rect 262128 438194 262180 438200
rect 262232 432290 262260 456078
rect 263520 439686 263548 476167
rect 263600 468512 263652 468518
rect 263600 468454 263652 468460
rect 263508 439680 263560 439686
rect 263508 439622 263560 439628
rect 263048 435804 263100 435810
rect 263048 435746 263100 435752
rect 262680 433424 262732 433430
rect 262680 433366 262732 433372
rect 262692 432614 262720 433366
rect 262680 432608 262732 432614
rect 262680 432550 262732 432556
rect 261404 432262 261878 432290
rect 262232 432262 262430 432290
rect 263060 432276 263088 435746
rect 263612 434586 263640 468454
rect 263692 450628 263744 450634
rect 263692 450570 263744 450576
rect 263600 434580 263652 434586
rect 263600 434522 263652 434528
rect 263704 432276 263732 450570
rect 264808 439754 264836 476167
rect 264796 439748 264848 439754
rect 264796 439690 264848 439696
rect 264888 437096 264940 437102
rect 264888 437038 264940 437044
rect 263784 436756 263836 436762
rect 263784 436698 263836 436704
rect 263796 435742 263824 436698
rect 263784 435736 263836 435742
rect 263784 435678 263836 435684
rect 263876 434580 263928 434586
rect 263876 434522 263928 434528
rect 263888 432290 263916 434522
rect 263888 432262 264270 432290
rect 264900 432276 264928 437038
rect 264992 434586 265020 478178
rect 266266 476368 266322 476377
rect 266266 476303 266322 476312
rect 266174 476232 266230 476241
rect 266174 476167 266230 476176
rect 266188 465934 266216 476167
rect 266176 465928 266228 465934
rect 266176 465870 266228 465876
rect 265072 451988 265124 451994
rect 265072 451930 265124 451936
rect 264980 434580 265032 434586
rect 264980 434522 265032 434528
rect 265084 432290 265112 451930
rect 266280 439822 266308 476303
rect 266268 439816 266320 439822
rect 266268 439758 266320 439764
rect 265716 434580 265768 434586
rect 265716 434522 265768 434528
rect 265728 432290 265756 434522
rect 266372 432290 266400 478314
rect 266464 441614 266492 478518
rect 267740 478508 267792 478514
rect 267740 478450 267792 478456
rect 267554 476368 267610 476377
rect 267554 476303 267610 476312
rect 267568 464506 267596 476303
rect 267646 476232 267702 476241
rect 267646 476167 267702 476176
rect 267556 464500 267608 464506
rect 267556 464442 267608 464448
rect 266464 441586 266952 441614
rect 266924 432290 266952 441586
rect 267660 439550 267688 476167
rect 267752 441614 267780 478450
rect 302240 478440 302292 478446
rect 302240 478382 302292 478388
rect 281540 478168 281592 478174
rect 281540 478110 281592 478116
rect 269026 477320 269082 477329
rect 269026 477255 269082 477264
rect 269040 476542 269068 477255
rect 281446 476912 281502 476921
rect 281446 476847 281502 476856
rect 269028 476536 269080 476542
rect 269028 476478 269080 476484
rect 274546 476504 274602 476513
rect 274546 476439 274602 476448
rect 271694 476368 271750 476377
rect 271694 476303 271750 476312
rect 274454 476368 274510 476377
rect 274454 476303 274510 476312
rect 268934 476232 268990 476241
rect 268934 476167 268990 476176
rect 270406 476232 270462 476241
rect 270406 476167 270462 476176
rect 267752 441586 268056 441614
rect 267648 439544 267700 439550
rect 267648 439486 267700 439492
rect 267924 436960 267976 436966
rect 267924 436902 267976 436908
rect 265084 432262 265466 432290
rect 265728 432262 266110 432290
rect 266372 432262 266754 432290
rect 266924 432262 267306 432290
rect 267936 432276 267964 436902
rect 268028 432290 268056 441586
rect 268948 439618 268976 476167
rect 269304 468648 269356 468654
rect 269304 468590 269356 468596
rect 269212 443828 269264 443834
rect 269212 443770 269264 443776
rect 268936 439612 268988 439618
rect 268936 439554 268988 439560
rect 269224 437474 269252 443770
rect 269316 441614 269344 468590
rect 270420 467294 270448 476167
rect 271708 468654 271736 476303
rect 271786 476232 271842 476241
rect 271786 476167 271842 476176
rect 273166 476232 273222 476241
rect 273166 476167 273222 476176
rect 274362 476232 274418 476241
rect 274362 476167 274418 476176
rect 271696 468648 271748 468654
rect 271696 468590 271748 468596
rect 270408 467288 270460 467294
rect 270408 467230 270460 467236
rect 271800 453422 271828 476167
rect 273180 458998 273208 476167
rect 273260 465792 273312 465798
rect 273260 465734 273312 465740
rect 273168 458992 273220 458998
rect 273168 458934 273220 458940
rect 271880 457496 271932 457502
rect 271880 457438 271932 457444
rect 270500 453416 270552 453422
rect 270500 453358 270552 453364
rect 271788 453416 271840 453422
rect 271788 453358 271840 453364
rect 269316 441586 269896 441614
rect 269224 437446 269344 437474
rect 268568 436824 268620 436830
rect 268568 436766 268620 436772
rect 268580 435810 268608 436766
rect 268568 435804 268620 435810
rect 268568 435746 268620 435752
rect 269120 434036 269172 434042
rect 269120 433978 269172 433984
rect 268028 432262 268502 432290
rect 269132 432276 269160 433978
rect 269316 432290 269344 437446
rect 269396 433968 269448 433974
rect 269396 433910 269448 433916
rect 269408 432750 269436 433910
rect 269396 432744 269448 432750
rect 269396 432686 269448 432692
rect 269868 432290 269896 441586
rect 270512 437474 270540 453358
rect 270592 446412 270644 446418
rect 270592 446354 270644 446360
rect 270604 441614 270632 446354
rect 270604 441586 271184 441614
rect 270512 437446 270632 437474
rect 270604 432290 270632 437446
rect 271156 432290 271184 441586
rect 271892 432290 271920 457438
rect 271972 445188 272024 445194
rect 271972 445130 272024 445136
rect 271984 441614 272012 445130
rect 271984 441586 272472 441614
rect 272248 433356 272300 433362
rect 272248 433298 272300 433304
rect 269316 432262 269790 432290
rect 269868 432262 270342 432290
rect 270604 432262 270986 432290
rect 271156 432262 271538 432290
rect 271892 432262 272182 432290
rect 249432 432210 249484 432216
rect 247592 432200 247644 432206
rect 237286 432168 237342 432177
rect 236946 432126 237286 432154
rect 241822 432138 242112 432154
rect 247250 432148 247592 432154
rect 247250 432142 247644 432148
rect 241822 432132 242124 432138
rect 241822 432126 242072 432132
rect 237286 432103 237342 432112
rect 247250 432126 247632 432142
rect 242072 432074 242124 432080
rect 245568 432064 245620 432070
rect 235446 432032 235502 432041
rect 233266 432002 233648 432018
rect 233266 431996 233660 432002
rect 233266 431990 233608 431996
rect 235106 431990 235446 432018
rect 245410 432012 245568 432018
rect 245410 432006 245620 432012
rect 245410 431990 245608 432006
rect 235446 431967 235502 431976
rect 233608 431938 233660 431944
rect 272260 431934 272288 433298
rect 272444 432290 272472 441586
rect 273272 436966 273300 465734
rect 273352 447908 273404 447914
rect 273352 447850 273404 447856
rect 273364 441614 273392 447850
rect 273364 441586 273484 441614
rect 273260 436960 273312 436966
rect 273260 436902 273312 436908
rect 273456 432290 273484 441586
rect 274376 438190 274404 476167
rect 274468 470014 274496 476303
rect 274560 474230 274588 476439
rect 277306 476368 277362 476377
rect 277306 476303 277362 476312
rect 278594 476368 278650 476377
rect 278594 476303 278650 476312
rect 275926 476232 275982 476241
rect 275926 476167 275982 476176
rect 277214 476232 277270 476241
rect 277214 476167 277270 476176
rect 274548 474224 274600 474230
rect 274548 474166 274600 474172
rect 274456 470008 274508 470014
rect 274456 469950 274508 469956
rect 274640 469872 274692 469878
rect 274640 469814 274692 469820
rect 274364 438184 274416 438190
rect 274364 438126 274416 438132
rect 274652 436966 274680 469814
rect 275940 454714 275968 476167
rect 277228 460358 277256 476167
rect 277216 460352 277268 460358
rect 277216 460294 277268 460300
rect 276020 456068 276072 456074
rect 276020 456010 276072 456016
rect 274732 454708 274784 454714
rect 274732 454650 274784 454656
rect 275928 454708 275980 454714
rect 275928 454650 275980 454656
rect 273628 436960 273680 436966
rect 273628 436902 273680 436908
rect 274640 436960 274692 436966
rect 274640 436902 274692 436908
rect 272444 432262 272826 432290
rect 273378 432262 273484 432290
rect 273640 432290 273668 436902
rect 274744 432290 274772 454650
rect 274824 450560 274876 450566
rect 274824 450502 274876 450508
rect 273640 432262 274022 432290
rect 274666 432262 274772 432290
rect 274836 432290 274864 450502
rect 275468 436960 275520 436966
rect 275468 436902 275520 436908
rect 275480 432290 275508 436902
rect 276032 432290 276060 456010
rect 277320 442474 277348 476303
rect 277400 464432 277452 464438
rect 277400 464374 277452 464380
rect 277308 442468 277360 442474
rect 277308 442410 277360 442416
rect 277032 440972 277084 440978
rect 277032 440914 277084 440920
rect 274836 432262 275218 432290
rect 275480 432262 275862 432290
rect 276032 432262 276414 432290
rect 277044 432276 277072 440914
rect 277412 432290 277440 464374
rect 278608 461786 278636 476303
rect 278686 476232 278742 476241
rect 278686 476167 278742 476176
rect 280066 476232 280122 476241
rect 280066 476167 280122 476176
rect 278596 461780 278648 461786
rect 278596 461722 278648 461728
rect 277492 458924 277544 458930
rect 277492 458866 277544 458872
rect 277504 441614 277532 458866
rect 278700 443834 278728 476167
rect 278780 460216 278832 460222
rect 278780 460158 278832 460164
rect 278688 443828 278740 443834
rect 278688 443770 278740 443776
rect 277504 441586 277808 441614
rect 277780 432290 277808 441586
rect 278792 436966 278820 460158
rect 280080 456074 280108 476167
rect 281460 475522 281488 476847
rect 281448 475516 281500 475522
rect 281448 475458 281500 475464
rect 280160 474020 280212 474026
rect 280160 473962 280212 473968
rect 280068 456068 280120 456074
rect 280068 456010 280120 456016
rect 278872 451920 278924 451926
rect 278872 451862 278924 451868
rect 278780 436960 278832 436966
rect 278780 436902 278832 436908
rect 277412 432262 277702 432290
rect 277780 432262 278254 432290
rect 278884 432276 278912 451862
rect 278964 442332 279016 442338
rect 278964 442274 279016 442280
rect 278976 441614 279004 442274
rect 278976 441586 279096 441614
rect 279068 432290 279096 441586
rect 279700 436960 279752 436966
rect 279700 436902 279752 436908
rect 279712 432290 279740 436902
rect 279976 434036 280028 434042
rect 279976 433978 280028 433984
rect 279988 432750 280016 433978
rect 280068 433356 280120 433362
rect 280068 433298 280120 433304
rect 279976 432744 280028 432750
rect 279976 432686 280028 432692
rect 280080 432682 280108 433298
rect 280068 432676 280120 432682
rect 280068 432618 280120 432624
rect 280172 432426 280200 473962
rect 280252 467220 280304 467226
rect 280252 467162 280304 467168
rect 280264 441614 280292 467162
rect 280264 441586 280936 441614
rect 280172 432398 280384 432426
rect 280356 432290 280384 432398
rect 280908 432290 280936 441586
rect 281552 436966 281580 478110
rect 284206 476232 284262 476241
rect 284206 476167 284262 476176
rect 286966 476232 287022 476241
rect 286966 476167 287022 476176
rect 288346 476232 288402 476241
rect 288346 476167 288402 476176
rect 291106 476232 291162 476241
rect 291106 476167 291162 476176
rect 293866 476232 293922 476241
rect 293866 476167 293922 476176
rect 296626 476232 296682 476241
rect 296626 476167 296682 476176
rect 299386 476232 299442 476241
rect 299386 476167 299442 476176
rect 302146 476232 302202 476241
rect 302146 476167 302202 476176
rect 282920 474768 282972 474774
rect 282920 474710 282972 474716
rect 281632 461712 281684 461718
rect 281632 461654 281684 461660
rect 281540 436960 281592 436966
rect 281540 436902 281592 436908
rect 281644 432290 281672 461654
rect 282932 436966 282960 474710
rect 284220 471306 284248 476167
rect 283012 471300 283064 471306
rect 283012 471242 283064 471248
rect 284208 471300 284260 471306
rect 284208 471242 284260 471248
rect 282092 436960 282144 436966
rect 282092 436902 282144 436908
rect 282920 436960 282972 436966
rect 282920 436902 282972 436908
rect 282104 432290 282132 436902
rect 282184 434852 282236 434858
rect 282184 434794 282236 434800
rect 282196 434110 282224 434794
rect 282184 434104 282236 434110
rect 282184 434046 282236 434052
rect 282920 433764 282972 433770
rect 282920 433706 282972 433712
rect 282932 432750 282960 433706
rect 282920 432744 282972 432750
rect 282920 432686 282972 432692
rect 283024 432290 283052 471242
rect 284484 462392 284536 462398
rect 284484 462334 284536 462340
rect 284392 448588 284444 448594
rect 284392 448530 284444 448536
rect 283380 436960 283432 436966
rect 283380 436902 283432 436908
rect 283392 432290 283420 436902
rect 284404 432290 284432 448530
rect 284496 441614 284524 462334
rect 284496 441586 284616 441614
rect 279068 432262 279450 432290
rect 279712 432262 280094 432290
rect 280356 432262 280738 432290
rect 280908 432262 281290 432290
rect 281644 432262 281934 432290
rect 282104 432262 282486 432290
rect 283024 432262 283130 432290
rect 283392 432262 283774 432290
rect 284326 432262 284432 432290
rect 284588 432290 284616 441586
rect 286980 440978 287008 476167
rect 288360 451926 288388 476167
rect 291120 468654 291148 476167
rect 289084 468648 289136 468654
rect 289084 468590 289136 468596
rect 291108 468648 291160 468654
rect 291108 468590 291160 468596
rect 288348 451920 288400 451926
rect 288348 451862 288400 451868
rect 286968 440972 287020 440978
rect 286968 440914 287020 440920
rect 286140 436688 286192 436694
rect 286140 436630 286192 436636
rect 285496 434920 285548 434926
rect 285496 434862 285548 434868
rect 285680 434920 285732 434926
rect 285680 434862 285732 434868
rect 284588 432262 284970 432290
rect 285508 432276 285536 434862
rect 285692 434178 285720 434862
rect 285680 434172 285732 434178
rect 285680 434114 285732 434120
rect 286152 432276 286180 436630
rect 287336 434988 287388 434994
rect 287336 434930 287388 434936
rect 286784 433696 286836 433702
rect 286784 433638 286836 433644
rect 286796 432276 286824 433638
rect 287348 432276 287376 434930
rect 289096 434042 289124 468590
rect 293880 449342 293908 476167
rect 293868 449336 293920 449342
rect 293868 449278 293920 449284
rect 296640 447914 296668 476167
rect 299400 469878 299428 476167
rect 302160 475590 302188 476167
rect 302148 475584 302200 475590
rect 302148 475526 302200 475532
rect 300860 471368 300912 471374
rect 300860 471310 300912 471316
rect 299388 469872 299440 469878
rect 299388 469814 299440 469820
rect 297364 465928 297416 465934
rect 297364 465870 297416 465876
rect 296628 447908 296680 447914
rect 296628 447850 296680 447856
rect 295892 436620 295944 436626
rect 295892 436562 295944 436568
rect 295248 436552 295300 436558
rect 295248 436494 295300 436500
rect 291660 436212 291712 436218
rect 291660 436154 291712 436160
rect 289176 435260 289228 435266
rect 289176 435202 289228 435208
rect 289084 434036 289136 434042
rect 289084 433978 289136 433984
rect 287980 433968 288032 433974
rect 287980 433910 288032 433916
rect 287992 432276 288020 433910
rect 288624 433628 288676 433634
rect 288624 433570 288676 433576
rect 288636 432276 288664 433570
rect 289188 432276 289216 435202
rect 291016 435192 291068 435198
rect 291016 435134 291068 435140
rect 290372 434240 290424 434246
rect 290372 434182 290424 434188
rect 289728 433832 289780 433838
rect 289728 433774 289780 433780
rect 289740 432818 289768 433774
rect 289820 433356 289872 433362
rect 289820 433298 289872 433304
rect 289728 432812 289780 432818
rect 289728 432754 289780 432760
rect 289832 432276 289860 433298
rect 290384 432276 290412 434182
rect 291028 432276 291056 435134
rect 291672 432276 291700 436154
rect 292212 436144 292264 436150
rect 292212 436086 292264 436092
rect 292224 432276 292252 436086
rect 294694 435296 294750 435305
rect 294694 435231 294750 435240
rect 292856 433560 292908 433566
rect 292856 433502 292908 433508
rect 292868 432276 292896 433502
rect 294052 433492 294104 433498
rect 294052 433434 294104 433440
rect 293408 432472 293460 432478
rect 293408 432414 293460 432420
rect 293420 432276 293448 432414
rect 294064 432276 294092 433434
rect 294708 432276 294736 435231
rect 295260 432276 295288 436494
rect 295904 432276 295932 436562
rect 296442 435024 296498 435033
rect 296442 434959 296498 434968
rect 296456 432276 296484 434959
rect 297376 434110 297404 465870
rect 298744 459060 298796 459066
rect 298744 459002 298796 459008
rect 297732 436484 297784 436490
rect 297732 436426 297784 436432
rect 297364 434104 297416 434110
rect 297364 434046 297416 434052
rect 297088 432404 297140 432410
rect 297088 432346 297140 432352
rect 297100 432276 297128 432346
rect 297744 432276 297772 436426
rect 298284 435124 298336 435130
rect 298284 435066 298336 435072
rect 298296 432276 298324 435066
rect 298756 434178 298784 459002
rect 300872 441614 300900 471310
rect 300872 441586 301544 441614
rect 300768 436280 300820 436286
rect 300768 436222 300820 436228
rect 300122 435160 300178 435169
rect 300122 435095 300178 435104
rect 298744 434172 298796 434178
rect 298744 434114 298796 434120
rect 298926 433936 298982 433945
rect 298926 433871 298982 433880
rect 298940 432276 298968 433871
rect 300136 432276 300164 435095
rect 300780 432276 300808 436222
rect 301044 432336 301096 432342
rect 301516 432290 301544 441586
rect 302252 434586 302280 478382
rect 357452 478378 357480 700334
rect 358820 700324 358872 700330
rect 358820 700266 358872 700272
rect 357440 478372 357492 478378
rect 357440 478314 357492 478320
rect 310520 478304 310572 478310
rect 310520 478246 310572 478252
rect 306102 477048 306158 477057
rect 306102 476983 306158 476992
rect 306116 476678 306144 476983
rect 309140 476808 309192 476814
rect 309046 476776 309102 476785
rect 309140 476750 309192 476756
rect 309046 476711 309102 476720
rect 305000 476672 305052 476678
rect 305000 476614 305052 476620
rect 306104 476672 306156 476678
rect 306104 476614 306156 476620
rect 303526 476368 303582 476377
rect 303526 476303 303528 476312
rect 303580 476303 303582 476312
rect 303528 476274 303580 476280
rect 303620 474156 303672 474162
rect 303620 474098 303672 474104
rect 302332 450696 302384 450702
rect 302332 450638 302384 450644
rect 302240 434580 302292 434586
rect 302240 434522 302292 434528
rect 302344 432290 302372 450638
rect 302884 434580 302936 434586
rect 302884 434522 302936 434528
rect 302896 432290 302924 434522
rect 303632 432290 303660 474098
rect 304356 438320 304408 438326
rect 304356 438262 304408 438268
rect 301096 432284 301346 432290
rect 301044 432278 301346 432284
rect 301056 432262 301346 432278
rect 301516 432262 301990 432290
rect 302344 432262 302634 432290
rect 302896 432262 303186 432290
rect 303632 432262 303830 432290
rect 304368 432276 304396 438262
rect 304908 433356 304960 433362
rect 304908 433298 304960 433304
rect 304920 432290 304948 433298
rect 305012 432698 305040 476614
rect 309060 476270 309088 476711
rect 309048 476264 309100 476270
rect 309048 476206 309100 476212
rect 307760 476196 307812 476202
rect 307760 476138 307812 476144
rect 305092 475448 305144 475454
rect 305092 475390 305144 475396
rect 305104 434586 305132 475390
rect 306380 460420 306432 460426
rect 306380 460362 306432 460368
rect 305184 453484 305236 453490
rect 305184 453426 305236 453432
rect 305092 434580 305144 434586
rect 305092 434522 305144 434528
rect 305196 433362 305224 453426
rect 306392 441614 306420 460362
rect 306392 441586 307064 441614
rect 306840 439884 306892 439890
rect 306840 439826 306892 439832
rect 305828 434580 305880 434586
rect 305828 434522 305880 434528
rect 305184 433356 305236 433362
rect 305184 433298 305236 433304
rect 305012 432670 305224 432698
rect 305196 432290 305224 432670
rect 305840 432290 305868 434522
rect 304920 432262 305026 432290
rect 305196 432262 305670 432290
rect 305840 432262 306222 432290
rect 306852 432276 306880 439826
rect 307036 432290 307064 441586
rect 307772 432290 307800 476138
rect 307852 472728 307904 472734
rect 307852 472670 307904 472676
rect 307864 441614 307892 472670
rect 307864 441586 308352 441614
rect 308324 432290 308352 441586
rect 309152 434654 309180 476750
rect 309232 476400 309284 476406
rect 309232 476342 309284 476348
rect 309140 434648 309192 434654
rect 309140 434590 309192 434596
rect 309244 434586 309272 476342
rect 309324 452056 309376 452062
rect 309324 451998 309376 452004
rect 309232 434580 309284 434586
rect 309232 434522 309284 434528
rect 309336 432290 309364 451998
rect 310532 437474 310560 478246
rect 358832 478242 358860 700266
rect 360844 670744 360896 670750
rect 360844 670686 360896 670692
rect 359464 563100 359516 563106
rect 359464 563042 359516 563048
rect 358820 478236 358872 478242
rect 358820 478178 358872 478184
rect 321466 477048 321522 477057
rect 321466 476983 321522 476992
rect 311900 476740 311952 476746
rect 311900 476682 311952 476688
rect 311806 476232 311862 476241
rect 311806 476167 311862 476176
rect 311820 476134 311848 476167
rect 311808 476128 311860 476134
rect 311808 476070 311860 476076
rect 310612 449268 310664 449274
rect 310612 449210 310664 449216
rect 310624 441614 310652 449210
rect 310624 441586 311296 441614
rect 310532 437446 310744 437474
rect 310060 434648 310112 434654
rect 310060 434590 310112 434596
rect 309508 434580 309560 434586
rect 309508 434522 309560 434528
rect 307036 432262 307418 432290
rect 307772 432262 308062 432290
rect 308324 432262 308706 432290
rect 309258 432262 309364 432290
rect 309520 432290 309548 434522
rect 310072 432290 310100 434590
rect 310716 432290 310744 437446
rect 311268 432290 311296 441586
rect 311912 436966 311940 476682
rect 314566 476640 314622 476649
rect 314566 476575 314622 476584
rect 317420 476604 317472 476610
rect 314580 474026 314608 476575
rect 317420 476546 317472 476552
rect 314660 476468 314712 476474
rect 314660 476410 314712 476416
rect 314568 474020 314620 474026
rect 314568 473962 314620 473968
rect 313280 469940 313332 469946
rect 313280 469882 313332 469888
rect 311992 461848 312044 461854
rect 311992 461790 312044 461796
rect 311900 436960 311952 436966
rect 311900 436902 311952 436908
rect 312004 432290 312032 461790
rect 312636 436960 312688 436966
rect 312636 436902 312688 436908
rect 312648 432290 312676 436902
rect 313292 432290 313320 469882
rect 314108 441040 314160 441046
rect 314108 440982 314160 440988
rect 309520 432262 309902 432290
rect 310072 432262 310454 432290
rect 310716 432262 311098 432290
rect 311268 432262 311742 432290
rect 312004 432262 312294 432290
rect 312648 432262 312938 432290
rect 313292 432262 313582 432290
rect 314120 432276 314148 440982
rect 314672 432290 314700 476410
rect 315946 476232 316002 476241
rect 315946 476167 316002 476176
rect 315960 472734 315988 476167
rect 316132 475380 316184 475386
rect 316132 475322 316184 475328
rect 315948 472728 316000 472734
rect 315948 472670 316000 472676
rect 314752 443760 314804 443766
rect 314752 443702 314804 443708
rect 314764 432698 314792 443702
rect 314844 442400 314896 442406
rect 314844 442342 314896 442348
rect 314856 441614 314884 442342
rect 316144 441614 316172 475322
rect 314856 441586 315528 441614
rect 316144 441586 316816 441614
rect 314764 432670 314976 432698
rect 314948 432290 314976 432670
rect 315500 432290 315528 441586
rect 316592 434172 316644 434178
rect 316592 434114 316644 434120
rect 314672 432262 314778 432290
rect 314948 432262 315330 432290
rect 315500 432262 315974 432290
rect 316604 432276 316632 434114
rect 316788 432290 316816 441586
rect 317432 436966 317460 476546
rect 318706 476504 318762 476513
rect 318706 476439 318762 476448
rect 318720 476406 318748 476439
rect 318708 476400 318760 476406
rect 318708 476342 318760 476348
rect 321480 476338 321508 476983
rect 322204 476672 322256 476678
rect 322204 476614 322256 476620
rect 321560 476536 321612 476542
rect 321560 476478 321612 476484
rect 320824 476332 320876 476338
rect 320824 476274 320876 476280
rect 321468 476332 321520 476338
rect 321468 476274 321520 476280
rect 318800 472796 318852 472802
rect 318800 472738 318852 472744
rect 317512 456204 317564 456210
rect 317512 456146 317564 456152
rect 317420 436960 317472 436966
rect 317420 436902 317472 436908
rect 317524 432290 317552 456146
rect 318812 436966 318840 472738
rect 318892 468580 318944 468586
rect 318892 468522 318944 468528
rect 317972 436960 318024 436966
rect 317972 436902 318024 436908
rect 318800 436960 318852 436966
rect 318800 436902 318852 436908
rect 317984 432290 318012 436902
rect 318904 432290 318932 468522
rect 320364 465860 320416 465866
rect 320364 465802 320416 465808
rect 320272 454844 320324 454850
rect 320272 454786 320324 454792
rect 320284 436966 320312 454786
rect 320376 441614 320404 465802
rect 320376 441586 320496 441614
rect 319260 436960 319312 436966
rect 319260 436902 319312 436908
rect 320272 436960 320324 436966
rect 320272 436902 320324 436908
rect 319272 432290 319300 436902
rect 320180 434104 320232 434110
rect 320180 434046 320232 434052
rect 316788 432262 317170 432290
rect 317524 432262 317814 432290
rect 317984 432262 318366 432290
rect 318904 432262 319010 432290
rect 319272 432262 319654 432290
rect 320192 432276 320220 434046
rect 320468 432290 320496 441586
rect 320836 434110 320864 476274
rect 321100 436960 321152 436966
rect 321100 436902 321152 436908
rect 320824 434104 320876 434110
rect 320824 434046 320876 434052
rect 321112 432290 321140 436902
rect 321572 432290 321600 476478
rect 321652 450764 321704 450770
rect 321652 450706 321704 450712
rect 321664 441614 321692 450706
rect 322216 441614 322244 476614
rect 327724 476400 327776 476406
rect 324226 476368 324282 476377
rect 327724 476342 327776 476348
rect 324226 476303 324282 476312
rect 324240 476270 324268 476303
rect 323584 476264 323636 476270
rect 323584 476206 323636 476212
rect 324228 476264 324280 476270
rect 324228 476206 324280 476212
rect 326986 476232 327042 476241
rect 323032 474088 323084 474094
rect 323032 474030 323084 474036
rect 323044 441614 323072 474030
rect 321664 441586 322152 441614
rect 322216 441586 322428 441614
rect 323044 441586 323440 441614
rect 322124 434602 322152 441586
rect 322124 434574 322336 434602
rect 322308 432290 322336 434574
rect 322400 434178 322428 441586
rect 322388 434172 322440 434178
rect 322388 434114 322440 434120
rect 323216 434036 323268 434042
rect 323216 433978 323268 433984
rect 320468 432262 320850 432290
rect 321112 432262 321402 432290
rect 321572 432262 322046 432290
rect 322308 432262 322690 432290
rect 323228 432276 323256 433978
rect 323412 432290 323440 441586
rect 323596 434042 323624 476206
rect 326986 476167 327042 476176
rect 327000 476134 327028 476167
rect 324964 476128 325016 476134
rect 324964 476070 325016 476076
rect 326988 476128 327040 476134
rect 326988 476070 327040 476076
rect 324320 474224 324372 474230
rect 324320 474166 324372 474172
rect 323584 434036 323636 434042
rect 323584 433978 323636 433984
rect 324332 432290 324360 474166
rect 324412 447976 324464 447982
rect 324412 447918 324464 447924
rect 324424 441614 324452 447918
rect 324424 441586 324728 441614
rect 324700 432290 324728 441586
rect 324976 434246 325004 476070
rect 327080 475516 327132 475522
rect 327080 475458 327132 475464
rect 325700 445120 325752 445126
rect 325700 445062 325752 445068
rect 325712 436694 325740 445062
rect 325792 443828 325844 443834
rect 325792 443770 325844 443776
rect 325804 436966 325832 443770
rect 325884 442468 325936 442474
rect 325884 442410 325936 442416
rect 325792 436960 325844 436966
rect 325792 436902 325844 436908
rect 325700 436688 325752 436694
rect 325700 436630 325752 436636
rect 324964 434240 325016 434246
rect 324964 434182 325016 434188
rect 325896 432290 325924 442410
rect 327092 436966 327120 475458
rect 327172 463004 327224 463010
rect 327172 462946 327224 462952
rect 326620 436960 326672 436966
rect 326620 436902 326672 436908
rect 327080 436960 327132 436966
rect 327080 436902 327132 436908
rect 325976 436688 326028 436694
rect 325976 436630 326028 436636
rect 323412 432262 323886 432290
rect 324332 432262 324438 432290
rect 324700 432262 325082 432290
rect 325726 432262 325924 432290
rect 325988 432290 326016 436630
rect 326632 432290 326660 436902
rect 327184 432290 327212 462946
rect 327736 441614 327764 476342
rect 329104 476332 329156 476338
rect 329104 476274 329156 476280
rect 328460 471300 328512 471306
rect 328460 471242 328512 471248
rect 327736 441586 327856 441614
rect 327724 436960 327776 436966
rect 327724 436902 327776 436908
rect 327736 432290 327764 436902
rect 327828 434450 327856 441586
rect 328472 436966 328500 471242
rect 328552 457564 328604 457570
rect 328552 457506 328604 457512
rect 328460 436960 328512 436966
rect 328460 436902 328512 436908
rect 327816 434444 327868 434450
rect 327816 434386 327868 434392
rect 328564 432290 328592 457506
rect 329012 436960 329064 436966
rect 329012 436902 329064 436908
rect 329024 432290 329052 436902
rect 329116 434382 329144 476274
rect 338764 476264 338816 476270
rect 338764 476206 338816 476212
rect 331864 476128 331916 476134
rect 331864 476070 331916 476076
rect 331220 451920 331272 451926
rect 331220 451862 331272 451868
rect 330024 446548 330076 446554
rect 330024 446490 330076 446496
rect 329104 434376 329156 434382
rect 329104 434318 329156 434324
rect 330036 432290 330064 446490
rect 331232 441614 331260 451862
rect 331232 441586 331352 441614
rect 330576 440972 330628 440978
rect 330576 440914 330628 440920
rect 325988 432262 326278 432290
rect 326632 432262 326922 432290
rect 327184 432262 327566 432290
rect 327736 432262 328118 432290
rect 328564 432262 328762 432290
rect 329024 432262 329314 432290
rect 329958 432262 330064 432290
rect 330588 432276 330616 440914
rect 331128 438252 331180 438258
rect 331128 438194 331180 438200
rect 331140 432276 331168 438194
rect 331324 432290 331352 441586
rect 331876 434314 331904 476070
rect 336740 475584 336792 475590
rect 336740 475526 336792 475532
rect 335360 469872 335412 469878
rect 335360 469814 335412 469820
rect 332600 468648 332652 468654
rect 332600 468590 332652 468596
rect 332324 439680 332376 439686
rect 332324 439622 332376 439628
rect 331864 434308 331916 434314
rect 331864 434250 331916 434256
rect 331324 432262 331798 432290
rect 332336 432276 332364 439622
rect 332612 432290 332640 468590
rect 333980 449336 334032 449342
rect 333980 449278 334032 449284
rect 333612 439748 333664 439754
rect 333612 439690 333664 439696
rect 332612 432262 332994 432290
rect 333624 432276 333652 439690
rect 333992 432290 334020 449278
rect 334808 439816 334860 439822
rect 334808 439758 334860 439764
rect 333992 432262 334190 432290
rect 334820 432276 334848 439758
rect 335372 434586 335400 469814
rect 335452 464500 335504 464506
rect 335452 464442 335504 464448
rect 335464 437474 335492 464442
rect 335544 447908 335596 447914
rect 335544 447850 335596 447856
rect 335556 441614 335584 447850
rect 336752 441614 336780 475526
rect 335556 441586 335768 441614
rect 336752 441586 337424 441614
rect 335464 437446 335676 437474
rect 335648 434654 335676 437446
rect 335636 434648 335688 434654
rect 335636 434590 335688 434596
rect 335360 434580 335412 434586
rect 335360 434522 335412 434528
rect 335740 432290 335768 441586
rect 337200 439544 337252 439550
rect 337200 439486 337252 439492
rect 336004 434648 336056 434654
rect 336004 434590 336056 434596
rect 335386 432262 335768 432290
rect 336016 432276 336044 434590
rect 336372 434580 336424 434586
rect 336372 434522 336424 434528
rect 336384 432290 336412 434522
rect 336384 432262 336674 432290
rect 337212 432276 337240 439486
rect 337396 432290 337424 441586
rect 338396 439612 338448 439618
rect 338396 439554 338448 439560
rect 337396 432262 337870 432290
rect 338408 432276 338436 439554
rect 338776 439550 338804 476206
rect 343640 474020 343692 474026
rect 343640 473962 343692 473968
rect 342352 470008 342404 470014
rect 342352 469950 342404 469956
rect 339592 467288 339644 467294
rect 339592 467230 339644 467236
rect 338764 439544 338816 439550
rect 338764 439486 338816 439492
rect 339040 434104 339092 434110
rect 339040 434046 339092 434052
rect 339052 432276 339080 434046
rect 339604 432290 339632 467230
rect 341064 458992 341116 458998
rect 341064 458934 341116 458940
rect 340972 453416 341024 453422
rect 340972 453358 341024 453364
rect 340236 434172 340288 434178
rect 340236 434114 340288 434120
rect 339604 432262 339710 432290
rect 340248 432276 340276 434114
rect 340984 432290 341012 453358
rect 341076 441614 341104 458934
rect 342364 441614 342392 469950
rect 341076 441586 341656 441614
rect 342364 441586 342944 441614
rect 341524 434036 341576 434042
rect 341524 433978 341576 433984
rect 340906 432262 341012 432290
rect 341536 432276 341564 433978
rect 341628 432290 341656 441586
rect 342720 434240 342772 434246
rect 342720 434182 342772 434188
rect 341628 432262 342102 432290
rect 342732 432276 342760 434182
rect 342916 432290 342944 441586
rect 343652 432290 343680 473962
rect 345204 472728 345256 472734
rect 345204 472670 345256 472676
rect 345112 454708 345164 454714
rect 345112 454650 345164 454656
rect 344560 438184 344612 438190
rect 344560 438126 344612 438132
rect 342916 432262 343298 432290
rect 343652 432262 343942 432290
rect 344572 432276 344600 438126
rect 345124 436966 345152 454650
rect 345112 436960 345164 436966
rect 345112 436902 345164 436908
rect 345216 432290 345244 472670
rect 347780 461780 347832 461786
rect 347780 461722 347832 461728
rect 346492 460352 346544 460358
rect 346492 460294 346544 460300
rect 346504 441614 346532 460294
rect 346504 441586 346624 441614
rect 345388 436960 345440 436966
rect 345388 436902 345440 436908
rect 345138 432262 345244 432290
rect 345400 432290 345428 436902
rect 346308 434444 346360 434450
rect 346308 434386 346360 434392
rect 345400 432262 345782 432290
rect 346320 432276 346348 434386
rect 346596 432290 346624 441586
rect 347596 434376 347648 434382
rect 347596 434318 347648 434324
rect 346596 432262 346978 432290
rect 347608 432276 347636 434318
rect 347792 432290 347820 461722
rect 349252 456068 349304 456074
rect 349252 456010 349304 456016
rect 348792 439544 348844 439550
rect 348792 439486 348844 439492
rect 347792 432262 348174 432290
rect 348804 432276 348832 439486
rect 349264 432290 349292 456010
rect 359476 442270 359504 563042
rect 360856 445058 360884 670686
rect 363604 590708 363656 590714
rect 363604 590650 363656 590656
rect 363616 453354 363644 590650
rect 363604 453348 363656 453354
rect 363604 453290 363656 453296
rect 364352 451994 364380 702406
rect 367744 700324 367796 700330
rect 367744 700266 367796 700272
rect 364340 451988 364392 451994
rect 364340 451930 364392 451936
rect 367756 446486 367784 700266
rect 397472 699718 397500 703520
rect 396724 699712 396776 699718
rect 396724 699654 396776 699660
rect 397460 699712 397512 699718
rect 397460 699654 397512 699660
rect 371884 696992 371936 696998
rect 371884 696934 371936 696940
rect 369124 643136 369176 643142
rect 369124 643078 369176 643084
rect 369136 454782 369164 643078
rect 369124 454776 369176 454782
rect 369124 454718 369176 454724
rect 371896 449206 371924 696934
rect 377404 630692 377456 630698
rect 377404 630634 377456 630640
rect 373264 576904 373316 576910
rect 373264 576846 373316 576852
rect 373276 472666 373304 576846
rect 373264 472660 373316 472666
rect 373264 472602 373316 472608
rect 377416 460290 377444 630634
rect 396736 468518 396764 699654
rect 396724 468512 396776 468518
rect 396724 468454 396776 468460
rect 377404 460284 377456 460290
rect 377404 460226 377456 460232
rect 371884 449200 371936 449206
rect 371884 449142 371936 449148
rect 367744 446480 367796 446486
rect 367744 446422 367796 446428
rect 360844 445052 360896 445058
rect 360844 444994 360896 445000
rect 359464 442264 359516 442270
rect 359464 442206 359516 442212
rect 412652 436898 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 429856 699718 429884 703520
rect 428464 699712 428516 699718
rect 428464 699654 428516 699660
rect 429844 699712 429896 699718
rect 429844 699654 429896 699660
rect 428476 450634 428504 699654
rect 432604 616888 432656 616894
rect 432604 616830 432656 616836
rect 428464 450628 428516 450634
rect 428464 450570 428516 450576
rect 432616 443698 432644 616830
rect 462332 456142 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 462320 456136 462372 456142
rect 462320 456078 462372 456084
rect 432604 443692 432656 443698
rect 432604 443634 432656 443640
rect 412640 436892 412692 436898
rect 412640 436834 412692 436840
rect 477512 436830 477540 702406
rect 494072 447846 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 527192 465730 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 527180 465724 527232 465730
rect 527180 465666 527232 465672
rect 494060 447840 494112 447846
rect 494060 447782 494112 447788
rect 477500 436824 477552 436830
rect 477500 436766 477552 436772
rect 542372 436762 542400 702406
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580262 683904 580318 683913
rect 580262 683839 580318 683848
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 579986 630864 580042 630873
rect 579986 630799 580042 630808
rect 580000 630698 580028 630799
rect 579988 630692 580040 630698
rect 579988 630634 580040 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580184 590714 580212 590951
rect 580172 590708 580224 590714
rect 580172 590650 580224 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563106 580212 564295
rect 580172 563100 580224 563106
rect 580172 563042 580224 563048
rect 579894 537840 579950 537849
rect 579894 537775 579950 537784
rect 579908 536858 579936 537775
rect 576124 536852 576176 536858
rect 576124 536794 576176 536800
rect 579896 536852 579948 536858
rect 579896 536794 579948 536800
rect 570604 524476 570656 524482
rect 570604 524418 570656 524424
rect 570616 458862 570644 524418
rect 574744 484424 574796 484430
rect 574744 484366 574796 484372
rect 574756 464370 574784 484366
rect 576136 467158 576164 536794
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 578882 511320 578938 511329
rect 578882 511255 578938 511264
rect 576124 467152 576176 467158
rect 576124 467094 576176 467100
rect 574744 464364 574796 464370
rect 574744 464306 574796 464312
rect 570604 458856 570656 458862
rect 570604 458798 570656 458804
rect 578896 440910 578924 511255
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 580184 470626 580212 471407
rect 580172 470620 580224 470626
rect 580172 470562 580224 470568
rect 580276 461650 580304 683839
rect 580264 461644 580316 461650
rect 580264 461586 580316 461592
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 578884 440904 578936 440910
rect 578884 440846 578936 440852
rect 542360 436756 542412 436762
rect 542360 436698 542412 436704
rect 353944 436416 353996 436422
rect 353944 436358 353996 436364
rect 352564 434512 352616 434518
rect 352564 434454 352616 434460
rect 349988 434308 350040 434314
rect 349988 434250 350040 434256
rect 349264 432262 349370 432290
rect 350000 432276 350028 434250
rect 350632 433492 350684 433498
rect 350632 433434 350684 433440
rect 350644 432276 350672 433434
rect 351184 433424 351236 433430
rect 351184 433366 351236 433372
rect 351196 432276 351224 433366
rect 351828 433356 351880 433362
rect 351828 433298 351880 433304
rect 351840 432276 351868 433298
rect 272248 431928 272300 431934
rect 272248 431870 272300 431876
rect 250536 431792 250588 431798
rect 243358 431760 243414 431769
rect 243018 431718 243358 431746
rect 250286 431740 250536 431746
rect 250286 431734 250588 431740
rect 299478 431760 299534 431769
rect 250286 431718 250576 431734
rect 243358 431695 243414 431704
rect 299534 431718 299598 431746
rect 299478 431695 299534 431704
rect 231216 398812 231268 398818
rect 231216 398754 231268 398760
rect 231124 376032 231176 376038
rect 231124 375974 231176 375980
rect 229744 374808 229796 374814
rect 229744 374750 229796 374756
rect 226984 374400 227036 374406
rect 226984 374342 227036 374348
rect 226996 310593 227024 374342
rect 228364 374332 228416 374338
rect 228364 374274 228416 374280
rect 227076 328500 227128 328506
rect 227076 328442 227128 328448
rect 226982 310584 227038 310593
rect 226982 310519 227038 310528
rect 227088 307698 227116 328442
rect 227076 307692 227128 307698
rect 227076 307634 227128 307640
rect 228376 307494 228404 374274
rect 228456 371272 228508 371278
rect 228456 371214 228508 371220
rect 228468 308718 228496 371214
rect 228548 322992 228600 322998
rect 228548 322934 228600 322940
rect 228560 309602 228588 322934
rect 228548 309596 228600 309602
rect 228548 309538 228600 309544
rect 228456 308712 228508 308718
rect 228456 308654 228508 308660
rect 229756 307766 229784 374750
rect 230020 374264 230072 374270
rect 230020 374206 230072 374212
rect 229836 374196 229888 374202
rect 229836 374138 229888 374144
rect 229848 308922 229876 374138
rect 229928 372700 229980 372706
rect 229928 372642 229980 372648
rect 229940 309097 229968 372642
rect 230032 309777 230060 374206
rect 231216 374128 231268 374134
rect 231216 374070 231268 374076
rect 231124 372768 231176 372774
rect 231124 372710 231176 372716
rect 230112 371544 230164 371550
rect 230112 371486 230164 371492
rect 230018 309768 230074 309777
rect 230018 309703 230074 309712
rect 229926 309088 229982 309097
rect 230124 309058 230152 371486
rect 230204 362976 230256 362982
rect 230204 362918 230256 362924
rect 230216 310486 230244 362918
rect 230296 357468 230348 357474
rect 230296 357410 230348 357416
rect 230204 310480 230256 310486
rect 230204 310422 230256 310428
rect 230308 309534 230336 357410
rect 230388 354748 230440 354754
rect 230388 354690 230440 354696
rect 230400 310214 230428 354690
rect 231032 320204 231084 320210
rect 231032 320146 231084 320152
rect 230940 311296 230992 311302
rect 230940 311238 230992 311244
rect 230388 310208 230440 310214
rect 230388 310150 230440 310156
rect 230952 310146 230980 311238
rect 230940 310140 230992 310146
rect 230940 310082 230992 310088
rect 230296 309528 230348 309534
rect 230296 309470 230348 309476
rect 231044 309398 231072 320146
rect 231032 309392 231084 309398
rect 231032 309334 231084 309340
rect 229926 309023 229982 309032
rect 230112 309052 230164 309058
rect 230112 308994 230164 309000
rect 229836 308916 229888 308922
rect 229836 308858 229888 308864
rect 231136 308446 231164 372710
rect 231228 310321 231256 374070
rect 231308 371476 231360 371482
rect 231308 371418 231360 371424
rect 231214 310312 231270 310321
rect 231214 310247 231270 310256
rect 231124 308440 231176 308446
rect 231320 308417 231348 371418
rect 231400 371340 231452 371346
rect 231400 371282 231452 371288
rect 231412 308854 231440 371282
rect 231490 370288 231546 370297
rect 231490 370223 231546 370232
rect 231400 308848 231452 308854
rect 231400 308790 231452 308796
rect 231504 308689 231532 370223
rect 231584 368552 231636 368558
rect 231584 368494 231636 368500
rect 231596 309466 231624 368494
rect 232228 342304 232280 342310
rect 232228 342246 232280 342252
rect 231676 339516 231728 339522
rect 231676 339458 231728 339464
rect 231688 309670 231716 339458
rect 232240 335354 232268 342246
rect 232240 335326 232360 335354
rect 231768 331288 231820 331294
rect 231768 331230 231820 331236
rect 231780 310078 231808 331230
rect 232332 325694 232360 335326
rect 231872 325666 232360 325694
rect 231872 313274 231900 325666
rect 231952 317484 232004 317490
rect 231952 317426 232004 317432
rect 231860 313268 231912 313274
rect 231860 313210 231912 313216
rect 231964 313154 231992 317426
rect 232136 314696 232188 314702
rect 232136 314638 232188 314644
rect 232044 313268 232096 313274
rect 232044 313210 232096 313216
rect 231872 313126 231992 313154
rect 231872 310457 231900 313126
rect 232056 313018 232084 313210
rect 231964 312990 232084 313018
rect 231858 310448 231914 310457
rect 231858 310383 231914 310392
rect 231860 310344 231912 310350
rect 231860 310286 231912 310292
rect 231768 310072 231820 310078
rect 231768 310014 231820 310020
rect 231676 309664 231728 309670
rect 231676 309606 231728 309612
rect 231584 309460 231636 309466
rect 231584 309402 231636 309408
rect 231490 308680 231546 308689
rect 231490 308615 231546 308624
rect 231124 308382 231176 308388
rect 231306 308408 231362 308417
rect 231306 308343 231362 308352
rect 231872 308106 231900 310286
rect 231964 309330 231992 312990
rect 232044 311908 232096 311914
rect 232044 311850 232096 311856
rect 232056 310282 232084 311850
rect 232148 310350 232176 314638
rect 232228 311228 232280 311234
rect 232228 311170 232280 311176
rect 232240 310622 232268 311170
rect 232320 311160 232372 311166
rect 232320 311102 232372 311108
rect 232228 310616 232280 310622
rect 232228 310558 232280 310564
rect 232332 310554 232360 311102
rect 233148 310616 233200 310622
rect 232778 310584 232834 310593
rect 232320 310548 232372 310554
rect 232320 310490 232372 310496
rect 232596 310548 232648 310554
rect 233148 310558 233200 310564
rect 233700 310616 233752 310622
rect 233700 310558 233752 310564
rect 232778 310519 232834 310528
rect 232964 310548 233016 310554
rect 232596 310490 232648 310496
rect 232226 310448 232282 310457
rect 232226 310383 232228 310392
rect 232280 310383 232282 310392
rect 232228 310354 232280 310360
rect 232136 310344 232188 310350
rect 232136 310286 232188 310292
rect 232044 310276 232096 310282
rect 232044 310218 232096 310224
rect 232044 310140 232096 310146
rect 232044 310082 232096 310088
rect 231952 309324 232004 309330
rect 231952 309266 232004 309272
rect 232056 308174 232084 310082
rect 232424 309126 232452 310420
rect 232516 310162 232544 310420
rect 232608 310298 232636 310490
rect 232700 310298 232728 310420
rect 232608 310270 232728 310298
rect 232792 310162 232820 310519
rect 232964 310490 233016 310496
rect 232976 310298 233004 310490
rect 233068 310298 233096 310420
rect 232976 310270 233096 310298
rect 232516 310134 232820 310162
rect 232412 309120 232464 309126
rect 232412 309062 232464 309068
rect 233160 308990 233188 310558
rect 233516 310480 233568 310486
rect 233516 310422 233568 310428
rect 233436 309058 233464 310420
rect 233528 310298 233556 310422
rect 233620 310298 233648 310420
rect 233528 310270 233648 310298
rect 233712 309126 233740 310558
rect 233700 309120 233752 309126
rect 233700 309062 233752 309068
rect 233424 309052 233476 309058
rect 233424 308994 233476 309000
rect 233148 308984 233200 308990
rect 233148 308926 233200 308932
rect 232044 308168 232096 308174
rect 232044 308110 232096 308116
rect 231860 308100 231912 308106
rect 231860 308042 231912 308048
rect 229744 307760 229796 307766
rect 229744 307702 229796 307708
rect 228364 307488 228416 307494
rect 228364 307430 228416 307436
rect 233332 306400 233384 306406
rect 233332 306342 233384 306348
rect 233344 299305 233372 306342
rect 233804 302234 233832 310420
rect 233988 309194 234016 310420
rect 233976 309188 234028 309194
rect 233976 309130 234028 309136
rect 234172 306406 234200 310420
rect 234356 309097 234384 310420
rect 234342 309088 234398 309097
rect 234342 309023 234398 309032
rect 234160 306400 234212 306406
rect 234160 306342 234212 306348
rect 233436 302206 233832 302234
rect 233436 300082 233464 302206
rect 233424 300076 233476 300082
rect 233424 300018 233476 300024
rect 233330 299296 233386 299305
rect 233330 299231 233386 299240
rect 234540 298586 234568 310420
rect 234724 299198 234752 310420
rect 234816 302734 234844 310420
rect 235000 310321 235028 310420
rect 235184 310350 235212 310420
rect 235172 310344 235224 310350
rect 234986 310312 235042 310321
rect 235172 310286 235224 310292
rect 234986 310247 235042 310256
rect 235368 309097 235396 310420
rect 235552 310010 235580 310420
rect 235540 310004 235592 310010
rect 235540 309946 235592 309952
rect 235354 309088 235410 309097
rect 235354 309023 235410 309032
rect 234804 302728 234856 302734
rect 234804 302670 234856 302676
rect 235736 302234 235764 310420
rect 235920 310282 235948 310420
rect 235908 310276 235960 310282
rect 235908 310218 235960 310224
rect 236104 304230 236132 310420
rect 236288 305454 236316 310420
rect 236472 309134 236500 310420
rect 236380 309106 236500 309134
rect 236276 305448 236328 305454
rect 236276 305390 236328 305396
rect 236380 304450 236408 309106
rect 236656 308514 236684 310420
rect 236644 308508 236696 308514
rect 236644 308450 236696 308456
rect 236840 307290 236868 310420
rect 236828 307284 236880 307290
rect 236828 307226 236880 307232
rect 236196 304422 236408 304450
rect 236092 304224 236144 304230
rect 236092 304166 236144 304172
rect 234816 302206 235764 302234
rect 234712 299192 234764 299198
rect 234712 299134 234764 299140
rect 234528 298580 234580 298586
rect 234528 298522 234580 298528
rect 234816 297770 234844 302206
rect 236196 299266 236224 304422
rect 236276 304224 236328 304230
rect 236276 304166 236328 304172
rect 236184 299260 236236 299266
rect 236184 299202 236236 299208
rect 236288 298722 236316 304166
rect 237024 303362 237052 310420
rect 236380 303334 237052 303362
rect 236276 298716 236328 298722
rect 236276 298658 236328 298664
rect 236380 297906 236408 303334
rect 236460 302728 236512 302734
rect 236460 302670 236512 302676
rect 236472 299441 236500 302670
rect 237208 300150 237236 310420
rect 237300 302734 237328 310420
rect 237380 307828 237432 307834
rect 237380 307770 237432 307776
rect 237288 302728 237340 302734
rect 237288 302670 237340 302676
rect 237392 300286 237420 307770
rect 237380 300280 237432 300286
rect 237380 300222 237432 300228
rect 237196 300144 237248 300150
rect 237196 300086 237248 300092
rect 236458 299432 236514 299441
rect 236458 299367 236514 299376
rect 237484 299334 237512 310420
rect 237668 308786 237696 310420
rect 237656 308780 237708 308786
rect 237656 308722 237708 308728
rect 237852 304502 237880 310420
rect 238036 309126 238064 310420
rect 238220 310214 238248 310420
rect 238208 310208 238260 310214
rect 238208 310150 238260 310156
rect 238404 309262 238432 310420
rect 238392 309256 238444 309262
rect 238392 309198 238444 309204
rect 238024 309120 238076 309126
rect 238024 309062 238076 309068
rect 238392 306196 238444 306202
rect 238392 306138 238444 306144
rect 238404 305318 238432 306138
rect 238392 305312 238444 305318
rect 238392 305254 238444 305260
rect 237840 304496 237892 304502
rect 237840 304438 237892 304444
rect 238588 302234 238616 310420
rect 238772 306354 238800 310420
rect 238956 309602 238984 310420
rect 238944 309596 238996 309602
rect 238944 309538 238996 309544
rect 239140 308854 239168 310420
rect 239128 308848 239180 308854
rect 239128 308790 239180 308796
rect 238772 306326 239168 306354
rect 239036 306196 239088 306202
rect 239036 306138 239088 306144
rect 238944 305448 238996 305454
rect 238944 305390 238996 305396
rect 238668 305380 238720 305386
rect 238668 305322 238720 305328
rect 237576 302206 238616 302234
rect 237472 299328 237524 299334
rect 237472 299270 237524 299276
rect 236368 297900 236420 297906
rect 236368 297842 236420 297848
rect 237576 297838 237604 302206
rect 238680 302190 238708 305322
rect 238668 302184 238720 302190
rect 238668 302126 238720 302132
rect 238956 300218 238984 305390
rect 239048 301209 239076 306138
rect 239034 301200 239090 301209
rect 239034 301135 239090 301144
rect 238944 300212 238996 300218
rect 238944 300154 238996 300160
rect 239140 298994 239168 306326
rect 239324 299402 239352 310420
rect 239402 308680 239458 308689
rect 239402 308615 239458 308624
rect 239416 308417 239444 308615
rect 239402 308408 239458 308417
rect 239402 308343 239458 308352
rect 239508 306202 239536 310420
rect 239600 308446 239628 310420
rect 239588 308440 239640 308446
rect 239588 308382 239640 308388
rect 239496 306196 239548 306202
rect 239496 306138 239548 306144
rect 239784 305386 239812 310420
rect 239968 305454 239996 310420
rect 239956 305448 240008 305454
rect 239956 305390 240008 305396
rect 239772 305380 239824 305386
rect 239772 305322 239824 305328
rect 240152 302234 240180 310420
rect 240336 306354 240364 310420
rect 240520 309641 240548 310420
rect 240506 309632 240562 309641
rect 240506 309567 240562 309576
rect 240704 307834 240732 310420
rect 240888 308990 240916 310420
rect 241072 310078 241100 310420
rect 241060 310072 241112 310078
rect 241060 310014 241112 310020
rect 240876 308984 240928 308990
rect 240876 308926 240928 308932
rect 240692 307828 240744 307834
rect 240692 307770 240744 307776
rect 241256 307698 241284 310420
rect 241440 308922 241468 310420
rect 241428 308916 241480 308922
rect 241428 308858 241480 308864
rect 241624 308378 241652 310420
rect 241612 308372 241664 308378
rect 241612 308314 241664 308320
rect 241244 307692 241296 307698
rect 241244 307634 241296 307640
rect 241808 307426 241836 310420
rect 241796 307420 241848 307426
rect 241796 307362 241848 307368
rect 241704 306400 241756 306406
rect 240336 306326 240640 306354
rect 241704 306342 241756 306348
rect 240152 302206 240364 302234
rect 239312 299396 239364 299402
rect 239312 299338 239364 299344
rect 239128 298988 239180 298994
rect 239128 298930 239180 298936
rect 237564 297832 237616 297838
rect 237564 297774 237616 297780
rect 234804 297764 234856 297770
rect 234804 297706 234856 297712
rect 240336 296682 240364 302206
rect 240612 300354 240640 306326
rect 240600 300348 240652 300354
rect 240600 300290 240652 300296
rect 241716 299470 241744 306342
rect 241992 300422 242020 310420
rect 242084 309534 242112 310420
rect 242072 309528 242124 309534
rect 242072 309470 242124 309476
rect 242268 305318 242296 310420
rect 242452 308281 242480 310420
rect 242438 308272 242494 308281
rect 242438 308207 242494 308216
rect 242636 306406 242664 310420
rect 242820 307986 242848 310420
rect 242728 307958 242848 307986
rect 242728 307562 242756 307958
rect 242808 307896 242860 307902
rect 242808 307838 242860 307844
rect 242716 307556 242768 307562
rect 242716 307498 242768 307504
rect 242624 306400 242676 306406
rect 242624 306342 242676 306348
rect 242256 305312 242308 305318
rect 242256 305254 242308 305260
rect 242820 300558 242848 307838
rect 243004 306354 243032 310420
rect 243004 306326 243124 306354
rect 242992 306196 243044 306202
rect 242992 306138 243044 306144
rect 242808 300552 242860 300558
rect 242808 300494 242860 300500
rect 241980 300416 242032 300422
rect 241980 300358 242032 300364
rect 241704 299464 241756 299470
rect 241704 299406 241756 299412
rect 243004 299130 243032 306138
rect 243096 300490 243124 306326
rect 243084 300484 243136 300490
rect 243084 300426 243136 300432
rect 242992 299124 243044 299130
rect 242992 299066 243044 299072
rect 240324 296676 240376 296682
rect 240324 296618 240376 296624
rect 243188 296614 243216 310420
rect 243372 308825 243400 310420
rect 243358 308816 243414 308825
rect 243358 308751 243414 308760
rect 243556 308394 243584 310420
rect 243740 308582 243768 310420
rect 243728 308576 243780 308582
rect 243728 308518 243780 308524
rect 243464 308366 243584 308394
rect 243464 308174 243492 308366
rect 243544 308236 243596 308242
rect 243544 308178 243596 308184
rect 243452 308168 243504 308174
rect 243452 308110 243504 308116
rect 243176 296608 243228 296614
rect 243176 296550 243228 296556
rect 225604 267708 225656 267714
rect 225604 267650 225656 267656
rect 243556 249082 243584 308178
rect 243924 307766 243952 310420
rect 243912 307760 243964 307766
rect 243912 307702 243964 307708
rect 244108 306202 244136 310420
rect 244096 306196 244148 306202
rect 244096 306138 244148 306144
rect 244292 304978 244320 310420
rect 244280 304972 244332 304978
rect 244280 304914 244332 304920
rect 244384 304434 244412 310420
rect 244568 306354 244596 310420
rect 244752 309670 244780 310420
rect 244740 309664 244792 309670
rect 244740 309606 244792 309612
rect 244568 306326 244688 306354
rect 244556 306196 244608 306202
rect 244556 306138 244608 306144
rect 244372 304428 244424 304434
rect 244372 304370 244424 304376
rect 244568 300626 244596 306138
rect 244660 300801 244688 306326
rect 244936 305998 244964 310420
rect 245120 306202 245148 310420
rect 245304 309505 245332 310420
rect 245290 309496 245346 309505
rect 245290 309431 245346 309440
rect 245488 309369 245516 310420
rect 245474 309360 245530 309369
rect 245474 309295 245530 309304
rect 245672 308650 245700 310420
rect 245660 308644 245712 308650
rect 245660 308586 245712 308592
rect 245856 307630 245884 310420
rect 245844 307624 245896 307630
rect 245844 307566 245896 307572
rect 246040 306950 246068 310420
rect 246224 309913 246252 310420
rect 246210 309904 246266 309913
rect 246210 309839 246266 309848
rect 246408 308106 246436 310420
rect 246396 308100 246448 308106
rect 246396 308042 246448 308048
rect 246028 306944 246080 306950
rect 246028 306886 246080 306892
rect 246592 306490 246620 310420
rect 245856 306462 246620 306490
rect 245108 306196 245160 306202
rect 245108 306138 245160 306144
rect 244924 305992 244976 305998
rect 244924 305934 244976 305940
rect 244646 300792 244702 300801
rect 244646 300727 244702 300736
rect 244556 300620 244608 300626
rect 244556 300562 244608 300568
rect 245856 297158 245884 306462
rect 246776 306354 246804 310420
rect 246868 309777 246896 310420
rect 246854 309768 246910 309777
rect 246854 309703 246910 309712
rect 247052 308961 247080 310420
rect 247038 308952 247094 308961
rect 247038 308887 247094 308896
rect 246948 308780 247000 308786
rect 246948 308722 247000 308728
rect 246856 308168 246908 308174
rect 246856 308110 246908 308116
rect 246132 306326 246804 306354
rect 246132 299062 246160 306326
rect 246868 306218 246896 308110
rect 246316 306190 246896 306218
rect 246120 299056 246172 299062
rect 246120 298998 246172 299004
rect 245844 297152 245896 297158
rect 245844 297094 245896 297100
rect 246316 250510 246344 306190
rect 246960 302234 246988 308722
rect 247040 307828 247092 307834
rect 247040 307770 247092 307776
rect 246408 302206 246988 302234
rect 246408 279546 246436 302206
rect 247052 300762 247080 307770
rect 247132 306400 247184 306406
rect 247132 306342 247184 306348
rect 247236 306354 247264 310420
rect 247040 300756 247092 300762
rect 247040 300698 247092 300704
rect 247144 296546 247172 306342
rect 247236 306326 247356 306354
rect 247224 304972 247276 304978
rect 247224 304914 247276 304920
rect 247236 297974 247264 304914
rect 247328 298654 247356 306326
rect 247316 298648 247368 298654
rect 247316 298590 247368 298596
rect 247224 297968 247276 297974
rect 247224 297910 247276 297916
rect 247132 296540 247184 296546
rect 247132 296482 247184 296488
rect 247420 296478 247448 310420
rect 247604 304366 247632 310420
rect 247788 309466 247816 310420
rect 247776 309460 247828 309466
rect 247776 309402 247828 309408
rect 247972 306406 248000 310420
rect 247960 306400 248012 306406
rect 247960 306342 248012 306348
rect 247592 304360 247644 304366
rect 247592 304302 247644 304308
rect 248156 302234 248184 310420
rect 248340 310350 248368 310420
rect 248328 310344 248380 310350
rect 248328 310286 248380 310292
rect 248524 309398 248552 310420
rect 248512 309392 248564 309398
rect 248512 309334 248564 309340
rect 248708 307494 248736 310420
rect 248696 307488 248748 307494
rect 248696 307430 248748 307436
rect 248604 306468 248656 306474
rect 248604 306410 248656 306416
rect 247512 302206 248184 302234
rect 247512 297090 247540 302206
rect 248616 300694 248644 306410
rect 248696 306400 248748 306406
rect 248696 306342 248748 306348
rect 248604 300688 248656 300694
rect 248604 300630 248656 300636
rect 248708 298790 248736 306342
rect 248892 300830 248920 310420
rect 249076 308854 249104 310420
rect 249064 308848 249116 308854
rect 249064 308790 249116 308796
rect 249064 307964 249116 307970
rect 249064 307906 249116 307912
rect 248880 300824 248932 300830
rect 248880 300766 248932 300772
rect 248696 298784 248748 298790
rect 248696 298726 248748 298732
rect 247500 297084 247552 297090
rect 247500 297026 247552 297032
rect 247408 296472 247460 296478
rect 247408 296414 247460 296420
rect 249076 283626 249104 307906
rect 249168 307358 249196 310420
rect 249156 307352 249208 307358
rect 249156 307294 249208 307300
rect 249352 306406 249380 310420
rect 249536 306474 249564 310420
rect 249524 306468 249576 306474
rect 249524 306410 249576 306416
rect 249340 306400 249392 306406
rect 249340 306342 249392 306348
rect 249720 304978 249748 310420
rect 249708 304972 249760 304978
rect 249708 304914 249760 304920
rect 249904 298926 249932 310420
rect 250088 306354 250116 310420
rect 250272 309233 250300 310420
rect 250258 309224 250314 309233
rect 250258 309159 250314 309168
rect 250456 307834 250484 310420
rect 250536 308100 250588 308106
rect 250536 308042 250588 308048
rect 250444 307828 250496 307834
rect 250444 307770 250496 307776
rect 249996 306326 250116 306354
rect 249996 301617 250024 306326
rect 250076 306196 250128 306202
rect 250076 306138 250128 306144
rect 249982 301608 250038 301617
rect 249982 301543 250038 301552
rect 249892 298920 249944 298926
rect 249892 298862 249944 298868
rect 250088 298858 250116 306138
rect 250548 305130 250576 308042
rect 250640 306202 250668 310420
rect 250824 308553 250852 310420
rect 250904 308712 250956 308718
rect 250904 308654 250956 308660
rect 250810 308544 250866 308553
rect 250810 308479 250866 308488
rect 250720 308032 250772 308038
rect 250720 307974 250772 307980
rect 250628 306196 250680 306202
rect 250628 306138 250680 306144
rect 250456 305102 250576 305130
rect 250076 298852 250128 298858
rect 250076 298794 250128 298800
rect 249064 283620 249116 283626
rect 249064 283562 249116 283568
rect 246396 279540 246448 279546
rect 246396 279482 246448 279488
rect 246304 250504 246356 250510
rect 246304 250446 246356 250452
rect 243544 249076 243596 249082
rect 243544 249018 243596 249024
rect 250456 245138 250484 305102
rect 250732 302234 250760 307974
rect 250548 302206 250760 302234
rect 250548 253230 250576 302206
rect 250916 296714 250944 308654
rect 251008 307902 251036 310420
rect 251192 308689 251220 310420
rect 251376 309330 251404 310420
rect 251364 309324 251416 309330
rect 251364 309266 251416 309272
rect 251178 308680 251234 308689
rect 251178 308615 251234 308624
rect 250996 307896 251048 307902
rect 250996 307838 251048 307844
rect 251560 307018 251588 310420
rect 251548 307012 251600 307018
rect 251548 306954 251600 306960
rect 251456 306808 251508 306814
rect 251456 306750 251508 306756
rect 251272 306400 251324 306406
rect 251272 306342 251324 306348
rect 250640 296686 250944 296714
rect 250640 260370 250668 296686
rect 250628 260364 250680 260370
rect 250628 260306 250680 260312
rect 250536 253224 250588 253230
rect 250536 253166 250588 253172
rect 251284 251870 251312 306342
rect 251364 301368 251416 301374
rect 251364 301310 251416 301316
rect 251376 260166 251404 301310
rect 251468 272542 251496 306750
rect 251548 306196 251600 306202
rect 251548 306138 251600 306144
rect 251456 272536 251508 272542
rect 251456 272478 251508 272484
rect 251364 260160 251416 260166
rect 251364 260102 251416 260108
rect 251272 251864 251324 251870
rect 251272 251806 251324 251812
rect 251560 246362 251588 306138
rect 251652 301374 251680 310420
rect 251836 308242 251864 310420
rect 251824 308236 251876 308242
rect 251824 308178 251876 308184
rect 251824 307828 251876 307834
rect 251824 307770 251876 307776
rect 251640 301368 251692 301374
rect 251640 301310 251692 301316
rect 251836 262954 251864 307770
rect 252020 303006 252048 310420
rect 252204 306202 252232 310420
rect 252284 308576 252336 308582
rect 252284 308518 252336 308524
rect 252192 306196 252244 306202
rect 252192 306138 252244 306144
rect 252008 303000 252060 303006
rect 252008 302942 252060 302948
rect 252296 302234 252324 308518
rect 252388 306406 252416 310420
rect 252572 306406 252600 310420
rect 252756 308174 252784 310420
rect 252744 308168 252796 308174
rect 252744 308110 252796 308116
rect 252744 306536 252796 306542
rect 252744 306478 252796 306484
rect 252652 306468 252704 306474
rect 252652 306410 252704 306416
rect 252376 306400 252428 306406
rect 252376 306342 252428 306348
rect 252560 306400 252612 306406
rect 252560 306342 252612 306348
rect 252112 302206 252324 302234
rect 252112 296714 252140 302206
rect 251928 296686 252140 296714
rect 251928 278050 251956 296686
rect 251916 278044 251968 278050
rect 251916 277986 251968 277992
rect 251824 262948 251876 262954
rect 251824 262890 251876 262896
rect 252664 261526 252692 306410
rect 252756 262886 252784 306478
rect 252836 306196 252888 306202
rect 252836 306138 252888 306144
rect 252848 269822 252876 306138
rect 252940 279478 252968 310420
rect 253124 302234 253152 310420
rect 253308 306474 253336 310420
rect 253296 306468 253348 306474
rect 253296 306410 253348 306416
rect 253204 306400 253256 306406
rect 253204 306342 253256 306348
rect 253032 302206 253152 302234
rect 253032 286346 253060 302206
rect 253020 286340 253072 286346
rect 253020 286282 253072 286288
rect 252928 279472 252980 279478
rect 252928 279414 252980 279420
rect 252836 269816 252888 269822
rect 252836 269758 252888 269764
rect 252744 262880 252796 262886
rect 252744 262822 252796 262828
rect 252652 261520 252704 261526
rect 252652 261462 252704 261468
rect 253216 260234 253244 306342
rect 253492 305697 253520 310420
rect 253676 306542 253704 310420
rect 253664 306536 253716 306542
rect 253664 306478 253716 306484
rect 253860 306202 253888 310420
rect 253952 306354 253980 310420
rect 254136 306524 254164 310420
rect 254320 306626 254348 310420
rect 254320 306598 254440 306626
rect 254136 306496 254348 306524
rect 253952 306326 254164 306354
rect 253848 306196 253900 306202
rect 253848 306138 253900 306144
rect 254032 306196 254084 306202
rect 254032 306138 254084 306144
rect 253478 305688 253534 305697
rect 253478 305623 253534 305632
rect 253204 260228 253256 260234
rect 253204 260170 253256 260176
rect 254044 252006 254072 306138
rect 254032 252000 254084 252006
rect 254032 251942 254084 251948
rect 254136 251938 254164 306326
rect 254320 306218 254348 306496
rect 254412 306354 254440 306598
rect 254504 306456 254532 310420
rect 254688 308038 254716 310420
rect 254676 308032 254728 308038
rect 254676 307974 254728 307980
rect 254504 306428 254624 306456
rect 254412 306326 254532 306354
rect 254320 306190 254440 306218
rect 254308 305992 254360 305998
rect 254308 305934 254360 305940
rect 254216 305448 254268 305454
rect 254216 305390 254268 305396
rect 254228 257378 254256 305390
rect 254320 260302 254348 305934
rect 254412 290494 254440 306190
rect 254400 290488 254452 290494
rect 254400 290430 254452 290436
rect 254308 260296 254360 260302
rect 254308 260238 254360 260244
rect 254216 257372 254268 257378
rect 254216 257314 254268 257320
rect 254124 251932 254176 251938
rect 254124 251874 254176 251880
rect 254504 247722 254532 306326
rect 254596 305454 254624 306428
rect 254584 305448 254636 305454
rect 254584 305390 254636 305396
rect 254872 304298 254900 310420
rect 255056 306202 255084 310420
rect 255044 306196 255096 306202
rect 255044 306138 255096 306144
rect 255240 305998 255268 310420
rect 255424 306354 255452 310420
rect 255608 306474 255636 310420
rect 255596 306468 255648 306474
rect 255596 306410 255648 306416
rect 255792 306354 255820 310420
rect 255976 307970 256004 310420
rect 255964 307964 256016 307970
rect 255964 307906 256016 307912
rect 255872 306468 255924 306474
rect 255872 306410 255924 306416
rect 255424 306326 255544 306354
rect 255228 305992 255280 305998
rect 255228 305934 255280 305940
rect 255412 305992 255464 305998
rect 255412 305934 255464 305940
rect 254860 304292 254912 304298
rect 254860 304234 254912 304240
rect 255424 256154 255452 305934
rect 255412 256148 255464 256154
rect 255412 256090 255464 256096
rect 255516 256018 255544 306326
rect 255608 306326 255820 306354
rect 255608 256086 255636 306326
rect 255688 306196 255740 306202
rect 255688 306138 255740 306144
rect 255700 257446 255728 306138
rect 255780 304156 255832 304162
rect 255780 304098 255832 304104
rect 255792 273970 255820 304098
rect 255884 300121 255912 306410
rect 256160 304162 256188 310420
rect 256344 305998 256372 310420
rect 256436 306202 256464 310420
rect 256424 306196 256476 306202
rect 256424 306138 256476 306144
rect 256332 305992 256384 305998
rect 256332 305934 256384 305940
rect 256148 304156 256200 304162
rect 256148 304098 256200 304104
rect 255870 300112 255926 300121
rect 255870 300047 255926 300056
rect 256620 296714 256648 310420
rect 256700 306400 256752 306406
rect 256700 306342 256752 306348
rect 255976 296686 256648 296714
rect 255780 273964 255832 273970
rect 255780 273906 255832 273912
rect 255688 257440 255740 257446
rect 255688 257382 255740 257388
rect 255596 256080 255648 256086
rect 255596 256022 255648 256028
rect 255504 256012 255556 256018
rect 255504 255954 255556 255960
rect 254492 247716 254544 247722
rect 254492 247658 254544 247664
rect 251548 246356 251600 246362
rect 251548 246298 251600 246304
rect 250444 245132 250496 245138
rect 250444 245074 250496 245080
rect 255976 244934 256004 296686
rect 256712 256222 256740 306342
rect 256804 305454 256832 310420
rect 256988 306354 257016 310420
rect 257172 306354 257200 310420
rect 257356 306406 257384 310420
rect 257436 307896 257488 307902
rect 257436 307838 257488 307844
rect 256896 306326 257016 306354
rect 257080 306326 257200 306354
rect 257344 306400 257396 306406
rect 257344 306342 257396 306348
rect 256792 305448 256844 305454
rect 256792 305390 256844 305396
rect 256792 305312 256844 305318
rect 256792 305254 256844 305260
rect 256804 257582 256832 305254
rect 256792 257576 256844 257582
rect 256792 257518 256844 257524
rect 256896 257514 256924 306326
rect 256976 306196 257028 306202
rect 256976 306138 257028 306144
rect 256988 264246 257016 306138
rect 257080 265674 257108 306326
rect 257160 305992 257212 305998
rect 257160 305934 257212 305940
rect 257172 282198 257200 305934
rect 257252 305448 257304 305454
rect 257252 305390 257304 305396
rect 257264 287706 257292 305390
rect 257448 302234 257476 307838
rect 257540 305318 257568 310420
rect 257724 306202 257752 310420
rect 257712 306196 257764 306202
rect 257712 306138 257764 306144
rect 257908 305998 257936 310420
rect 258092 308786 258120 310420
rect 258080 308780 258132 308786
rect 258080 308722 258132 308728
rect 258172 306468 258224 306474
rect 258172 306410 258224 306416
rect 257896 305992 257948 305998
rect 257896 305934 257948 305940
rect 257528 305312 257580 305318
rect 257528 305254 257580 305260
rect 257356 302206 257476 302234
rect 257252 287700 257304 287706
rect 257252 287642 257304 287648
rect 257160 282192 257212 282198
rect 257160 282134 257212 282140
rect 257356 271182 257384 302206
rect 257344 271176 257396 271182
rect 257344 271118 257396 271124
rect 257068 265668 257120 265674
rect 257068 265610 257120 265616
rect 256976 264240 257028 264246
rect 256976 264182 257028 264188
rect 256884 257508 256936 257514
rect 256884 257450 256936 257456
rect 256700 256216 256752 256222
rect 256700 256158 256752 256164
rect 258184 246430 258212 306410
rect 258276 306202 258304 310420
rect 258356 306400 258408 306406
rect 258356 306342 258408 306348
rect 258264 306196 258316 306202
rect 258264 306138 258316 306144
rect 258264 305992 258316 305998
rect 258264 305934 258316 305940
rect 258276 246498 258304 305934
rect 258368 248198 258396 306342
rect 258460 249150 258488 310420
rect 258644 306354 258672 310420
rect 258736 306474 258764 310420
rect 258724 306468 258776 306474
rect 258724 306410 258776 306416
rect 258920 306406 258948 310420
rect 259104 307834 259132 310420
rect 259092 307828 259144 307834
rect 259092 307770 259144 307776
rect 258552 306326 258672 306354
rect 258908 306400 258960 306406
rect 258908 306342 258960 306348
rect 258552 261594 258580 306326
rect 258632 306196 258684 306202
rect 258632 306138 258684 306144
rect 258540 261588 258592 261594
rect 258540 261530 258592 261536
rect 258448 249144 258500 249150
rect 258448 249086 258500 249092
rect 258356 248192 258408 248198
rect 258356 248134 258408 248140
rect 258264 246492 258316 246498
rect 258264 246434 258316 246440
rect 258172 246424 258224 246430
rect 258172 246366 258224 246372
rect 258644 245002 258672 306138
rect 259288 305998 259316 310420
rect 259472 306202 259500 310420
rect 259656 309134 259684 310420
rect 259656 309106 259776 309134
rect 259552 306400 259604 306406
rect 259552 306342 259604 306348
rect 259460 306196 259512 306202
rect 259460 306138 259512 306144
rect 259276 305992 259328 305998
rect 259276 305934 259328 305940
rect 259460 305448 259512 305454
rect 259460 305390 259512 305396
rect 259472 246566 259500 305390
rect 259564 247790 259592 306342
rect 259644 305992 259696 305998
rect 259644 305934 259696 305940
rect 259656 249286 259684 305934
rect 259644 249280 259696 249286
rect 259644 249222 259696 249228
rect 259748 249218 259776 309106
rect 259840 306406 259868 310420
rect 259828 306400 259880 306406
rect 259828 306342 259880 306348
rect 259920 306400 259972 306406
rect 259920 306342 259972 306348
rect 259828 306196 259880 306202
rect 259828 306138 259880 306144
rect 259840 250578 259868 306138
rect 259932 253298 259960 306342
rect 260024 305454 260052 310420
rect 260012 305448 260064 305454
rect 260012 305390 260064 305396
rect 260208 302234 260236 310420
rect 260392 305998 260420 310420
rect 260576 306406 260604 310420
rect 260564 306400 260616 306406
rect 260564 306342 260616 306348
rect 260380 305992 260432 305998
rect 260380 305934 260432 305940
rect 260024 302206 260236 302234
rect 260024 265742 260052 302206
rect 260760 296714 260788 310420
rect 260944 306354 260972 310420
rect 260116 296686 260788 296714
rect 260852 306326 260972 306354
rect 261128 306354 261156 310420
rect 261220 308990 261248 310420
rect 261208 308984 261260 308990
rect 261208 308926 261260 308932
rect 261404 306882 261432 310420
rect 261484 308984 261536 308990
rect 261484 308926 261536 308932
rect 261392 306876 261444 306882
rect 261392 306818 261444 306824
rect 261392 306672 261444 306678
rect 261392 306614 261444 306620
rect 261128 306326 261248 306354
rect 260116 267034 260144 296686
rect 260852 293282 260880 306326
rect 261116 305992 261168 305998
rect 261116 305934 261168 305940
rect 260932 305448 260984 305454
rect 260932 305390 260984 305396
rect 260840 293276 260892 293282
rect 260840 293218 260892 293224
rect 260104 267028 260156 267034
rect 260104 266970 260156 266976
rect 260012 265736 260064 265742
rect 260012 265678 260064 265684
rect 260944 253366 260972 305390
rect 261024 302524 261076 302530
rect 261024 302466 261076 302472
rect 261036 254590 261064 302466
rect 261128 265810 261156 305934
rect 261220 272610 261248 306326
rect 261300 306196 261352 306202
rect 261300 306138 261352 306144
rect 261312 276690 261340 306138
rect 261404 287774 261432 306614
rect 261392 287768 261444 287774
rect 261392 287710 261444 287716
rect 261300 276684 261352 276690
rect 261300 276626 261352 276632
rect 261208 272604 261260 272610
rect 261208 272546 261260 272552
rect 261116 265804 261168 265810
rect 261116 265746 261168 265752
rect 261024 254584 261076 254590
rect 261024 254526 261076 254532
rect 260932 253360 260984 253366
rect 260932 253302 260984 253308
rect 259920 253292 259972 253298
rect 259920 253234 259972 253240
rect 259828 250572 259880 250578
rect 259828 250514 259880 250520
rect 259736 249212 259788 249218
rect 259736 249154 259788 249160
rect 261496 247858 261524 308926
rect 261588 305454 261616 310420
rect 261772 305998 261800 310420
rect 261956 306202 261984 310420
rect 261944 306196 261996 306202
rect 261944 306138 261996 306144
rect 261760 305992 261812 305998
rect 261760 305934 261812 305940
rect 261576 305448 261628 305454
rect 261576 305390 261628 305396
rect 262140 302530 262168 310420
rect 262220 306468 262272 306474
rect 262220 306410 262272 306416
rect 262128 302524 262180 302530
rect 262128 302466 262180 302472
rect 262232 302234 262260 306410
rect 262324 304978 262352 310420
rect 262404 306400 262456 306406
rect 262404 306342 262456 306348
rect 262312 304972 262364 304978
rect 262312 304914 262364 304920
rect 262232 302206 262352 302234
rect 262324 250714 262352 302206
rect 262416 252074 262444 306342
rect 262508 305046 262536 310420
rect 262692 306354 262720 310420
rect 262876 306474 262904 310420
rect 262864 306468 262916 306474
rect 262864 306410 262916 306416
rect 263060 306406 263088 310420
rect 262600 306326 262720 306354
rect 263048 306400 263100 306406
rect 263048 306342 263100 306348
rect 262496 305040 262548 305046
rect 262496 304982 262548 304988
rect 262496 304904 262548 304910
rect 262496 304846 262548 304852
rect 262508 253434 262536 304846
rect 262600 254658 262628 306326
rect 263244 305130 263272 310420
rect 263428 307902 263456 310420
rect 263416 307896 263468 307902
rect 263416 307838 263468 307844
rect 262692 305102 263272 305130
rect 262692 256290 262720 305102
rect 262864 305040 262916 305046
rect 262864 304982 262916 304988
rect 262772 304972 262824 304978
rect 262772 304914 262824 304920
rect 262784 264314 262812 304914
rect 262772 264308 262824 264314
rect 262772 264250 262824 264256
rect 262680 256284 262732 256290
rect 262680 256226 262732 256232
rect 262588 254652 262640 254658
rect 262588 254594 262640 254600
rect 262496 253428 262548 253434
rect 262496 253370 262548 253376
rect 262404 252068 262456 252074
rect 262404 252010 262456 252016
rect 262312 250708 262364 250714
rect 262312 250650 262364 250656
rect 262876 250646 262904 304982
rect 263520 304910 263548 310420
rect 263600 306536 263652 306542
rect 263600 306478 263652 306484
rect 263508 304904 263560 304910
rect 263508 304846 263560 304852
rect 262864 250640 262916 250646
rect 262864 250582 262916 250588
rect 263612 249354 263640 306478
rect 263704 306406 263732 310420
rect 263888 306746 263916 310420
rect 263876 306740 263928 306746
rect 263876 306682 263928 306688
rect 264072 306610 264100 310420
rect 264152 306740 264204 306746
rect 264152 306682 264204 306688
rect 263876 306604 263928 306610
rect 263876 306546 263928 306552
rect 264060 306604 264112 306610
rect 264060 306546 264112 306552
rect 263784 306468 263836 306474
rect 263784 306410 263836 306416
rect 263692 306400 263744 306406
rect 263692 306342 263744 306348
rect 263692 306196 263744 306202
rect 263692 306138 263744 306144
rect 263704 252142 263732 306138
rect 263796 254726 263824 306410
rect 263888 261662 263916 306546
rect 264164 306490 264192 306682
rect 264072 306462 264192 306490
rect 263968 305992 264020 305998
rect 263968 305934 264020 305940
rect 263980 272678 264008 305934
rect 264072 274038 264100 306462
rect 264152 306400 264204 306406
rect 264152 306342 264204 306348
rect 264164 276758 264192 306342
rect 264256 306202 264284 310420
rect 264244 306196 264296 306202
rect 264244 306138 264296 306144
rect 264440 305998 264468 310420
rect 264624 306542 264652 310420
rect 264612 306536 264664 306542
rect 264612 306478 264664 306484
rect 264808 306474 264836 310420
rect 264992 306474 265020 310420
rect 264796 306468 264848 306474
rect 264796 306410 264848 306416
rect 264980 306468 265032 306474
rect 264980 306410 265032 306416
rect 265176 306354 265204 310420
rect 264992 306326 265204 306354
rect 264428 305992 264480 305998
rect 264428 305934 264480 305940
rect 264152 276752 264204 276758
rect 264152 276694 264204 276700
rect 264060 274032 264112 274038
rect 264060 273974 264112 273980
rect 263968 272672 264020 272678
rect 263968 272614 264020 272620
rect 263876 261656 263928 261662
rect 263876 261598 263928 261604
rect 264992 254794 265020 306326
rect 265360 306218 265388 310420
rect 265440 306468 265492 306474
rect 265440 306410 265492 306416
rect 265072 306196 265124 306202
rect 265072 306138 265124 306144
rect 265176 306190 265388 306218
rect 265084 257650 265112 306138
rect 265176 258738 265204 306190
rect 265256 305992 265308 305998
rect 265256 305934 265308 305940
rect 265268 261730 265296 305934
rect 265348 305448 265400 305454
rect 265348 305390 265400 305396
rect 265360 264382 265388 305390
rect 265452 268394 265480 306410
rect 265544 268462 265572 310420
rect 265728 306202 265756 310420
rect 265716 306196 265768 306202
rect 265716 306138 265768 306144
rect 265912 305998 265940 310420
rect 265900 305992 265952 305998
rect 265900 305934 265952 305940
rect 266004 296714 266032 310420
rect 266188 305454 266216 310420
rect 266372 305998 266400 310420
rect 266556 306354 266584 310420
rect 266636 306468 266688 306474
rect 266636 306410 266688 306416
rect 266464 306326 266584 306354
rect 266360 305992 266412 305998
rect 266360 305934 266412 305940
rect 266176 305448 266228 305454
rect 266176 305390 266228 305396
rect 265636 296686 266032 296714
rect 265636 269890 265664 296686
rect 265624 269884 265676 269890
rect 265624 269826 265676 269832
rect 265532 268456 265584 268462
rect 265532 268398 265584 268404
rect 265440 268388 265492 268394
rect 265440 268330 265492 268336
rect 265348 264376 265400 264382
rect 265348 264318 265400 264324
rect 265256 261724 265308 261730
rect 265256 261666 265308 261672
rect 265164 258732 265216 258738
rect 265164 258674 265216 258680
rect 265072 257644 265124 257650
rect 265072 257586 265124 257592
rect 266464 254862 266492 306326
rect 266648 306218 266676 306410
rect 266740 306354 266768 310420
rect 266924 306474 266952 310420
rect 266912 306468 266964 306474
rect 266912 306410 266964 306416
rect 266740 306326 266952 306354
rect 266556 306190 266676 306218
rect 266728 306196 266780 306202
rect 266556 263022 266584 306190
rect 266728 306138 266780 306144
rect 266636 305448 266688 305454
rect 266636 305390 266688 305396
rect 266648 269958 266676 305390
rect 266740 276826 266768 306138
rect 266820 305992 266872 305998
rect 266820 305934 266872 305940
rect 266832 279614 266860 305934
rect 266924 284986 266952 306326
rect 267108 306202 267136 310420
rect 267096 306196 267148 306202
rect 267096 306138 267148 306144
rect 267292 305454 267320 310420
rect 267280 305448 267332 305454
rect 267280 305390 267332 305396
rect 267476 296714 267504 310420
rect 267660 308650 267688 310420
rect 267648 308644 267700 308650
rect 267648 308586 267700 308592
rect 267844 306626 267872 310420
rect 267752 306598 267872 306626
rect 267752 305386 267780 306598
rect 268028 306490 268056 310420
rect 267844 306462 268056 306490
rect 267844 305454 267872 306462
rect 268212 306354 268240 310420
rect 267936 306326 268240 306354
rect 267832 305448 267884 305454
rect 267832 305390 267884 305396
rect 267740 305380 267792 305386
rect 267740 305322 267792 305328
rect 267832 305312 267884 305318
rect 267832 305254 267884 305260
rect 267016 296686 267504 296714
rect 266912 284980 266964 284986
rect 266912 284922 266964 284928
rect 266820 279608 266872 279614
rect 266820 279550 266872 279556
rect 266728 276820 266780 276826
rect 266728 276762 266780 276768
rect 266636 269952 266688 269958
rect 266636 269894 266688 269900
rect 266544 263016 266596 263022
rect 266544 262958 266596 262964
rect 266452 254856 266504 254862
rect 266452 254798 266504 254804
rect 264980 254788 265032 254794
rect 264980 254730 265032 254736
rect 263784 254720 263836 254726
rect 263784 254662 263836 254668
rect 263692 252136 263744 252142
rect 263692 252078 263744 252084
rect 263600 249348 263652 249354
rect 263600 249290 263652 249296
rect 261484 247852 261536 247858
rect 261484 247794 261536 247800
rect 259552 247784 259604 247790
rect 259552 247726 259604 247732
rect 259460 246560 259512 246566
rect 259460 246502 259512 246508
rect 267016 245070 267044 296686
rect 267844 253502 267872 305254
rect 267936 263090 267964 306326
rect 268304 306218 268332 310420
rect 268028 306190 268332 306218
rect 268028 267102 268056 306190
rect 268488 305538 268516 310420
rect 268672 308514 268700 310420
rect 268660 308508 268712 308514
rect 268660 308450 268712 308456
rect 268120 305510 268516 305538
rect 268120 268530 268148 305510
rect 268292 305448 268344 305454
rect 268292 305390 268344 305396
rect 268200 305380 268252 305386
rect 268200 305322 268252 305328
rect 268212 280838 268240 305322
rect 268304 283694 268332 305390
rect 268856 305318 268884 310420
rect 268844 305312 268896 305318
rect 268844 305254 268896 305260
rect 269040 296714 269068 310420
rect 269224 308446 269252 310420
rect 269212 308440 269264 308446
rect 269212 308382 269264 308388
rect 269408 307018 269436 310420
rect 269592 309134 269620 310420
rect 269500 309106 269620 309134
rect 269396 307012 269448 307018
rect 269396 306954 269448 306960
rect 269500 306490 269528 309106
rect 269672 307012 269724 307018
rect 269672 306954 269724 306960
rect 269684 306762 269712 306954
rect 268396 296686 269068 296714
rect 269224 306462 269528 306490
rect 269592 306734 269712 306762
rect 268292 283688 268344 283694
rect 268292 283630 268344 283636
rect 268200 280832 268252 280838
rect 268200 280774 268252 280780
rect 268108 268524 268160 268530
rect 268108 268466 268160 268472
rect 268016 267096 268068 267102
rect 268016 267038 268068 267044
rect 267924 263084 267976 263090
rect 267924 263026 267976 263032
rect 267832 253496 267884 253502
rect 267832 253438 267884 253444
rect 268396 246634 268424 296686
rect 269224 267170 269252 306462
rect 269304 306400 269356 306406
rect 269304 306342 269356 306348
rect 269316 270026 269344 306342
rect 269488 306196 269540 306202
rect 269488 306138 269540 306144
rect 269396 305992 269448 305998
rect 269396 305934 269448 305940
rect 269408 274106 269436 305934
rect 269500 283762 269528 306138
rect 269488 283756 269540 283762
rect 269488 283698 269540 283704
rect 269396 274100 269448 274106
rect 269396 274042 269448 274048
rect 269304 270020 269356 270026
rect 269304 269962 269356 269968
rect 269212 267164 269264 267170
rect 269212 267106 269264 267112
rect 269592 253570 269620 306734
rect 269776 306474 269804 310420
rect 269764 306468 269816 306474
rect 269764 306410 269816 306416
rect 269960 306354 269988 310420
rect 270040 307828 270092 307834
rect 270040 307770 270092 307776
rect 269684 306326 269988 306354
rect 269684 296002 269712 306326
rect 270052 306218 270080 307770
rect 269776 306190 270080 306218
rect 270144 306202 270172 310420
rect 270224 308576 270276 308582
rect 270224 308518 270276 308524
rect 270132 306196 270184 306202
rect 269672 295996 269724 296002
rect 269672 295938 269724 295944
rect 269776 291854 269804 306190
rect 270132 306138 270184 306144
rect 270236 302234 270264 308518
rect 270328 305998 270356 310420
rect 270512 307834 270540 310420
rect 270592 307964 270644 307970
rect 270592 307906 270644 307912
rect 270500 307828 270552 307834
rect 270500 307770 270552 307776
rect 270316 305992 270368 305998
rect 270316 305934 270368 305940
rect 270052 302206 270264 302234
rect 270052 300257 270080 302206
rect 270038 300248 270094 300257
rect 270038 300183 270094 300192
rect 269764 291848 269816 291854
rect 269764 291790 269816 291796
rect 270604 270094 270632 307906
rect 270696 275330 270724 310420
rect 270788 282266 270816 310420
rect 270868 306400 270920 306406
rect 270868 306342 270920 306348
rect 270880 285054 270908 306342
rect 270972 306082 271000 310420
rect 271156 307970 271184 310420
rect 271144 307964 271196 307970
rect 271144 307906 271196 307912
rect 271340 306406 271368 310420
rect 271328 306400 271380 306406
rect 271328 306342 271380 306348
rect 270972 306054 271276 306082
rect 270960 305992 271012 305998
rect 270960 305934 271012 305940
rect 270972 289134 271000 305934
rect 271052 304292 271104 304298
rect 271052 304234 271104 304240
rect 270960 289128 271012 289134
rect 270960 289070 271012 289076
rect 270868 285048 270920 285054
rect 270868 284990 270920 284996
rect 270776 282260 270828 282266
rect 270776 282202 270828 282208
rect 270684 275324 270736 275330
rect 270684 275266 270736 275272
rect 270592 270088 270644 270094
rect 270592 270030 270644 270036
rect 271064 268598 271092 304234
rect 271144 299804 271196 299810
rect 271144 299746 271196 299752
rect 271156 294642 271184 299746
rect 271144 294636 271196 294642
rect 271144 294578 271196 294584
rect 271248 290562 271276 306054
rect 271524 305998 271552 310420
rect 271604 306468 271656 306474
rect 271604 306410 271656 306416
rect 271512 305992 271564 305998
rect 271512 305934 271564 305940
rect 271616 299810 271644 306410
rect 271708 304298 271736 310420
rect 271892 306354 271920 310420
rect 272076 306474 272104 310420
rect 272064 306468 272116 306474
rect 272064 306410 272116 306416
rect 272156 306468 272208 306474
rect 272156 306410 272208 306416
rect 271892 306326 272104 306354
rect 271972 306196 272024 306202
rect 271972 306138 272024 306144
rect 271696 304292 271748 304298
rect 271696 304234 271748 304240
rect 271604 299804 271656 299810
rect 271604 299746 271656 299752
rect 271236 290556 271288 290562
rect 271236 290498 271288 290504
rect 271052 268592 271104 268598
rect 271052 268534 271104 268540
rect 271984 264450 272012 306138
rect 272076 265878 272104 306326
rect 272168 271250 272196 306410
rect 272260 280906 272288 310420
rect 272340 306400 272392 306406
rect 272340 306342 272392 306348
rect 272352 287842 272380 306342
rect 272340 287836 272392 287842
rect 272340 287778 272392 287784
rect 272248 280900 272300 280906
rect 272248 280842 272300 280848
rect 272156 271244 272208 271250
rect 272156 271186 272208 271192
rect 272064 265872 272116 265878
rect 272064 265814 272116 265820
rect 271972 264444 272024 264450
rect 271972 264386 272024 264392
rect 269580 253564 269632 253570
rect 269580 253506 269632 253512
rect 272444 250782 272472 310420
rect 272524 307896 272576 307902
rect 272524 307838 272576 307844
rect 272536 258942 272564 307838
rect 272628 296070 272656 310420
rect 272812 306474 272840 310420
rect 272800 306468 272852 306474
rect 272800 306410 272852 306416
rect 272996 306202 273024 310420
rect 273088 306406 273116 310420
rect 273272 308666 273300 310420
rect 273456 309134 273484 310420
rect 273180 308638 273300 308666
rect 273364 309106 273484 309134
rect 273180 308310 273208 308638
rect 273168 308304 273220 308310
rect 273168 308246 273220 308252
rect 273260 306468 273312 306474
rect 273260 306410 273312 306416
rect 273076 306400 273128 306406
rect 273076 306342 273128 306348
rect 272984 306196 273036 306202
rect 272984 306138 273036 306144
rect 272616 296064 272668 296070
rect 272616 296006 272668 296012
rect 273272 293350 273300 306410
rect 273364 296138 273392 309106
rect 273640 306474 273668 310420
rect 273720 308304 273772 308310
rect 273720 308246 273772 308252
rect 273628 306468 273680 306474
rect 273628 306410 273680 306416
rect 273536 306400 273588 306406
rect 273536 306342 273588 306348
rect 273444 306060 273496 306066
rect 273444 306002 273496 306008
rect 273352 296132 273404 296138
rect 273352 296074 273404 296080
rect 273260 293344 273312 293350
rect 273260 293286 273312 293292
rect 273456 271318 273484 306002
rect 273548 276894 273576 306342
rect 273732 306218 273760 308246
rect 273824 306406 273852 310420
rect 273812 306400 273864 306406
rect 273812 306342 273864 306348
rect 273640 306190 273760 306218
rect 273812 306196 273864 306202
rect 273640 278118 273668 306190
rect 273812 306138 273864 306144
rect 273720 305448 273772 305454
rect 273720 305390 273772 305396
rect 273732 286414 273760 305390
rect 273720 286408 273772 286414
rect 273720 286350 273772 286356
rect 273628 278112 273680 278118
rect 273628 278054 273680 278060
rect 273536 276888 273588 276894
rect 273536 276830 273588 276836
rect 273444 271312 273496 271318
rect 273444 271254 273496 271260
rect 272524 258936 272576 258942
rect 272524 258878 272576 258884
rect 272432 250776 272484 250782
rect 272432 250718 272484 250724
rect 273824 247926 273852 306138
rect 274008 306066 274036 310420
rect 273996 306060 274048 306066
rect 273996 306002 274048 306008
rect 274192 305454 274220 310420
rect 274180 305448 274232 305454
rect 274180 305390 274232 305396
rect 274376 296714 274404 310420
rect 274560 306202 274588 310420
rect 274744 306456 274772 310420
rect 274652 306428 274772 306456
rect 274652 306202 274680 306428
rect 274928 306354 274956 310420
rect 274744 306326 274956 306354
rect 275008 306400 275060 306406
rect 275008 306342 275060 306348
rect 275112 306354 275140 310420
rect 275296 308582 275324 310420
rect 275284 308576 275336 308582
rect 275284 308518 275336 308524
rect 275284 308032 275336 308038
rect 275284 307974 275336 307980
rect 274548 306196 274600 306202
rect 274548 306138 274600 306144
rect 274640 306196 274692 306202
rect 274640 306138 274692 306144
rect 274640 305652 274692 305658
rect 274640 305594 274692 305600
rect 274652 305454 274680 305594
rect 274640 305448 274692 305454
rect 274640 305390 274692 305396
rect 273916 296686 274404 296714
rect 273916 263158 273944 296686
rect 273904 263152 273956 263158
rect 273904 263094 273956 263100
rect 273812 247920 273864 247926
rect 273812 247862 273864 247868
rect 268384 246628 268436 246634
rect 268384 246570 268436 246576
rect 274744 245274 274772 306326
rect 274824 306060 274876 306066
rect 274824 306002 274876 306008
rect 274836 265946 274864 306002
rect 274916 305652 274968 305658
rect 274916 305594 274968 305600
rect 274928 281042 274956 305594
rect 275020 282334 275048 306342
rect 275112 306326 275232 306354
rect 275100 306196 275152 306202
rect 275100 306138 275152 306144
rect 275112 285122 275140 306138
rect 275100 285116 275152 285122
rect 275100 285058 275152 285064
rect 275008 282328 275060 282334
rect 275008 282270 275060 282276
rect 274916 281036 274968 281042
rect 274916 280978 274968 280984
rect 274824 265940 274876 265946
rect 274824 265882 274876 265888
rect 275204 245342 275232 306326
rect 275296 270162 275324 307974
rect 275376 307828 275428 307834
rect 275376 307770 275428 307776
rect 275388 302938 275416 307770
rect 275480 306406 275508 310420
rect 275468 306400 275520 306406
rect 275468 306342 275520 306348
rect 275572 306066 275600 310420
rect 275560 306060 275612 306066
rect 275560 306002 275612 306008
rect 275376 302932 275428 302938
rect 275376 302874 275428 302880
rect 275756 296714 275784 310420
rect 275940 305658 275968 310420
rect 276020 306400 276072 306406
rect 276020 306342 276072 306348
rect 275928 305652 275980 305658
rect 275928 305594 275980 305600
rect 275480 296686 275784 296714
rect 275480 294710 275508 296686
rect 275468 294704 275520 294710
rect 275468 294646 275520 294652
rect 275284 270156 275336 270162
rect 275284 270098 275336 270104
rect 276032 247994 276060 306342
rect 276124 302234 276152 310420
rect 276204 306468 276256 306474
rect 276204 306410 276256 306416
rect 276216 306116 276244 306410
rect 276308 306354 276336 310420
rect 276492 306474 276520 310420
rect 276480 306468 276532 306474
rect 276480 306410 276532 306416
rect 276308 306326 276520 306354
rect 276216 306088 276336 306116
rect 276124 302206 276244 302234
rect 276216 272746 276244 302206
rect 276308 279682 276336 306088
rect 276388 306060 276440 306066
rect 276388 306002 276440 306008
rect 276400 291922 276428 306002
rect 276492 300393 276520 306326
rect 276478 300384 276534 300393
rect 276478 300319 276534 300328
rect 276676 296714 276704 310420
rect 276860 305454 276888 310420
rect 277044 306066 277072 310420
rect 277228 306406 277256 310420
rect 277412 307834 277440 310420
rect 277400 307828 277452 307834
rect 277400 307770 277452 307776
rect 277492 306468 277544 306474
rect 277492 306410 277544 306416
rect 277216 306400 277268 306406
rect 277216 306342 277268 306348
rect 277032 306060 277084 306066
rect 277032 306002 277084 306008
rect 276848 305448 276900 305454
rect 276848 305390 276900 305396
rect 276584 296686 276704 296714
rect 276388 291916 276440 291922
rect 276388 291858 276440 291864
rect 276296 279676 276348 279682
rect 276296 279618 276348 279624
rect 276204 272740 276256 272746
rect 276204 272682 276256 272688
rect 276584 264518 276612 296686
rect 276572 264512 276624 264518
rect 276572 264454 276624 264460
rect 277504 248062 277532 306410
rect 277596 258806 277624 310420
rect 277676 306400 277728 306406
rect 277676 306342 277728 306348
rect 277688 258874 277716 306342
rect 277780 306252 277808 310420
rect 277872 306354 277900 310420
rect 278056 306406 278084 310420
rect 278136 307828 278188 307834
rect 278136 307770 278188 307776
rect 278044 306400 278096 306406
rect 277872 306326 277992 306354
rect 278044 306342 278096 306348
rect 277780 306224 277900 306252
rect 277768 306060 277820 306066
rect 277768 306002 277820 306008
rect 277780 261798 277808 306002
rect 277872 279750 277900 306224
rect 277860 279744 277912 279750
rect 277860 279686 277912 279692
rect 277768 261792 277820 261798
rect 277768 261734 277820 261740
rect 277676 258868 277728 258874
rect 277676 258810 277728 258816
rect 277584 258800 277636 258806
rect 277584 258742 277636 258748
rect 277492 248056 277544 248062
rect 277492 247998 277544 248004
rect 276020 247988 276072 247994
rect 276020 247930 276072 247936
rect 277964 246702 277992 306326
rect 278044 306196 278096 306202
rect 278044 306138 278096 306144
rect 278056 270230 278084 306138
rect 278148 275398 278176 307770
rect 278240 306066 278268 310420
rect 278320 307896 278372 307902
rect 278320 307838 278372 307844
rect 278332 306202 278360 307838
rect 278424 306474 278452 310420
rect 278608 307970 278636 310420
rect 278596 307964 278648 307970
rect 278596 307906 278648 307912
rect 278792 307834 278820 310420
rect 278780 307828 278832 307834
rect 278780 307770 278832 307776
rect 278412 306468 278464 306474
rect 278412 306410 278464 306416
rect 278872 306400 278924 306406
rect 278872 306342 278924 306348
rect 278320 306196 278372 306202
rect 278320 306138 278372 306144
rect 278228 306060 278280 306066
rect 278228 306002 278280 306008
rect 278136 275392 278188 275398
rect 278136 275334 278188 275340
rect 278044 270224 278096 270230
rect 278044 270166 278096 270172
rect 278884 249422 278912 306342
rect 278976 305658 279004 310420
rect 279160 306354 279188 310420
rect 279344 306354 279372 310420
rect 279528 306406 279556 310420
rect 279068 306326 279188 306354
rect 279252 306326 279372 306354
rect 279516 306400 279568 306406
rect 279516 306342 279568 306348
rect 278964 305652 279016 305658
rect 278964 305594 279016 305600
rect 278964 305448 279016 305454
rect 278964 305390 279016 305396
rect 278976 253706 279004 305390
rect 279068 260506 279096 306326
rect 279148 306060 279200 306066
rect 279148 306002 279200 306008
rect 279160 260574 279188 306002
rect 279252 267238 279280 306326
rect 279712 306066 279740 310420
rect 279700 306060 279752 306066
rect 279700 306002 279752 306008
rect 279896 305946 279924 310420
rect 279344 305918 279924 305946
rect 279344 268666 279372 305918
rect 279424 305652 279476 305658
rect 279424 305594 279476 305600
rect 279332 268660 279384 268666
rect 279332 268602 279384 268608
rect 279240 267232 279292 267238
rect 279240 267174 279292 267180
rect 279148 260568 279200 260574
rect 279148 260510 279200 260516
rect 279056 260500 279108 260506
rect 279056 260442 279108 260448
rect 278964 253700 279016 253706
rect 278964 253642 279016 253648
rect 278872 249416 278924 249422
rect 278872 249358 278924 249364
rect 279436 248130 279464 305594
rect 280080 305454 280108 310420
rect 280264 306354 280292 310420
rect 280356 308038 280384 310420
rect 280344 308032 280396 308038
rect 280344 307974 280396 307980
rect 280540 307086 280568 310420
rect 280528 307080 280580 307086
rect 280528 307022 280580 307028
rect 280528 306468 280580 306474
rect 280528 306410 280580 306416
rect 280436 306400 280488 306406
rect 280264 306326 280384 306354
rect 280436 306342 280488 306348
rect 280252 306196 280304 306202
rect 280252 306138 280304 306144
rect 280068 305448 280120 305454
rect 280068 305390 280120 305396
rect 280264 261934 280292 306138
rect 280252 261928 280304 261934
rect 280252 261870 280304 261876
rect 280356 261866 280384 306326
rect 280448 263226 280476 306342
rect 280540 268734 280568 306410
rect 280724 306202 280752 310420
rect 280908 307902 280936 310420
rect 280896 307896 280948 307902
rect 280896 307838 280948 307844
rect 280712 306196 280764 306202
rect 280712 306138 280764 306144
rect 281092 296714 281120 310420
rect 281276 306406 281304 310420
rect 281460 306474 281488 310420
rect 281448 306468 281500 306474
rect 281448 306410 281500 306416
rect 281264 306400 281316 306406
rect 281644 306354 281672 310420
rect 281724 306468 281776 306474
rect 281724 306410 281776 306416
rect 281264 306342 281316 306348
rect 280632 296686 281120 296714
rect 281552 306326 281672 306354
rect 280528 268728 280580 268734
rect 280528 268670 280580 268676
rect 280436 263220 280488 263226
rect 280436 263162 280488 263168
rect 280344 261860 280396 261866
rect 280344 261802 280396 261808
rect 280632 254930 280660 296686
rect 281552 254998 281580 306326
rect 281736 306252 281764 306410
rect 281828 306354 281856 310420
rect 282012 306354 282040 310420
rect 282196 306474 282224 310420
rect 282184 306468 282236 306474
rect 282184 306410 282236 306416
rect 281828 306326 281948 306354
rect 282012 306326 282224 306354
rect 281644 306224 281764 306252
rect 281644 256426 281672 306224
rect 281816 306060 281868 306066
rect 281816 306002 281868 306008
rect 281724 305448 281776 305454
rect 281724 305390 281776 305396
rect 281736 257718 281764 305390
rect 281828 264654 281856 306002
rect 281816 264648 281868 264654
rect 281816 264590 281868 264596
rect 281920 264586 281948 306326
rect 282092 306196 282144 306202
rect 282092 306138 282144 306144
rect 282000 305652 282052 305658
rect 282000 305594 282052 305600
rect 282012 265577 282040 305594
rect 282104 271454 282132 306138
rect 282092 271448 282144 271454
rect 282092 271390 282144 271396
rect 282196 271386 282224 306326
rect 282380 306066 282408 310420
rect 282564 306202 282592 310420
rect 282552 306196 282604 306202
rect 282552 306138 282604 306144
rect 282368 306060 282420 306066
rect 282368 306002 282420 306008
rect 282656 305454 282684 310420
rect 282736 306536 282788 306542
rect 282736 306478 282788 306484
rect 282748 306270 282776 306478
rect 282736 306264 282788 306270
rect 282736 306206 282788 306212
rect 282840 305658 282868 310420
rect 283024 306354 283052 310420
rect 283208 306882 283236 310420
rect 283196 306876 283248 306882
rect 283196 306818 283248 306824
rect 283392 306354 283420 310420
rect 282932 306326 283052 306354
rect 283116 306326 283420 306354
rect 282828 305652 282880 305658
rect 282828 305594 282880 305600
rect 282644 305448 282696 305454
rect 282644 305390 282696 305396
rect 282184 271380 282236 271386
rect 282184 271322 282236 271328
rect 281998 265568 282054 265577
rect 281998 265503 282054 265512
rect 281908 264580 281960 264586
rect 281908 264522 281960 264528
rect 282932 262857 282960 306326
rect 283012 306264 283064 306270
rect 283012 306206 283064 306212
rect 283024 283830 283052 306206
rect 283116 284889 283144 306326
rect 283576 306218 283604 310420
rect 283656 306876 283708 306882
rect 283656 306818 283708 306824
rect 283300 306190 283604 306218
rect 283196 306128 283248 306134
rect 283196 306070 283248 306076
rect 283208 293185 283236 306070
rect 283300 295254 283328 306190
rect 283668 306082 283696 306818
rect 283760 306134 283788 310420
rect 283944 306270 283972 310420
rect 283932 306264 283984 306270
rect 283932 306206 283984 306212
rect 283392 306054 283696 306082
rect 283748 306128 283800 306134
rect 283748 306070 283800 306076
rect 283392 301753 283420 306054
rect 284128 303249 284156 310420
rect 284312 306105 284340 310420
rect 284298 306096 284354 306105
rect 284298 306031 284354 306040
rect 284114 303240 284170 303249
rect 284114 303175 284170 303184
rect 284496 302977 284524 310420
rect 284680 303113 284708 310420
rect 284864 306241 284892 310420
rect 284850 306232 284906 306241
rect 284850 306167 284906 306176
rect 285048 303385 285076 310420
rect 285034 303376 285090 303385
rect 285034 303311 285090 303320
rect 284666 303104 284722 303113
rect 284666 303039 284722 303048
rect 284482 302968 284538 302977
rect 284482 302903 284538 302912
rect 285140 302802 285168 310420
rect 285324 305522 285352 310420
rect 285312 305516 285364 305522
rect 285312 305458 285364 305464
rect 285508 303550 285536 310420
rect 285496 303544 285548 303550
rect 285496 303486 285548 303492
rect 285692 302870 285720 310420
rect 285876 305833 285904 310420
rect 286060 306490 286088 310420
rect 285968 306462 286088 306490
rect 285862 305824 285918 305833
rect 285862 305759 285918 305768
rect 285968 303618 285996 306462
rect 286048 306332 286100 306338
rect 286048 306274 286100 306280
rect 285956 303612 286008 303618
rect 285956 303554 286008 303560
rect 285680 302864 285732 302870
rect 285680 302806 285732 302812
rect 285128 302796 285180 302802
rect 285128 302738 285180 302744
rect 283378 301744 283434 301753
rect 283378 301679 283434 301688
rect 286060 299946 286088 306274
rect 286244 302234 286272 310420
rect 286428 305590 286456 310420
rect 286416 305584 286468 305590
rect 286416 305526 286468 305532
rect 286612 303346 286640 310420
rect 286796 306338 286824 310420
rect 286784 306332 286836 306338
rect 286784 306274 286836 306280
rect 286980 305969 287008 310420
rect 286966 305960 287022 305969
rect 286966 305895 287022 305904
rect 287164 303482 287192 310420
rect 287152 303476 287204 303482
rect 287152 303418 287204 303424
rect 286600 303340 286652 303346
rect 286600 303282 286652 303288
rect 286152 302206 286272 302234
rect 287348 302234 287376 310420
rect 287440 306474 287468 310420
rect 287428 306468 287480 306474
rect 287428 306410 287480 306416
rect 287624 303278 287652 310420
rect 287612 303272 287664 303278
rect 287612 303214 287664 303220
rect 287808 303090 287836 310420
rect 287992 306066 288020 310420
rect 287980 306060 288032 306066
rect 287980 306002 288032 306008
rect 288176 303414 288204 310420
rect 288164 303408 288216 303414
rect 288164 303350 288216 303356
rect 287532 303062 287836 303090
rect 287348 302206 287468 302234
rect 286152 300529 286180 302206
rect 286138 300520 286194 300529
rect 286138 300455 286194 300464
rect 286048 299940 286100 299946
rect 286048 299882 286100 299888
rect 287440 297673 287468 302206
rect 287532 297809 287560 303062
rect 288360 302234 288388 310420
rect 288544 306202 288572 310420
rect 288532 306196 288584 306202
rect 288532 306138 288584 306144
rect 288728 302841 288756 310420
rect 288912 306354 288940 310420
rect 289096 306542 289124 310420
rect 289084 306536 289136 306542
rect 289084 306478 289136 306484
rect 288820 306326 288940 306354
rect 288714 302832 288770 302841
rect 288714 302767 288770 302776
rect 288820 302234 288848 306326
rect 288900 306264 288952 306270
rect 288900 306206 288952 306212
rect 287624 302206 288388 302234
rect 288636 302206 288848 302234
rect 287624 297945 287652 302206
rect 288636 301481 288664 302206
rect 288622 301472 288678 301481
rect 288622 301407 288678 301416
rect 287610 297936 287666 297945
rect 287610 297871 287666 297880
rect 287518 297800 287574 297809
rect 287518 297735 287574 297744
rect 287426 297664 287482 297673
rect 287426 297599 287482 297608
rect 288912 297401 288940 306206
rect 289280 297537 289308 310420
rect 289464 306270 289492 310420
rect 289452 306264 289504 306270
rect 289452 306206 289504 306212
rect 289648 305726 289676 310420
rect 289636 305720 289688 305726
rect 289636 305662 289688 305668
rect 289832 302234 289860 310420
rect 289924 306338 289952 310420
rect 289912 306332 289964 306338
rect 289912 306274 289964 306280
rect 290108 305794 290136 310420
rect 290292 306490 290320 310420
rect 290476 307222 290504 310420
rect 290464 307216 290516 307222
rect 290464 307158 290516 307164
rect 290292 306462 290504 306490
rect 290372 306332 290424 306338
rect 290372 306274 290424 306280
rect 290188 306264 290240 306270
rect 290188 306206 290240 306212
rect 290096 305788 290148 305794
rect 290096 305730 290148 305736
rect 289832 302206 290044 302234
rect 289266 297528 289322 297537
rect 289266 297463 289322 297472
rect 288898 297392 288954 297401
rect 290016 297362 290044 302206
rect 288898 297327 288954 297336
rect 290004 297356 290056 297362
rect 290004 297298 290056 297304
rect 290200 297226 290228 306206
rect 290280 306196 290332 306202
rect 290280 306138 290332 306144
rect 290292 301646 290320 306138
rect 290280 301640 290332 301646
rect 290280 301582 290332 301588
rect 290384 297634 290412 306274
rect 290476 303142 290504 306462
rect 290660 305930 290688 310420
rect 290844 306270 290872 310420
rect 290832 306264 290884 306270
rect 290832 306206 290884 306212
rect 291028 306202 291056 310420
rect 291016 306196 291068 306202
rect 291016 306138 291068 306144
rect 290648 305924 290700 305930
rect 290648 305866 290700 305872
rect 291212 305862 291240 310420
rect 291396 306406 291424 310420
rect 291580 306626 291608 310420
rect 291764 306626 291792 310420
rect 291580 306598 291700 306626
rect 291764 306598 291884 306626
rect 291384 306400 291436 306406
rect 291384 306342 291436 306348
rect 291476 306332 291528 306338
rect 291476 306274 291528 306280
rect 291200 305856 291252 305862
rect 291200 305798 291252 305804
rect 290464 303136 290516 303142
rect 290464 303078 290516 303084
rect 290372 297628 290424 297634
rect 290372 297570 290424 297576
rect 291488 297294 291516 306274
rect 291568 306264 291620 306270
rect 291568 306206 291620 306212
rect 291476 297288 291528 297294
rect 291476 297230 291528 297236
rect 290188 297220 290240 297226
rect 290188 297162 290240 297168
rect 283288 295248 283340 295254
rect 283288 295190 283340 295196
rect 291580 294846 291608 306206
rect 291672 294982 291700 306598
rect 291752 306400 291804 306406
rect 291752 306342 291804 306348
rect 291764 297702 291792 306342
rect 291856 303074 291884 306598
rect 291844 303068 291896 303074
rect 291844 303010 291896 303016
rect 291752 297696 291804 297702
rect 291752 297638 291804 297644
rect 291948 297430 291976 310420
rect 292132 306270 292160 310420
rect 292120 306264 292172 306270
rect 292120 306206 292172 306212
rect 292316 303210 292344 310420
rect 292408 306338 292436 310420
rect 292396 306332 292448 306338
rect 292396 306274 292448 306280
rect 292304 303204 292356 303210
rect 292304 303146 292356 303152
rect 291936 297424 291988 297430
rect 291936 297366 291988 297372
rect 292592 295050 292620 310420
rect 292776 306320 292804 310420
rect 292684 306292 292804 306320
rect 292856 306332 292908 306338
rect 292684 300014 292712 306292
rect 292960 306320 292988 310420
rect 293144 306320 293172 310420
rect 293328 306338 293356 310420
rect 293316 306332 293368 306338
rect 292960 306292 293080 306320
rect 293144 306292 293264 306320
rect 292856 306274 292908 306280
rect 292764 306060 292816 306066
rect 292764 306002 292816 306008
rect 292672 300008 292724 300014
rect 292672 299950 292724 299956
rect 292580 295044 292632 295050
rect 292580 294986 292632 294992
rect 291660 294976 291712 294982
rect 291660 294918 291712 294924
rect 292776 294914 292804 306002
rect 292764 294908 292816 294914
rect 292764 294850 292816 294856
rect 291568 294840 291620 294846
rect 291568 294782 291620 294788
rect 292868 294778 292896 306274
rect 292948 306128 293000 306134
rect 292948 306070 293000 306076
rect 292960 295118 292988 306070
rect 293052 295186 293080 306292
rect 293132 306196 293184 306202
rect 293132 306138 293184 306144
rect 293040 295180 293092 295186
rect 293040 295122 293092 295128
rect 292948 295112 293000 295118
rect 292948 295054 293000 295060
rect 292856 294772 292908 294778
rect 292856 294714 292908 294720
rect 283194 293176 283250 293185
rect 283194 293111 283250 293120
rect 283102 284880 283158 284889
rect 283102 284815 283158 284824
rect 283012 283824 283064 283830
rect 283012 283766 283064 283772
rect 282918 262848 282974 262857
rect 282918 262783 282974 262792
rect 281724 257712 281776 257718
rect 281724 257654 281776 257660
rect 281632 256420 281684 256426
rect 281632 256362 281684 256368
rect 281540 254992 281592 254998
rect 281540 254934 281592 254940
rect 280620 254924 280672 254930
rect 280620 254866 280672 254872
rect 279424 248124 279476 248130
rect 279424 248066 279476 248072
rect 277952 246696 278004 246702
rect 277952 246638 278004 246644
rect 275192 245336 275244 245342
rect 275192 245278 275244 245284
rect 274732 245268 274784 245274
rect 274732 245210 274784 245216
rect 267004 245064 267056 245070
rect 267004 245006 267056 245012
rect 258632 244996 258684 245002
rect 258632 244938 258684 244944
rect 255964 244928 256016 244934
rect 255964 244870 256016 244876
rect 293144 243574 293172 306138
rect 293236 243778 293264 306292
rect 293316 306274 293368 306280
rect 293512 306066 293540 310420
rect 293696 306202 293724 310420
rect 293684 306196 293736 306202
rect 293684 306138 293736 306144
rect 293880 306134 293908 310420
rect 294064 306882 294092 310420
rect 294052 306876 294104 306882
rect 294052 306818 294104 306824
rect 294052 306672 294104 306678
rect 294052 306614 294104 306620
rect 293960 306332 294012 306338
rect 293960 306274 294012 306280
rect 293868 306128 293920 306134
rect 293868 306070 293920 306076
rect 293500 306060 293552 306066
rect 293500 306002 293552 306008
rect 293224 243772 293276 243778
rect 293224 243714 293276 243720
rect 293972 243710 294000 306274
rect 293960 243704 294012 243710
rect 293960 243646 294012 243652
rect 294064 243642 294092 306614
rect 294248 306338 294276 310420
rect 294432 306490 294460 310420
rect 294616 308582 294644 310420
rect 294604 308576 294656 308582
rect 294604 308518 294656 308524
rect 294340 306462 294460 306490
rect 294236 306332 294288 306338
rect 294236 306274 294288 306280
rect 294236 306196 294288 306202
rect 294236 306138 294288 306144
rect 294144 306128 294196 306134
rect 294144 306070 294196 306076
rect 294156 300150 294184 306070
rect 294248 300529 294276 306138
rect 294340 302841 294368 306462
rect 294326 302832 294382 302841
rect 294326 302767 294382 302776
rect 294234 300520 294290 300529
rect 294234 300455 294290 300464
rect 294708 300393 294736 310420
rect 294788 308576 294840 308582
rect 294788 308518 294840 308524
rect 294694 300384 294750 300393
rect 294694 300319 294750 300328
rect 294800 300257 294828 308518
rect 294892 306202 294920 310420
rect 294880 306196 294932 306202
rect 294880 306138 294932 306144
rect 295076 305697 295104 310420
rect 295260 306134 295288 310420
rect 295340 306400 295392 306406
rect 295340 306342 295392 306348
rect 295248 306128 295300 306134
rect 295248 306070 295300 306076
rect 295062 305688 295118 305697
rect 295062 305623 295118 305632
rect 294786 300248 294842 300257
rect 294786 300183 294842 300192
rect 294144 300144 294196 300150
rect 294144 300086 294196 300092
rect 294052 243636 294104 243642
rect 294052 243578 294104 243584
rect 295352 243574 295380 306342
rect 293132 243568 293184 243574
rect 293132 243510 293184 243516
rect 295340 243568 295392 243574
rect 295444 243545 295472 310420
rect 295524 306332 295576 306338
rect 295524 306274 295576 306280
rect 295536 243642 295564 306274
rect 295628 243710 295656 310420
rect 295812 302234 295840 310420
rect 295996 308446 296024 310420
rect 295984 308440 296036 308446
rect 295984 308382 296036 308388
rect 296180 306338 296208 310420
rect 296364 306406 296392 310420
rect 296352 306400 296404 306406
rect 296352 306342 296404 306348
rect 296168 306332 296220 306338
rect 296168 306274 296220 306280
rect 295720 302206 295840 302234
rect 295720 243778 295748 302206
rect 296548 296714 296576 310420
rect 296732 306406 296760 310420
rect 296720 306400 296772 306406
rect 296720 306342 296772 306348
rect 296720 306264 296772 306270
rect 296720 306206 296772 306212
rect 295812 296686 296576 296714
rect 295812 245138 295840 296686
rect 295800 245132 295852 245138
rect 295800 245074 295852 245080
rect 296732 245002 296760 306206
rect 296916 306184 296944 310420
rect 297100 306270 297128 310420
rect 297192 309534 297220 310420
rect 297180 309528 297232 309534
rect 297180 309470 297232 309476
rect 297376 309466 297404 310420
rect 297364 309460 297416 309466
rect 297364 309402 297416 309408
rect 297180 306400 297232 306406
rect 297180 306342 297232 306348
rect 297088 306264 297140 306270
rect 297088 306206 297140 306212
rect 296916 306156 297036 306184
rect 296812 306060 296864 306066
rect 296812 306002 296864 306008
rect 296824 245274 296852 306002
rect 296904 305992 296956 305998
rect 296904 305934 296956 305940
rect 296916 245342 296944 305934
rect 297008 248033 297036 306156
rect 297192 296714 297220 306342
rect 297560 305998 297588 310420
rect 297744 306066 297772 310420
rect 297928 309262 297956 310420
rect 297916 309256 297968 309262
rect 297916 309198 297968 309204
rect 298112 306320 298140 310420
rect 298296 309330 298324 310420
rect 298284 309324 298336 309330
rect 298284 309266 298336 309272
rect 298480 308689 298508 310420
rect 298664 309398 298692 310420
rect 298652 309392 298704 309398
rect 298652 309334 298704 309340
rect 298466 308680 298522 308689
rect 298466 308615 298522 308624
rect 298848 308417 298876 310420
rect 298834 308408 298890 308417
rect 298834 308343 298890 308352
rect 298112 306292 298324 306320
rect 298100 306196 298152 306202
rect 298100 306138 298152 306144
rect 297732 306060 297784 306066
rect 297732 306002 297784 306008
rect 297548 305992 297600 305998
rect 297548 305934 297600 305940
rect 297100 296686 297220 296714
rect 296994 248024 297050 248033
rect 296994 247959 297050 247968
rect 297100 247926 297128 296686
rect 297088 247920 297140 247926
rect 297088 247862 297140 247868
rect 296904 245336 296956 245342
rect 296904 245278 296956 245284
rect 296812 245268 296864 245274
rect 296812 245210 296864 245216
rect 298112 245070 298140 306138
rect 298192 305652 298244 305658
rect 298192 305594 298244 305600
rect 298204 248169 298232 305594
rect 298296 250986 298324 306292
rect 299032 305658 299060 310420
rect 299216 309194 299244 310420
rect 299204 309188 299256 309194
rect 299204 309130 299256 309136
rect 299400 306202 299428 310420
rect 299492 306338 299520 310420
rect 299676 308553 299704 310420
rect 299662 308544 299718 308553
rect 299662 308479 299718 308488
rect 299860 306490 299888 310420
rect 299676 306462 299888 306490
rect 299480 306332 299532 306338
rect 299480 306274 299532 306280
rect 299388 306196 299440 306202
rect 299388 306138 299440 306144
rect 299572 306196 299624 306202
rect 299572 306138 299624 306144
rect 299480 306128 299532 306134
rect 299480 306070 299532 306076
rect 299020 305652 299072 305658
rect 299020 305594 299072 305600
rect 298284 250980 298336 250986
rect 298284 250922 298336 250928
rect 298190 248160 298246 248169
rect 298190 248095 298246 248104
rect 299492 245478 299520 306070
rect 299480 245472 299532 245478
rect 299480 245414 299532 245420
rect 299584 245410 299612 306138
rect 299676 245546 299704 306462
rect 299756 306332 299808 306338
rect 300044 306320 300072 310420
rect 299756 306274 299808 306280
rect 299860 306292 300072 306320
rect 299768 247654 299796 306274
rect 299860 248062 299888 306292
rect 300228 306202 300256 310420
rect 300216 306196 300268 306202
rect 300216 306138 300268 306144
rect 300412 302234 300440 310420
rect 299952 302206 300440 302234
rect 299848 248056 299900 248062
rect 299848 247998 299900 248004
rect 299952 247994 299980 302206
rect 300596 296714 300624 310420
rect 300780 306134 300808 310420
rect 300860 306604 300912 306610
rect 300860 306546 300912 306552
rect 300872 306252 300900 306546
rect 300964 306320 300992 310420
rect 301148 306406 301176 310420
rect 301332 306610 301360 310420
rect 301320 306604 301372 306610
rect 301320 306546 301372 306552
rect 301516 306490 301544 310420
rect 301240 306462 301544 306490
rect 301136 306400 301188 306406
rect 301136 306342 301188 306348
rect 300964 306292 301084 306320
rect 300872 306224 300992 306252
rect 300768 306128 300820 306134
rect 300768 306070 300820 306076
rect 300860 306060 300912 306066
rect 300860 306002 300912 306008
rect 300044 296686 300624 296714
rect 300044 250918 300072 296686
rect 300032 250912 300084 250918
rect 300032 250854 300084 250860
rect 299940 247988 299992 247994
rect 299940 247930 299992 247936
rect 299756 247648 299808 247654
rect 299756 247590 299808 247596
rect 299664 245540 299716 245546
rect 299664 245482 299716 245488
rect 299572 245404 299624 245410
rect 299572 245346 299624 245352
rect 298100 245064 298152 245070
rect 298100 245006 298152 245012
rect 296720 244996 296772 245002
rect 296720 244938 296772 244944
rect 300872 244866 300900 306002
rect 300964 245614 300992 306224
rect 301056 248198 301084 306292
rect 301240 306252 301268 306462
rect 301320 306400 301372 306406
rect 301320 306342 301372 306348
rect 301148 306224 301268 306252
rect 301044 248192 301096 248198
rect 301044 248134 301096 248140
rect 301148 248130 301176 306224
rect 301228 306128 301280 306134
rect 301228 306070 301280 306076
rect 301240 248266 301268 306070
rect 301332 251122 301360 306342
rect 301412 304700 301464 304706
rect 301412 304642 301464 304648
rect 301320 251116 301372 251122
rect 301320 251058 301372 251064
rect 301424 251054 301452 304642
rect 301700 296714 301728 310420
rect 301884 306066 301912 310420
rect 301976 306134 302004 310420
rect 301964 306128 302016 306134
rect 301964 306070 302016 306076
rect 301872 306060 301924 306066
rect 301872 306002 301924 306008
rect 302160 304706 302188 310420
rect 302344 306354 302372 310420
rect 302252 306326 302372 306354
rect 302528 306354 302556 310420
rect 302528 306326 302648 306354
rect 302148 304700 302200 304706
rect 302148 304642 302200 304648
rect 301516 296686 301728 296714
rect 301516 251190 301544 296686
rect 301504 251184 301556 251190
rect 301504 251126 301556 251132
rect 301412 251048 301464 251054
rect 301412 250990 301464 250996
rect 301228 248260 301280 248266
rect 301228 248202 301280 248208
rect 301136 248124 301188 248130
rect 301136 248066 301188 248072
rect 300952 245608 301004 245614
rect 300952 245550 301004 245556
rect 302252 245449 302280 306326
rect 302516 306264 302568 306270
rect 302516 306206 302568 306212
rect 302332 306196 302384 306202
rect 302332 306138 302384 306144
rect 302238 245440 302294 245449
rect 302238 245375 302294 245384
rect 300860 244860 300912 244866
rect 300860 244802 300912 244808
rect 302344 244798 302372 306138
rect 302424 303748 302476 303754
rect 302424 303690 302476 303696
rect 302436 245585 302464 303690
rect 302528 247586 302556 306206
rect 302620 248334 302648 306326
rect 302712 250617 302740 310420
rect 302896 303754 302924 310420
rect 303080 306270 303108 310420
rect 303068 306264 303120 306270
rect 303068 306206 303120 306212
rect 302884 303748 302936 303754
rect 302884 303690 302936 303696
rect 303264 296714 303292 310420
rect 303448 306202 303476 310420
rect 303632 306354 303660 310420
rect 303816 306490 303844 310420
rect 304000 308825 304028 310420
rect 303986 308816 304042 308825
rect 303986 308751 304042 308760
rect 303816 306462 304120 306490
rect 303988 306400 304040 306406
rect 303632 306326 303844 306354
rect 303988 306342 304040 306348
rect 303712 306264 303764 306270
rect 303712 306206 303764 306212
rect 303436 306196 303488 306202
rect 303436 306138 303488 306144
rect 303620 306196 303672 306202
rect 303620 306138 303672 306144
rect 302896 296686 303292 296714
rect 302698 250608 302754 250617
rect 302698 250543 302754 250552
rect 302896 250481 302924 296686
rect 302882 250472 302938 250481
rect 302882 250407 302938 250416
rect 302608 248328 302660 248334
rect 302608 248270 302660 248276
rect 302516 247580 302568 247586
rect 302516 247522 302568 247528
rect 303632 246265 303660 306138
rect 303724 248305 303752 306206
rect 303816 248402 303844 306326
rect 303896 306332 303948 306338
rect 303896 306274 303948 306280
rect 303908 250889 303936 306274
rect 304000 279750 304028 306342
rect 303988 279744 304040 279750
rect 303988 279686 304040 279692
rect 303894 250880 303950 250889
rect 303894 250815 303950 250824
rect 304092 250753 304120 306462
rect 304184 306270 304212 310420
rect 304276 306338 304304 310420
rect 304460 308514 304488 310420
rect 304448 308508 304500 308514
rect 304448 308450 304500 308456
rect 304264 306332 304316 306338
rect 304264 306274 304316 306280
rect 304172 306264 304224 306270
rect 304172 306206 304224 306212
rect 304644 306202 304672 310420
rect 304828 306406 304856 310420
rect 305012 306406 305040 310420
rect 305196 308718 305224 310420
rect 305380 309134 305408 310420
rect 305288 309106 305408 309134
rect 305184 308712 305236 308718
rect 305184 308654 305236 308660
rect 304816 306400 304868 306406
rect 304816 306342 304868 306348
rect 305000 306400 305052 306406
rect 305288 306354 305316 309106
rect 305460 308712 305512 308718
rect 305460 308654 305512 308660
rect 305000 306342 305052 306348
rect 305092 306332 305144 306338
rect 305092 306274 305144 306280
rect 305196 306326 305316 306354
rect 304632 306196 304684 306202
rect 304632 306138 304684 306144
rect 305000 306128 305052 306134
rect 305000 306070 305052 306076
rect 305012 265577 305040 306070
rect 305104 267073 305132 306274
rect 305196 280809 305224 306326
rect 305276 306264 305328 306270
rect 305276 306206 305328 306212
rect 305288 283529 305316 306206
rect 305368 306196 305420 306202
rect 305368 306138 305420 306144
rect 305380 294545 305408 306138
rect 305472 296041 305500 308654
rect 305564 306490 305592 310420
rect 305564 306462 305684 306490
rect 305552 306400 305604 306406
rect 305552 306342 305604 306348
rect 305564 300665 305592 306342
rect 305656 302977 305684 306462
rect 305748 306338 305776 310420
rect 305736 306332 305788 306338
rect 305736 306274 305788 306280
rect 305932 306270 305960 310420
rect 305920 306264 305972 306270
rect 305920 306206 305972 306212
rect 306116 306202 306144 310420
rect 306104 306196 306156 306202
rect 306104 306138 306156 306144
rect 306300 306134 306328 310420
rect 306484 306490 306512 310420
rect 306484 306462 306604 306490
rect 306380 306332 306432 306338
rect 306380 306274 306432 306280
rect 306288 306128 306340 306134
rect 306288 306070 306340 306076
rect 305642 302968 305698 302977
rect 305642 302903 305698 302912
rect 305550 300656 305606 300665
rect 305550 300591 305606 300600
rect 305458 296032 305514 296041
rect 305458 295967 305514 295976
rect 305366 294536 305422 294545
rect 305366 294471 305422 294480
rect 305274 283520 305330 283529
rect 305274 283455 305330 283464
rect 305182 280800 305238 280809
rect 305182 280735 305238 280744
rect 305090 267064 305146 267073
rect 305090 266999 305146 267008
rect 304998 265568 305054 265577
rect 304998 265503 305054 265512
rect 306392 263158 306420 306274
rect 306576 306218 306604 306462
rect 306668 306377 306696 310420
rect 306654 306368 306710 306377
rect 306654 306303 306710 306312
rect 306576 306190 306696 306218
rect 306564 306128 306616 306134
rect 306470 306096 306526 306105
rect 306564 306070 306616 306076
rect 306470 306031 306526 306040
rect 306380 263152 306432 263158
rect 306380 263094 306432 263100
rect 306484 262857 306512 306031
rect 306576 264586 306604 306070
rect 306668 272513 306696 306190
rect 306760 282606 306788 310420
rect 306944 307834 306972 310420
rect 306932 307828 306984 307834
rect 306932 307770 306984 307776
rect 307128 306338 307156 310420
rect 307116 306332 307168 306338
rect 307116 306274 307168 306280
rect 307312 302234 307340 310420
rect 306852 302206 307340 302234
rect 306748 282600 306800 282606
rect 306748 282542 306800 282548
rect 306852 282538 306880 302206
rect 307496 296714 307524 310420
rect 307680 306134 307708 310420
rect 307864 306474 307892 310420
rect 307852 306468 307904 306474
rect 307852 306410 307904 306416
rect 308048 306354 308076 310420
rect 307772 306326 308076 306354
rect 307668 306128 307720 306134
rect 307668 306070 307720 306076
rect 306944 296686 307524 296714
rect 306944 286686 306972 296686
rect 306932 286680 306984 286686
rect 306932 286622 306984 286628
rect 306840 282532 306892 282538
rect 306840 282474 306892 282480
rect 306654 272504 306710 272513
rect 306654 272439 306710 272448
rect 306564 264580 306616 264586
rect 306564 264522 306616 264528
rect 306470 262848 306526 262857
rect 306470 262783 306526 262792
rect 307772 254930 307800 306326
rect 308232 306218 308260 310420
rect 307864 306190 308260 306218
rect 307864 264518 307892 306190
rect 308416 305402 308444 310420
rect 308496 306468 308548 306474
rect 308496 306410 308548 306416
rect 308048 305374 308444 305402
rect 307944 305244 307996 305250
rect 307944 305186 307996 305192
rect 307956 265946 307984 305186
rect 308048 278254 308076 305374
rect 308508 305266 308536 306410
rect 308232 305238 308536 305266
rect 308128 304428 308180 304434
rect 308128 304370 308180 304376
rect 308140 283694 308168 304370
rect 308232 283762 308260 305238
rect 308600 302234 308628 310420
rect 308680 307828 308732 307834
rect 308680 307770 308732 307776
rect 308324 302206 308628 302234
rect 308324 288046 308352 302206
rect 308692 296714 308720 307770
rect 308784 305250 308812 310420
rect 308772 305244 308824 305250
rect 308772 305186 308824 305192
rect 308968 304434 308996 310420
rect 309060 307834 309088 310420
rect 309048 307828 309100 307834
rect 309048 307770 309100 307776
rect 309140 306536 309192 306542
rect 309140 306478 309192 306484
rect 308956 304428 309008 304434
rect 308956 304370 309008 304376
rect 308508 296686 308720 296714
rect 308312 288040 308364 288046
rect 308312 287982 308364 287988
rect 308508 285258 308536 296686
rect 308496 285252 308548 285258
rect 308496 285194 308548 285200
rect 308220 283756 308272 283762
rect 308220 283698 308272 283704
rect 308128 283688 308180 283694
rect 308128 283630 308180 283636
rect 308036 278248 308088 278254
rect 308036 278190 308088 278196
rect 307944 265940 307996 265946
rect 307944 265882 307996 265888
rect 307852 264512 307904 264518
rect 307852 264454 307904 264460
rect 307760 254924 307812 254930
rect 307760 254866 307812 254872
rect 309152 254862 309180 306478
rect 309244 265878 309272 310420
rect 309324 306468 309376 306474
rect 309324 306410 309376 306416
rect 309336 267306 309364 306410
rect 309428 306354 309456 310420
rect 309612 306542 309640 310420
rect 309600 306536 309652 306542
rect 309600 306478 309652 306484
rect 309796 306474 309824 310420
rect 309784 306468 309836 306474
rect 309784 306410 309836 306416
rect 309980 306354 310008 310420
rect 310060 307828 310112 307834
rect 310060 307770 310112 307776
rect 309428 306326 309640 306354
rect 309508 306264 309560 306270
rect 309508 306206 309560 306212
rect 309416 306196 309468 306202
rect 309416 306138 309468 306144
rect 309324 267300 309376 267306
rect 309324 267242 309376 267248
rect 309428 267238 309456 306138
rect 309520 275670 309548 306206
rect 309612 283626 309640 306326
rect 309704 306326 310008 306354
rect 309704 285190 309732 306326
rect 310072 302234 310100 307770
rect 310164 306270 310192 310420
rect 310152 306264 310204 306270
rect 310152 306206 310204 306212
rect 310348 306202 310376 310420
rect 310532 306626 310560 310420
rect 310532 306598 310652 306626
rect 310520 306468 310572 306474
rect 310520 306410 310572 306416
rect 310336 306196 310388 306202
rect 310336 306138 310388 306144
rect 309796 302206 310100 302234
rect 309796 287978 309824 302206
rect 309784 287972 309836 287978
rect 309784 287914 309836 287920
rect 309692 285184 309744 285190
rect 309692 285126 309744 285132
rect 309600 283620 309652 283626
rect 309600 283562 309652 283568
rect 309508 275664 309560 275670
rect 309508 275606 309560 275612
rect 310532 268734 310560 306410
rect 310624 304162 310652 306598
rect 310716 306270 310744 310420
rect 310900 306474 310928 310420
rect 310888 306468 310940 306474
rect 310888 306410 310940 306416
rect 311084 306354 311112 310420
rect 311268 308038 311296 310420
rect 311256 308032 311308 308038
rect 311256 307974 311308 307980
rect 310808 306326 311112 306354
rect 310704 306264 310756 306270
rect 310704 306206 310756 306212
rect 310704 306128 310756 306134
rect 310704 306070 310756 306076
rect 310612 304156 310664 304162
rect 310612 304098 310664 304104
rect 310612 304020 310664 304026
rect 310612 303962 310664 303968
rect 310624 270162 310652 303962
rect 310716 282470 310744 306070
rect 310808 285054 310836 306326
rect 310980 306264 311032 306270
rect 310980 306206 311032 306212
rect 310888 304156 310940 304162
rect 310888 304098 310940 304104
rect 310900 285122 310928 304098
rect 310992 286618 311020 306206
rect 311452 304026 311480 310420
rect 311544 306134 311572 310420
rect 311532 306128 311584 306134
rect 311532 306070 311584 306076
rect 311440 304020 311492 304026
rect 311440 303962 311492 303968
rect 311728 296714 311756 310420
rect 311912 308394 311940 310420
rect 312096 308394 312124 310420
rect 312280 308802 312308 310420
rect 312280 308774 312400 308802
rect 312372 308530 312400 308774
rect 312464 308666 312492 310420
rect 312464 308638 312584 308666
rect 312372 308502 312492 308530
rect 311912 308366 312032 308394
rect 312096 308366 312308 308394
rect 311900 308304 311952 308310
rect 311900 308246 311952 308252
rect 311084 296686 311756 296714
rect 311084 287842 311112 296686
rect 311072 287836 311124 287842
rect 311072 287778 311124 287784
rect 310980 286612 311032 286618
rect 310980 286554 311032 286560
rect 310888 285116 310940 285122
rect 310888 285058 310940 285064
rect 310796 285048 310848 285054
rect 310796 284990 310848 284996
rect 310704 282464 310756 282470
rect 310704 282406 310756 282412
rect 310612 270156 310664 270162
rect 310612 270098 310664 270104
rect 310520 268728 310572 268734
rect 310520 268670 310572 268676
rect 309416 267232 309468 267238
rect 309416 267174 309468 267180
rect 309232 265872 309284 265878
rect 309232 265814 309284 265820
rect 309140 254856 309192 254862
rect 309140 254798 309192 254804
rect 311912 250850 311940 308246
rect 312004 265810 312032 308366
rect 312084 308236 312136 308242
rect 312084 308178 312136 308184
rect 312096 271454 312124 308178
rect 312176 308168 312228 308174
rect 312176 308110 312228 308116
rect 312188 272678 312216 308110
rect 312280 272746 312308 308366
rect 312360 308372 312412 308378
rect 312360 308314 312412 308320
rect 312372 284986 312400 308314
rect 312464 289474 312492 308502
rect 312556 308242 312584 308638
rect 312648 308310 312676 310420
rect 312636 308304 312688 308310
rect 312636 308246 312688 308252
rect 312544 308236 312596 308242
rect 312544 308178 312596 308184
rect 312832 308122 312860 310420
rect 313016 308174 313044 310420
rect 313200 308378 313228 310420
rect 313280 308576 313332 308582
rect 313280 308518 313332 308524
rect 313188 308372 313240 308378
rect 313188 308314 313240 308320
rect 312556 308094 312860 308122
rect 313004 308168 313056 308174
rect 313004 308110 313056 308116
rect 312452 289468 312504 289474
rect 312452 289410 312504 289416
rect 312556 289338 312584 308094
rect 312636 308032 312688 308038
rect 312636 307974 312688 307980
rect 312544 289332 312596 289338
rect 312544 289274 312596 289280
rect 312648 287910 312676 307974
rect 312636 287904 312688 287910
rect 312636 287846 312688 287852
rect 312360 284980 312412 284986
rect 312360 284922 312412 284928
rect 312268 272740 312320 272746
rect 312268 272682 312320 272688
rect 312176 272672 312228 272678
rect 312176 272614 312228 272620
rect 312084 271448 312136 271454
rect 312084 271390 312136 271396
rect 311992 265804 312044 265810
rect 311992 265746 312044 265752
rect 313292 252142 313320 308518
rect 313384 308310 313412 310420
rect 313568 308394 313596 310420
rect 313476 308366 313596 308394
rect 313648 308372 313700 308378
rect 313372 308304 313424 308310
rect 313372 308246 313424 308252
rect 313372 308168 313424 308174
rect 313372 308110 313424 308116
rect 313384 256426 313412 308110
rect 313476 274310 313504 308366
rect 313648 308314 313700 308320
rect 313556 308236 313608 308242
rect 313556 308178 313608 308184
rect 313568 275534 313596 308178
rect 313660 275602 313688 308314
rect 313752 286550 313780 310420
rect 313844 289202 313872 310420
rect 314028 308378 314056 310420
rect 314212 308582 314240 310420
rect 314200 308576 314252 308582
rect 314200 308518 314252 308524
rect 314016 308372 314068 308378
rect 314016 308314 314068 308320
rect 313924 308304 313976 308310
rect 313924 308246 313976 308252
rect 313936 289270 313964 308246
rect 314396 308174 314424 310420
rect 314580 308242 314608 310420
rect 314660 308644 314712 308650
rect 314660 308586 314712 308592
rect 314568 308236 314620 308242
rect 314568 308178 314620 308184
rect 314384 308168 314436 308174
rect 314384 308110 314436 308116
rect 313924 289264 313976 289270
rect 313924 289206 313976 289212
rect 313832 289196 313884 289202
rect 313832 289138 313884 289144
rect 313740 286544 313792 286550
rect 313740 286486 313792 286492
rect 313648 275596 313700 275602
rect 313648 275538 313700 275544
rect 313556 275528 313608 275534
rect 313556 275470 313608 275476
rect 313464 274304 313516 274310
rect 313464 274246 313516 274252
rect 313372 256420 313424 256426
rect 313372 256362 313424 256368
rect 313280 252136 313332 252142
rect 313280 252078 313332 252084
rect 311900 250844 311952 250850
rect 311900 250786 311952 250792
rect 304078 250744 304134 250753
rect 304078 250679 304134 250688
rect 303804 248396 303856 248402
rect 303804 248338 303856 248344
rect 303710 248296 303766 248305
rect 303710 248231 303766 248240
rect 303618 246256 303674 246265
rect 303618 246191 303674 246200
rect 302422 245576 302478 245585
rect 302422 245511 302478 245520
rect 314672 244934 314700 308586
rect 314764 308582 314792 310420
rect 314752 308576 314804 308582
rect 314752 308518 314804 308524
rect 314844 308372 314896 308378
rect 314844 308314 314896 308320
rect 314752 308236 314804 308242
rect 314752 308178 314804 308184
rect 314764 256290 314792 308178
rect 314856 267170 314884 308314
rect 314948 308310 314976 310420
rect 315132 308394 315160 310420
rect 315212 308576 315264 308582
rect 315212 308518 315264 308524
rect 315040 308366 315160 308394
rect 314936 308304 314988 308310
rect 314936 308246 314988 308252
rect 314936 308168 314988 308174
rect 314936 308110 314988 308116
rect 314948 279682 314976 308110
rect 315040 281042 315068 308366
rect 315120 308304 315172 308310
rect 315120 308246 315172 308252
rect 315132 289406 315160 308246
rect 315224 291922 315252 308518
rect 315316 308378 315344 310420
rect 315304 308372 315356 308378
rect 315304 308314 315356 308320
rect 315500 308242 315528 310420
rect 315488 308236 315540 308242
rect 315488 308178 315540 308184
rect 315684 308174 315712 310420
rect 315868 308650 315896 310420
rect 315856 308644 315908 308650
rect 315856 308586 315908 308592
rect 316052 308242 316080 310420
rect 316236 308650 316264 310420
rect 316224 308644 316276 308650
rect 316224 308586 316276 308592
rect 316132 308576 316184 308582
rect 316328 308530 316356 310420
rect 316512 308582 316540 310420
rect 316132 308518 316184 308524
rect 316040 308236 316092 308242
rect 316040 308178 316092 308184
rect 315672 308168 315724 308174
rect 316144 308122 316172 308518
rect 315672 308110 315724 308116
rect 316052 308094 316172 308122
rect 316236 308502 316356 308530
rect 316500 308576 316552 308582
rect 316500 308518 316552 308524
rect 315212 291916 315264 291922
rect 315212 291858 315264 291864
rect 315120 289400 315172 289406
rect 315120 289342 315172 289348
rect 315028 281036 315080 281042
rect 315028 280978 315080 280984
rect 314936 279676 314988 279682
rect 314936 279618 314988 279624
rect 314844 267164 314896 267170
rect 314844 267106 314896 267112
rect 314752 256284 314804 256290
rect 314752 256226 314804 256232
rect 316052 256222 316080 308094
rect 316132 308032 316184 308038
rect 316132 307974 316184 307980
rect 316144 265742 316172 307974
rect 316236 275466 316264 308502
rect 316408 308372 316460 308378
rect 316408 308314 316460 308320
rect 316316 308304 316368 308310
rect 316316 308246 316368 308252
rect 316328 278186 316356 308246
rect 316420 280906 316448 308314
rect 316500 308236 316552 308242
rect 316500 308178 316552 308184
rect 316512 290494 316540 308178
rect 316696 307222 316724 310420
rect 316880 308038 316908 310420
rect 317064 308378 317092 310420
rect 317052 308372 317104 308378
rect 317052 308314 317104 308320
rect 317248 308310 317276 310420
rect 317432 308378 317460 310420
rect 317512 308576 317564 308582
rect 317512 308518 317564 308524
rect 317420 308372 317472 308378
rect 317420 308314 317472 308320
rect 317236 308304 317288 308310
rect 317236 308246 317288 308252
rect 317420 308236 317472 308242
rect 317420 308178 317472 308184
rect 316868 308032 316920 308038
rect 316868 307974 316920 307980
rect 316684 307216 316736 307222
rect 316684 307158 316736 307164
rect 316500 290488 316552 290494
rect 316500 290430 316552 290436
rect 316408 280900 316460 280906
rect 316408 280842 316460 280848
rect 316316 278180 316368 278186
rect 316316 278122 316368 278128
rect 316224 275460 316276 275466
rect 316224 275402 316276 275408
rect 316132 265736 316184 265742
rect 316132 265678 316184 265684
rect 316040 256216 316092 256222
rect 316040 256158 316092 256164
rect 317432 247858 317460 308178
rect 317524 250782 317552 308518
rect 317616 256154 317644 310420
rect 317696 308372 317748 308378
rect 317696 308314 317748 308320
rect 317708 263090 317736 308314
rect 317696 263084 317748 263090
rect 317696 263026 317748 263032
rect 317800 263022 317828 310420
rect 317984 308582 318012 310420
rect 317972 308576 318024 308582
rect 317972 308518 318024 308524
rect 318168 308394 318196 310420
rect 318248 308644 318300 308650
rect 318248 308586 318300 308592
rect 317880 308372 317932 308378
rect 317880 308314 317932 308320
rect 317984 308366 318196 308394
rect 317892 264450 317920 308314
rect 317984 268666 318012 308366
rect 318260 296714 318288 308586
rect 318352 308378 318380 310420
rect 318340 308372 318392 308378
rect 318340 308314 318392 308320
rect 318536 308242 318564 310420
rect 318524 308236 318576 308242
rect 318524 308178 318576 308184
rect 318628 307970 318656 310420
rect 318812 308378 318840 310420
rect 318800 308372 318852 308378
rect 318800 308314 318852 308320
rect 318996 308292 319024 310420
rect 319180 308310 319208 310420
rect 319260 308372 319312 308378
rect 319260 308314 319312 308320
rect 318904 308264 319024 308292
rect 319168 308304 319220 308310
rect 318800 308236 318852 308242
rect 318800 308178 318852 308184
rect 318616 307964 318668 307970
rect 318616 307906 318668 307912
rect 318168 296686 318288 296714
rect 318168 277030 318196 296686
rect 318156 277024 318208 277030
rect 318156 276966 318208 276972
rect 317972 268660 318024 268666
rect 317972 268602 318024 268608
rect 317880 264444 317932 264450
rect 317880 264386 317932 264392
rect 317788 263016 317840 263022
rect 317788 262958 317840 262964
rect 317604 256148 317656 256154
rect 317604 256090 317656 256096
rect 317512 250776 317564 250782
rect 317512 250718 317564 250724
rect 317420 247852 317472 247858
rect 317420 247794 317472 247800
rect 318812 247790 318840 308178
rect 318904 249354 318932 308264
rect 319168 308246 319220 308252
rect 319168 308168 319220 308174
rect 319168 308110 319220 308116
rect 318984 308100 319036 308106
rect 318984 308042 319036 308048
rect 318892 249348 318944 249354
rect 318892 249290 318944 249296
rect 318996 249286 319024 308042
rect 319076 308032 319128 308038
rect 319076 307974 319128 307980
rect 319088 252074 319116 307974
rect 319180 253570 319208 308110
rect 319272 267102 319300 308314
rect 319364 268598 319392 310420
rect 319444 308372 319496 308378
rect 319444 308314 319496 308320
rect 319456 270094 319484 308314
rect 319548 308106 319576 310420
rect 319732 308174 319760 310420
rect 319916 308378 319944 310420
rect 319904 308372 319956 308378
rect 319904 308314 319956 308320
rect 319720 308168 319772 308174
rect 319720 308110 319772 308116
rect 319536 308100 319588 308106
rect 319536 308042 319588 308048
rect 320100 308038 320128 310420
rect 320180 308304 320232 308310
rect 320180 308246 320232 308252
rect 320088 308032 320140 308038
rect 320088 307974 320140 307980
rect 319536 307964 319588 307970
rect 319536 307906 319588 307912
rect 319548 272610 319576 307906
rect 319536 272604 319588 272610
rect 319536 272546 319588 272552
rect 319444 270088 319496 270094
rect 319444 270030 319496 270036
rect 319352 268592 319404 268598
rect 319352 268534 319404 268540
rect 319260 267096 319312 267102
rect 319260 267038 319312 267044
rect 319168 253564 319220 253570
rect 319168 253506 319220 253512
rect 319076 252068 319128 252074
rect 319076 252010 319128 252016
rect 318984 249280 319036 249286
rect 318984 249222 319036 249228
rect 318800 247784 318852 247790
rect 318800 247726 318852 247732
rect 320192 245313 320220 308246
rect 320284 254794 320312 310420
rect 320364 308644 320416 308650
rect 320364 308586 320416 308592
rect 320376 261662 320404 308586
rect 320468 261730 320496 310420
rect 320652 308650 320680 310420
rect 320640 308644 320692 308650
rect 320640 308586 320692 308592
rect 320836 308530 320864 310420
rect 320652 308502 320864 308530
rect 320548 308372 320600 308378
rect 320548 308314 320600 308320
rect 320560 262954 320588 308314
rect 320652 270026 320680 308502
rect 321020 308394 321048 310420
rect 320744 308366 321048 308394
rect 321112 308378 321140 310420
rect 321100 308372 321152 308378
rect 320744 271386 320772 308366
rect 321100 308314 321152 308320
rect 321296 308310 321324 310420
rect 321284 308304 321336 308310
rect 321284 308246 321336 308252
rect 321480 296714 321508 310420
rect 321664 306338 321692 310420
rect 321848 307834 321876 310420
rect 321836 307828 321888 307834
rect 321836 307770 321888 307776
rect 321836 306400 321888 306406
rect 321836 306342 321888 306348
rect 321652 306332 321704 306338
rect 321652 306274 321704 306280
rect 321560 306264 321612 306270
rect 321560 306206 321612 306212
rect 320836 296686 321508 296714
rect 320836 274242 320864 296686
rect 320824 274236 320876 274242
rect 320824 274178 320876 274184
rect 320732 271380 320784 271386
rect 320732 271322 320784 271328
rect 320640 270020 320692 270026
rect 320640 269962 320692 269968
rect 320548 262948 320600 262954
rect 320548 262890 320600 262896
rect 320456 261724 320508 261730
rect 320456 261666 320508 261672
rect 320364 261656 320416 261662
rect 320364 261598 320416 261604
rect 320272 254788 320324 254794
rect 320272 254730 320324 254736
rect 321572 247722 321600 306206
rect 321744 306196 321796 306202
rect 321744 306138 321796 306144
rect 321652 306128 321704 306134
rect 321652 306070 321704 306076
rect 321664 261594 321692 306070
rect 321756 274174 321784 306138
rect 321848 282334 321876 306342
rect 322032 302234 322060 310420
rect 322112 306332 322164 306338
rect 322112 306274 322164 306280
rect 321940 302206 322060 302234
rect 321940 294642 321968 302206
rect 322124 300121 322152 306274
rect 322216 306202 322244 310420
rect 322204 306196 322256 306202
rect 322204 306138 322256 306144
rect 322400 306134 322428 310420
rect 322584 306406 322612 310420
rect 322572 306400 322624 306406
rect 322572 306342 322624 306348
rect 322768 306270 322796 310420
rect 322952 306474 322980 310420
rect 322940 306468 322992 306474
rect 322940 306410 322992 306416
rect 323136 306354 323164 310420
rect 323320 307290 323348 310420
rect 323308 307284 323360 307290
rect 323308 307226 323360 307232
rect 323412 306354 323440 310420
rect 323492 307284 323544 307290
rect 323492 307226 323544 307232
rect 322952 306326 323164 306354
rect 323228 306326 323440 306354
rect 322756 306264 322808 306270
rect 322756 306206 322808 306212
rect 322388 306128 322440 306134
rect 322388 306070 322440 306076
rect 322110 300112 322166 300121
rect 322110 300047 322166 300056
rect 321928 294636 321980 294642
rect 321928 294578 321980 294584
rect 321836 282328 321888 282334
rect 321836 282270 321888 282276
rect 321744 274168 321796 274174
rect 321744 274110 321796 274116
rect 321652 261588 321704 261594
rect 321652 261530 321704 261536
rect 321560 247716 321612 247722
rect 321560 247658 321612 247664
rect 320178 245304 320234 245313
rect 320178 245239 320234 245248
rect 322952 245177 322980 306326
rect 323228 306184 323256 306326
rect 323308 306264 323360 306270
rect 323308 306206 323360 306212
rect 323136 306156 323256 306184
rect 323032 306128 323084 306134
rect 323032 306070 323084 306076
rect 323044 247897 323072 306070
rect 323030 247888 323086 247897
rect 323030 247823 323086 247832
rect 322938 245168 322994 245177
rect 322938 245103 322994 245112
rect 323136 245041 323164 306156
rect 323216 306060 323268 306066
rect 323216 306002 323268 306008
rect 323228 253502 323256 306002
rect 323320 271318 323348 306206
rect 323400 306196 323452 306202
rect 323400 306138 323452 306144
rect 323412 274106 323440 306138
rect 323504 280838 323532 307226
rect 323596 306134 323624 310420
rect 323676 307828 323728 307834
rect 323676 307770 323728 307776
rect 323584 306128 323636 306134
rect 323584 306070 323636 306076
rect 323688 287774 323716 307770
rect 323780 306270 323808 310420
rect 323768 306264 323820 306270
rect 323768 306206 323820 306212
rect 323964 306066 323992 310420
rect 324148 307834 324176 310420
rect 324136 307828 324188 307834
rect 324136 307770 324188 307776
rect 324332 306354 324360 310420
rect 324240 306326 324360 306354
rect 324516 306338 324544 310420
rect 324700 306490 324728 310420
rect 324608 306462 324728 306490
rect 324504 306332 324556 306338
rect 323952 306060 324004 306066
rect 323952 306002 324004 306008
rect 324240 305930 324268 306326
rect 324504 306274 324556 306280
rect 324608 306218 324636 306462
rect 324884 306354 324912 310420
rect 324332 306190 324636 306218
rect 324700 306326 324912 306354
rect 324228 305924 324280 305930
rect 324228 305866 324280 305872
rect 323676 287768 323728 287774
rect 323676 287710 323728 287716
rect 323492 280832 323544 280838
rect 323492 280774 323544 280780
rect 323400 274100 323452 274106
rect 323400 274042 323452 274048
rect 323308 271312 323360 271318
rect 323308 271254 323360 271260
rect 323216 253496 323268 253502
rect 323216 253438 323268 253444
rect 324332 249218 324360 306190
rect 324596 306128 324648 306134
rect 324596 306070 324648 306076
rect 324412 305992 324464 305998
rect 324412 305934 324464 305940
rect 324504 305992 324556 305998
rect 324504 305934 324556 305940
rect 324424 253434 324452 305934
rect 324516 261526 324544 305934
rect 324608 269958 324636 306070
rect 324700 279614 324728 306326
rect 325068 306218 325096 310420
rect 325252 307834 325280 310420
rect 325148 307828 325200 307834
rect 325148 307770 325200 307776
rect 325240 307828 325292 307834
rect 325240 307770 325292 307776
rect 324792 306190 325096 306218
rect 324792 286414 324820 306190
rect 324872 305924 324924 305930
rect 324872 305866 324924 305872
rect 324884 287706 324912 305866
rect 325160 302234 325188 307770
rect 325436 306134 325464 310420
rect 325424 306128 325476 306134
rect 325424 306070 325476 306076
rect 325620 305998 325648 310420
rect 325804 307902 325832 310420
rect 325792 307896 325844 307902
rect 325792 307838 325844 307844
rect 325896 307018 325924 310420
rect 325884 307012 325936 307018
rect 325884 306954 325936 306960
rect 326080 306354 326108 310420
rect 326264 307086 326292 310420
rect 326252 307080 326304 307086
rect 326252 307022 326304 307028
rect 326160 307012 326212 307018
rect 326160 306954 326212 306960
rect 325804 306326 326108 306354
rect 325608 305992 325660 305998
rect 325608 305934 325660 305940
rect 325700 304904 325752 304910
rect 325700 304846 325752 304852
rect 325068 302206 325188 302234
rect 324872 287700 324924 287706
rect 324872 287642 324924 287648
rect 324780 286408 324832 286414
rect 324780 286350 324832 286356
rect 324688 279608 324740 279614
rect 324688 279550 324740 279556
rect 324596 269952 324648 269958
rect 324596 269894 324648 269900
rect 324504 261520 324556 261526
rect 324504 261462 324556 261468
rect 324412 253428 324464 253434
rect 324412 253370 324464 253376
rect 325068 250714 325096 302206
rect 325712 256086 325740 304846
rect 325804 264382 325832 306326
rect 325976 306264 326028 306270
rect 325976 306206 326028 306212
rect 325884 306196 325936 306202
rect 325884 306138 325936 306144
rect 325896 268530 325924 306138
rect 325884 268524 325936 268530
rect 325884 268466 325936 268472
rect 325988 268462 326016 306206
rect 326172 299474 326200 306954
rect 326448 306202 326476 310420
rect 326632 306270 326660 310420
rect 326620 306264 326672 306270
rect 326620 306206 326672 306212
rect 326436 306196 326488 306202
rect 326436 306138 326488 306144
rect 326816 304910 326844 310420
rect 326804 304904 326856 304910
rect 326804 304846 326856 304852
rect 326080 299446 326200 299474
rect 326080 275398 326108 299446
rect 327000 296714 327028 310420
rect 327184 306474 327212 310420
rect 327172 306468 327224 306474
rect 327172 306410 327224 306416
rect 327368 306354 327396 310420
rect 327448 306468 327500 306474
rect 327448 306410 327500 306416
rect 327080 306332 327132 306338
rect 327080 306274 327132 306280
rect 327184 306326 327396 306354
rect 326172 296686 327028 296714
rect 326172 276962 326200 296686
rect 326160 276956 326212 276962
rect 326160 276898 326212 276904
rect 326068 275392 326120 275398
rect 326068 275334 326120 275340
rect 325976 268456 326028 268462
rect 325976 268398 326028 268404
rect 325792 264376 325844 264382
rect 325792 264318 325844 264324
rect 325700 256080 325752 256086
rect 325700 256022 325752 256028
rect 325056 250708 325108 250714
rect 325056 250650 325108 250656
rect 324320 249212 324372 249218
rect 324320 249154 324372 249160
rect 327092 246634 327120 306274
rect 327184 253366 327212 306326
rect 327264 306196 327316 306202
rect 327264 306138 327316 306144
rect 327276 256018 327304 306138
rect 327356 306128 327408 306134
rect 327356 306070 327408 306076
rect 327368 267034 327396 306070
rect 327460 269890 327488 306410
rect 327552 306354 327580 310420
rect 327552 306326 327672 306354
rect 327736 306338 327764 310420
rect 327816 307828 327868 307834
rect 327816 307770 327868 307776
rect 327540 306264 327592 306270
rect 327540 306206 327592 306212
rect 327552 276894 327580 306206
rect 327644 286346 327672 306326
rect 327724 306332 327776 306338
rect 327724 306274 327776 306280
rect 327632 286340 327684 286346
rect 327632 286282 327684 286288
rect 327540 276888 327592 276894
rect 327540 276830 327592 276836
rect 327448 269884 327500 269890
rect 327448 269826 327500 269832
rect 327356 267028 327408 267034
rect 327356 266970 327408 266976
rect 327264 256012 327316 256018
rect 327264 255954 327316 255960
rect 327172 253360 327224 253366
rect 327172 253302 327224 253308
rect 327828 250646 327856 307770
rect 327920 306202 327948 310420
rect 328104 306270 328132 310420
rect 328092 306264 328144 306270
rect 328092 306206 328144 306212
rect 327908 306196 327960 306202
rect 327908 306138 327960 306144
rect 328196 306134 328224 310420
rect 328380 307834 328408 310420
rect 328368 307828 328420 307834
rect 328368 307770 328420 307776
rect 328460 306332 328512 306338
rect 328460 306274 328512 306280
rect 328184 306128 328236 306134
rect 328184 306070 328236 306076
rect 327816 250640 327868 250646
rect 327816 250582 327868 250588
rect 328472 247761 328500 306274
rect 328564 305998 328592 310420
rect 328748 306354 328776 310420
rect 328656 306326 328776 306354
rect 328552 305992 328604 305998
rect 328552 305934 328604 305940
rect 328552 305856 328604 305862
rect 328552 305798 328604 305804
rect 328564 249150 328592 305798
rect 328656 250578 328684 306326
rect 328932 306218 328960 310420
rect 329012 307896 329064 307902
rect 329012 307838 329064 307844
rect 328748 306190 328960 306218
rect 329024 306218 329052 307838
rect 329116 306338 329144 310420
rect 329104 306332 329156 306338
rect 329104 306274 329156 306280
rect 329024 306190 329144 306218
rect 328748 252006 328776 306190
rect 328828 306128 328880 306134
rect 328828 306070 328880 306076
rect 328840 257446 328868 306070
rect 328920 306060 328972 306066
rect 328920 306002 328972 306008
rect 328932 264314 328960 306002
rect 329012 305992 329064 305998
rect 329012 305934 329064 305940
rect 329024 274038 329052 305934
rect 329012 274032 329064 274038
rect 329012 273974 329064 273980
rect 328920 264308 328972 264314
rect 328920 264250 328972 264256
rect 328828 257440 328880 257446
rect 328828 257382 328880 257388
rect 329116 254726 329144 306190
rect 329300 306066 329328 310420
rect 329380 307828 329432 307834
rect 329380 307770 329432 307776
rect 329288 306060 329340 306066
rect 329288 306002 329340 306008
rect 329392 302234 329420 307770
rect 329484 306134 329512 310420
rect 329472 306128 329524 306134
rect 329472 306070 329524 306076
rect 329668 305862 329696 310420
rect 329852 306270 329880 310420
rect 330036 307970 330064 310420
rect 330024 307964 330076 307970
rect 330024 307906 330076 307912
rect 329932 306536 329984 306542
rect 329932 306478 329984 306484
rect 329840 306264 329892 306270
rect 329840 306206 329892 306212
rect 329944 306082 329972 306478
rect 330116 306468 330168 306474
rect 330116 306410 330168 306416
rect 330024 306332 330076 306338
rect 330024 306274 330076 306280
rect 329852 306054 329972 306082
rect 329656 305856 329708 305862
rect 329656 305798 329708 305804
rect 329208 302206 329420 302234
rect 329208 257514 329236 302206
rect 329852 258738 329880 306054
rect 329932 305992 329984 305998
rect 329932 305934 329984 305940
rect 329944 260370 329972 305934
rect 330036 265674 330064 306274
rect 330128 271250 330156 306410
rect 330220 275330 330248 310420
rect 330404 306474 330432 310420
rect 330588 306542 330616 310420
rect 330576 306536 330628 306542
rect 330576 306478 330628 306484
rect 330392 306468 330444 306474
rect 330392 306410 330444 306416
rect 330680 306354 330708 310420
rect 330312 306326 330708 306354
rect 330864 306338 330892 310420
rect 330852 306332 330904 306338
rect 330312 276826 330340 306326
rect 330852 306274 330904 306280
rect 330392 306264 330444 306270
rect 330392 306206 330444 306212
rect 330404 282266 330432 306206
rect 331048 305998 331076 310420
rect 331232 307834 331260 310420
rect 331220 307828 331272 307834
rect 331220 307770 331272 307776
rect 331416 306320 331444 310420
rect 331600 306490 331628 310420
rect 331232 306292 331444 306320
rect 331508 306462 331628 306490
rect 331036 305992 331088 305998
rect 331036 305934 331088 305940
rect 330392 282260 330444 282266
rect 330392 282202 330444 282208
rect 330300 276820 330352 276826
rect 330300 276762 330352 276768
rect 330208 275324 330260 275330
rect 330208 275266 330260 275272
rect 330116 271244 330168 271250
rect 330116 271186 330168 271192
rect 330024 265668 330076 265674
rect 330024 265610 330076 265616
rect 329932 260364 329984 260370
rect 329932 260306 329984 260312
rect 329840 258732 329892 258738
rect 329840 258674 329892 258680
rect 329196 257508 329248 257514
rect 329196 257450 329248 257456
rect 329104 254720 329156 254726
rect 329104 254662 329156 254668
rect 331232 253298 331260 306292
rect 331508 306252 331536 306462
rect 331784 306320 331812 310420
rect 331864 307964 331916 307970
rect 331864 307906 331916 307912
rect 331324 306224 331536 306252
rect 331600 306292 331812 306320
rect 331324 260302 331352 306224
rect 331496 306128 331548 306134
rect 331496 306070 331548 306076
rect 331404 306060 331456 306066
rect 331404 306002 331456 306008
rect 331312 260296 331364 260302
rect 331312 260238 331364 260244
rect 331416 260234 331444 306002
rect 331508 264246 331536 306070
rect 331600 273970 331628 306292
rect 331680 306196 331732 306202
rect 331680 306138 331732 306144
rect 331692 276758 331720 306138
rect 331772 305924 331824 305930
rect 331772 305866 331824 305872
rect 331784 278050 331812 305866
rect 331876 302234 331904 307906
rect 331968 306134 331996 310420
rect 331956 306128 332008 306134
rect 331956 306070 332008 306076
rect 332152 306066 332180 310420
rect 332140 306060 332192 306066
rect 332140 306002 332192 306008
rect 332336 305930 332364 310420
rect 332520 306202 332548 310420
rect 332704 306746 332732 310420
rect 332692 306740 332744 306746
rect 332692 306682 332744 306688
rect 332888 306490 332916 310420
rect 332612 306462 332916 306490
rect 332508 306196 332560 306202
rect 332508 306138 332560 306144
rect 332324 305924 332376 305930
rect 332324 305866 332376 305872
rect 331876 302206 331996 302234
rect 331772 278044 331824 278050
rect 331772 277986 331824 277992
rect 331680 276752 331732 276758
rect 331680 276694 331732 276700
rect 331588 273964 331640 273970
rect 331588 273906 331640 273912
rect 331496 264240 331548 264246
rect 331496 264182 331548 264188
rect 331404 260228 331456 260234
rect 331404 260170 331456 260176
rect 331968 258806 331996 302206
rect 331956 258800 332008 258806
rect 331956 258742 332008 258748
rect 331220 253292 331272 253298
rect 331220 253234 331272 253240
rect 328736 252000 328788 252006
rect 328736 251942 328788 251948
rect 328644 250572 328696 250578
rect 328644 250514 328696 250520
rect 328552 249144 328604 249150
rect 328552 249086 328604 249092
rect 328458 247752 328514 247761
rect 328458 247687 328514 247696
rect 327080 246628 327132 246634
rect 327080 246570 327132 246576
rect 323122 245032 323178 245041
rect 323122 244967 323178 244976
rect 314660 244928 314712 244934
rect 332612 244905 332640 306462
rect 332784 306400 332836 306406
rect 332784 306342 332836 306348
rect 332796 305980 332824 306342
rect 332980 306320 333008 310420
rect 333060 306740 333112 306746
rect 333060 306682 333112 306688
rect 333072 306354 333100 306682
rect 333164 306513 333192 310420
rect 333150 306504 333206 306513
rect 333150 306439 333206 306448
rect 333072 306326 333192 306354
rect 332704 305952 332824 305980
rect 332888 306292 333008 306320
rect 332704 251938 332732 305952
rect 332784 305856 332836 305862
rect 332784 305798 332836 305804
rect 332796 271182 332824 305798
rect 332888 276690 332916 306292
rect 333058 306232 333114 306241
rect 332968 306196 333020 306202
rect 333058 306167 333114 306176
rect 332968 306138 333020 306144
rect 332980 279546 333008 306138
rect 333072 291854 333100 306167
rect 333164 293350 333192 306326
rect 333244 306332 333296 306338
rect 333244 306274 333296 306280
rect 333256 298790 333284 306274
rect 333348 306202 333376 310420
rect 333428 307828 333480 307834
rect 333428 307770 333480 307776
rect 333336 306196 333388 306202
rect 333336 306138 333388 306144
rect 333244 298784 333296 298790
rect 333244 298726 333296 298732
rect 333152 293344 333204 293350
rect 333152 293286 333204 293292
rect 333440 292574 333468 307770
rect 333532 306474 333560 310420
rect 333520 306468 333572 306474
rect 333520 306410 333572 306416
rect 333716 306338 333744 310420
rect 333704 306332 333756 306338
rect 333704 306274 333756 306280
rect 333900 305862 333928 310420
rect 334084 306320 334112 310420
rect 333992 306292 334112 306320
rect 333888 305856 333940 305862
rect 333888 305798 333940 305804
rect 333348 292546 333468 292574
rect 333060 291848 333112 291854
rect 333060 291790 333112 291796
rect 332968 279540 333020 279546
rect 332968 279482 333020 279488
rect 333348 278118 333376 292546
rect 333336 278112 333388 278118
rect 333336 278054 333388 278060
rect 332876 276684 332928 276690
rect 332876 276626 332928 276632
rect 332784 271176 332836 271182
rect 332784 271118 332836 271124
rect 332692 251932 332744 251938
rect 332692 251874 332744 251880
rect 333992 246566 334020 306292
rect 334268 306252 334296 310420
rect 334348 306332 334400 306338
rect 334348 306274 334400 306280
rect 334084 306224 334296 306252
rect 333980 246560 334032 246566
rect 333980 246502 334032 246508
rect 334084 246498 334112 306224
rect 334164 306060 334216 306066
rect 334164 306002 334216 306008
rect 334176 247625 334204 306002
rect 334256 305992 334308 305998
rect 334256 305934 334308 305940
rect 334268 254590 334296 305934
rect 334360 254658 334388 306274
rect 334452 306218 334480 310420
rect 334636 306338 334664 310420
rect 334624 306332 334676 306338
rect 334624 306274 334676 306280
rect 334452 306190 334572 306218
rect 334440 306128 334492 306134
rect 334440 306070 334492 306076
rect 334452 269822 334480 306070
rect 334544 279478 334572 306190
rect 334820 306066 334848 310420
rect 335004 306134 335032 310420
rect 334992 306128 335044 306134
rect 334992 306070 335044 306076
rect 334808 306060 334860 306066
rect 334808 306002 334860 306008
rect 335188 305998 335216 310420
rect 335372 306490 335400 310420
rect 335280 306462 335400 306490
rect 335280 306202 335308 306462
rect 335464 306320 335492 310420
rect 335648 306320 335676 310420
rect 335832 306320 335860 310420
rect 335372 306292 335492 306320
rect 335556 306292 335676 306320
rect 335740 306292 335860 306320
rect 335268 306196 335320 306202
rect 335268 306138 335320 306144
rect 335176 305992 335228 305998
rect 335176 305934 335228 305940
rect 334532 279472 334584 279478
rect 334532 279414 334584 279420
rect 334440 269816 334492 269822
rect 334440 269758 334492 269764
rect 334348 254652 334400 254658
rect 334348 254594 334400 254600
rect 334256 254584 334308 254590
rect 334256 254526 334308 254532
rect 334162 247616 334218 247625
rect 334162 247551 334218 247560
rect 334072 246492 334124 246498
rect 334072 246434 334124 246440
rect 335372 246430 335400 306292
rect 335452 306128 335504 306134
rect 335452 306070 335504 306076
rect 335464 249082 335492 306070
rect 335556 251870 335584 306292
rect 335636 306196 335688 306202
rect 335636 306138 335688 306144
rect 335648 253230 335676 306138
rect 335740 257378 335768 306292
rect 335820 306196 335872 306202
rect 335820 306138 335872 306144
rect 335832 260166 335860 306138
rect 336016 302234 336044 310420
rect 336200 306134 336228 310420
rect 336384 306202 336412 310420
rect 336372 306196 336424 306202
rect 336372 306138 336424 306144
rect 336188 306128 336240 306134
rect 336188 306070 336240 306076
rect 335924 302206 336044 302234
rect 335924 268394 335952 302206
rect 336568 292574 336596 310420
rect 336752 306338 336780 310420
rect 336832 306400 336884 306406
rect 336936 306377 336964 310420
rect 337120 307018 337148 310420
rect 337108 307012 337160 307018
rect 337108 306954 337160 306960
rect 337200 306808 337252 306814
rect 337200 306750 337252 306756
rect 337016 306468 337068 306474
rect 337016 306410 337068 306416
rect 336832 306342 336884 306348
rect 336922 306368 336978 306377
rect 336740 306332 336792 306338
rect 336740 306274 336792 306280
rect 336740 306196 336792 306202
rect 336740 306138 336792 306144
rect 336016 292546 336596 292574
rect 336016 272542 336044 292546
rect 336004 272536 336056 272542
rect 336004 272478 336056 272484
rect 335912 268388 335964 268394
rect 335912 268330 335964 268336
rect 335820 260160 335872 260166
rect 335820 260102 335872 260108
rect 335728 257372 335780 257378
rect 335728 257314 335780 257320
rect 335636 253224 335688 253230
rect 335636 253166 335688 253172
rect 335544 251864 335596 251870
rect 335544 251806 335596 251812
rect 335452 249076 335504 249082
rect 335452 249018 335504 249024
rect 335360 246424 335412 246430
rect 335360 246366 335412 246372
rect 336752 245206 336780 306138
rect 336844 250510 336872 306342
rect 336922 306303 336978 306312
rect 336924 306264 336976 306270
rect 336924 306206 336976 306212
rect 336936 262886 336964 306206
rect 337028 282198 337056 306410
rect 337108 304156 337160 304162
rect 337108 304098 337160 304104
rect 337120 289134 337148 304098
rect 337212 293282 337240 306750
rect 337304 306474 337332 310420
rect 337292 306468 337344 306474
rect 337292 306410 337344 306416
rect 337292 306332 337344 306338
rect 337292 306274 337344 306280
rect 337304 297430 337332 306274
rect 337488 304162 337516 310420
rect 337672 306406 337700 310420
rect 337660 306400 337712 306406
rect 337660 306342 337712 306348
rect 337764 306270 337792 310420
rect 337752 306264 337804 306270
rect 337752 306206 337804 306212
rect 337948 306202 337976 310420
rect 338132 306202 338160 310420
rect 338316 309134 338344 310420
rect 338224 309106 338344 309134
rect 337936 306196 337988 306202
rect 337936 306138 337988 306144
rect 338120 306196 338172 306202
rect 338120 306138 338172 306144
rect 338224 306082 338252 309106
rect 338500 308281 338528 310420
rect 338684 309097 338712 310420
rect 338670 309088 338726 309097
rect 338670 309023 338726 309032
rect 338486 308272 338542 308281
rect 338486 308207 338542 308216
rect 338132 306054 338252 306082
rect 337476 304156 337528 304162
rect 337476 304098 337528 304104
rect 337292 297424 337344 297430
rect 337292 297366 337344 297372
rect 337200 293276 337252 293282
rect 337200 293218 337252 293224
rect 337108 289128 337160 289134
rect 337108 289070 337160 289076
rect 337016 282192 337068 282198
rect 337016 282134 337068 282140
rect 336924 262880 336976 262886
rect 336924 262822 336976 262828
rect 338132 260438 338160 306054
rect 338212 305992 338264 305998
rect 338212 305934 338264 305940
rect 338224 286482 338252 305934
rect 338868 303113 338896 310420
rect 338854 303104 338910 303113
rect 338854 303039 338910 303048
rect 339052 302954 339080 310420
rect 339236 308961 339264 310420
rect 339222 308952 339278 308961
rect 339222 308887 339278 308896
rect 339420 308582 339448 310420
rect 339408 308576 339460 308582
rect 339408 308518 339460 308524
rect 339604 306490 339632 310420
rect 339512 306462 339632 306490
rect 339512 303249 339540 306462
rect 339788 306320 339816 310420
rect 339972 307154 340000 310420
rect 339960 307148 340012 307154
rect 339960 307090 340012 307096
rect 340156 306377 340184 310420
rect 339604 306292 339816 306320
rect 340142 306368 340198 306377
rect 340142 306303 340198 306312
rect 339498 303240 339554 303249
rect 339498 303175 339554 303184
rect 338500 302926 339080 302954
rect 338500 302274 338528 302926
rect 338408 302246 338528 302274
rect 338408 297566 338436 302246
rect 338396 297560 338448 297566
rect 338396 297502 338448 297508
rect 339604 297498 339632 306292
rect 340248 302410 340276 310420
rect 339696 302382 340276 302410
rect 339696 300218 339724 302382
rect 339960 302320 340012 302326
rect 339960 302262 340012 302268
rect 339684 300212 339736 300218
rect 339684 300154 339736 300160
rect 339592 297492 339644 297498
rect 339592 297434 339644 297440
rect 338212 286476 338264 286482
rect 338212 286418 338264 286424
rect 339972 280974 340000 302262
rect 340432 301578 340460 310420
rect 340616 302326 340644 310420
rect 340800 306105 340828 310420
rect 340984 308378 341012 310420
rect 341168 309134 341196 310420
rect 341076 309106 341196 309134
rect 340972 308372 341024 308378
rect 340972 308314 341024 308320
rect 340972 306264 341024 306270
rect 340972 306206 341024 306212
rect 340786 306096 340842 306105
rect 340786 306031 340842 306040
rect 340604 302320 340656 302326
rect 340604 302262 340656 302268
rect 340420 301572 340472 301578
rect 340420 301514 340472 301520
rect 339960 280968 340012 280974
rect 339960 280910 340012 280916
rect 338120 260432 338172 260438
rect 338120 260374 338172 260380
rect 340984 253638 341012 306206
rect 341076 301510 341104 309106
rect 341156 306332 341208 306338
rect 341156 306274 341208 306280
rect 341064 301504 341116 301510
rect 341064 301446 341116 301452
rect 341168 300490 341196 306274
rect 341352 302234 341380 310420
rect 341536 305969 341564 310420
rect 341616 307828 341668 307834
rect 341616 307770 341668 307776
rect 341522 305960 341578 305969
rect 341522 305895 341578 305904
rect 341352 302206 341472 302234
rect 341156 300484 341208 300490
rect 341156 300426 341208 300432
rect 340972 253632 341024 253638
rect 340972 253574 341024 253580
rect 341444 252210 341472 302206
rect 341628 296714 341656 307770
rect 341720 306338 341748 310420
rect 341708 306332 341760 306338
rect 341708 306274 341760 306280
rect 341904 306270 341932 310420
rect 341892 306264 341944 306270
rect 341892 306206 341944 306212
rect 342088 305658 342116 310420
rect 342272 306354 342300 310420
rect 342456 307834 342484 310420
rect 342444 307828 342496 307834
rect 342444 307770 342496 307776
rect 342548 306490 342576 310420
rect 342548 306462 342668 306490
rect 342272 306326 342576 306354
rect 342352 306264 342404 306270
rect 342352 306206 342404 306212
rect 342076 305652 342128 305658
rect 342076 305594 342128 305600
rect 341536 296686 341656 296714
rect 341536 293418 341564 296686
rect 341524 293412 341576 293418
rect 341524 293354 341576 293360
rect 342364 282402 342392 306206
rect 342444 304496 342496 304502
rect 342444 304438 342496 304444
rect 342456 300558 342484 304438
rect 342444 300552 342496 300558
rect 342444 300494 342496 300500
rect 342548 300354 342576 306326
rect 342640 305794 342668 306462
rect 342628 305788 342680 305794
rect 342628 305730 342680 305736
rect 342732 304502 342760 310420
rect 342916 306270 342944 310420
rect 342904 306264 342956 306270
rect 342904 306206 342956 306212
rect 343100 305726 343128 310420
rect 343088 305720 343140 305726
rect 343088 305662 343140 305668
rect 342720 304496 342772 304502
rect 342720 304438 342772 304444
rect 343284 302234 343312 310420
rect 343364 308372 343416 308378
rect 343364 308314 343416 308320
rect 342640 302206 343312 302234
rect 342640 300626 342668 302206
rect 342628 300620 342680 300626
rect 342628 300562 342680 300568
rect 342536 300348 342588 300354
rect 342536 300290 342588 300296
rect 343376 300286 343404 308314
rect 343364 300280 343416 300286
rect 343364 300222 343416 300228
rect 343468 296714 343496 310420
rect 343652 306490 343680 310420
rect 343652 306462 343772 306490
rect 343640 306332 343692 306338
rect 343640 306274 343692 306280
rect 343652 300422 343680 306274
rect 343744 306241 343772 306462
rect 343730 306232 343786 306241
rect 343730 306167 343786 306176
rect 343836 302234 343864 310420
rect 344020 305930 344048 310420
rect 344204 306338 344232 310420
rect 344388 308378 344416 310420
rect 344376 308372 344428 308378
rect 344376 308314 344428 308320
rect 344192 306332 344244 306338
rect 344192 306274 344244 306280
rect 344008 305924 344060 305930
rect 344008 305866 344060 305872
rect 344572 305862 344600 310420
rect 344756 308650 344784 310420
rect 344744 308644 344796 308650
rect 344744 308586 344796 308592
rect 344560 305856 344612 305862
rect 344560 305798 344612 305804
rect 344940 303521 344968 310420
rect 345032 308922 345060 310420
rect 345020 308916 345072 308922
rect 345020 308858 345072 308864
rect 344926 303512 344982 303521
rect 344926 303447 344982 303456
rect 345216 303385 345244 310420
rect 345400 308854 345428 310420
rect 345388 308848 345440 308854
rect 345388 308790 345440 308796
rect 345202 303376 345258 303385
rect 345202 303311 345258 303320
rect 345584 302938 345612 310420
rect 345768 307970 345796 310420
rect 345756 307964 345808 307970
rect 345756 307906 345808 307912
rect 345952 303006 345980 310420
rect 346136 308786 346164 310420
rect 346124 308780 346176 308786
rect 346124 308722 346176 308728
rect 346320 303074 346348 310420
rect 346504 308990 346532 310420
rect 346492 308984 346544 308990
rect 346492 308926 346544 308932
rect 346688 303346 346716 310420
rect 346872 309058 346900 310420
rect 346860 309052 346912 309058
rect 346860 308994 346912 309000
rect 346676 303340 346728 303346
rect 346676 303282 346728 303288
rect 347056 303142 347084 310420
rect 347240 309126 347268 310420
rect 347228 309120 347280 309126
rect 347228 309062 347280 309068
rect 347136 308508 347188 308514
rect 347136 308450 347188 308456
rect 347044 303136 347096 303142
rect 347044 303078 347096 303084
rect 346308 303068 346360 303074
rect 346308 303010 346360 303016
rect 345940 303000 345992 303006
rect 345940 302942 345992 302948
rect 345572 302932 345624 302938
rect 345572 302874 345624 302880
rect 343744 302206 343864 302234
rect 343744 300830 343772 302206
rect 343732 300824 343784 300830
rect 343732 300766 343784 300772
rect 343640 300416 343692 300422
rect 343640 300358 343692 300364
rect 342916 296686 343496 296714
rect 342352 282396 342404 282402
rect 342352 282338 342404 282344
rect 342916 256358 342944 296686
rect 342904 256352 342956 256358
rect 342904 256294 342956 256300
rect 341432 252204 341484 252210
rect 341432 252146 341484 252152
rect 336832 250504 336884 250510
rect 336832 250446 336884 250452
rect 347148 247518 347176 308450
rect 347332 303210 347360 310420
rect 347516 307902 347544 310420
rect 347504 307896 347556 307902
rect 347504 307838 347556 307844
rect 347700 303414 347728 310420
rect 347884 308106 347912 310420
rect 347872 308100 347924 308106
rect 347872 308042 347924 308048
rect 347688 303408 347740 303414
rect 347688 303350 347740 303356
rect 347320 303204 347372 303210
rect 347320 303146 347372 303152
rect 348068 302734 348096 310420
rect 348252 308718 348280 310420
rect 348240 308712 348292 308718
rect 348240 308654 348292 308660
rect 348436 303482 348464 310420
rect 348620 305998 348648 310420
rect 348608 305992 348660 305998
rect 348608 305934 348660 305940
rect 348424 303476 348476 303482
rect 348424 303418 348476 303424
rect 348804 302870 348832 310420
rect 348988 306134 349016 310420
rect 349172 306490 349200 310420
rect 349172 306462 349292 306490
rect 349160 306264 349212 306270
rect 349160 306206 349212 306212
rect 348976 306128 349028 306134
rect 348976 306070 349028 306076
rect 348792 302864 348844 302870
rect 348792 302806 348844 302812
rect 348056 302728 348108 302734
rect 348056 302670 348108 302676
rect 349172 300694 349200 306206
rect 349264 303618 349292 306462
rect 349356 306066 349384 310420
rect 349344 306060 349396 306066
rect 349344 306002 349396 306008
rect 349252 303612 349304 303618
rect 349252 303554 349304 303560
rect 349540 303278 349568 310420
rect 349724 306474 349752 310420
rect 349712 306468 349764 306474
rect 349712 306410 349764 306416
rect 349816 303550 349844 310420
rect 349896 308440 349948 308446
rect 349896 308382 349948 308388
rect 349804 303544 349856 303550
rect 349804 303486 349856 303492
rect 349528 303272 349580 303278
rect 349528 303214 349580 303220
rect 349160 300688 349212 300694
rect 349160 300630 349212 300636
rect 347136 247512 347188 247518
rect 347136 247454 347188 247460
rect 349908 245206 349936 308382
rect 350000 306202 350028 310420
rect 350184 306270 350212 310420
rect 350368 306270 350396 310420
rect 350552 308394 350580 310420
rect 350736 308514 350764 310420
rect 350724 308508 350776 308514
rect 350724 308450 350776 308456
rect 350552 308366 350856 308394
rect 350540 308304 350592 308310
rect 350540 308246 350592 308252
rect 350172 306264 350224 306270
rect 350172 306206 350224 306212
rect 350356 306264 350408 306270
rect 350356 306206 350408 306212
rect 349988 306196 350040 306202
rect 349988 306138 350040 306144
rect 350552 300762 350580 308246
rect 350724 308236 350776 308242
rect 350724 308178 350776 308184
rect 350632 307148 350684 307154
rect 350632 307090 350684 307096
rect 350540 300756 350592 300762
rect 350540 300698 350592 300704
rect 350644 300082 350672 307090
rect 350632 300076 350684 300082
rect 350632 300018 350684 300024
rect 350736 300014 350764 308178
rect 350724 300008 350776 300014
rect 350724 299950 350776 299956
rect 350828 299946 350856 308366
rect 350920 308310 350948 310420
rect 351104 308394 351132 310420
rect 351012 308366 351132 308394
rect 350908 308304 350960 308310
rect 350908 308246 350960 308252
rect 350908 308168 350960 308174
rect 350908 308110 350960 308116
rect 350920 305590 350948 308110
rect 350908 305584 350960 305590
rect 350908 305526 350960 305532
rect 351012 305522 351040 308366
rect 351288 308242 351316 310420
rect 351276 308236 351328 308242
rect 351276 308178 351328 308184
rect 351000 305516 351052 305522
rect 351000 305458 351052 305464
rect 351472 305454 351500 310420
rect 351656 307154 351684 310420
rect 351840 308174 351868 310420
rect 351828 308168 351880 308174
rect 351828 308110 351880 308116
rect 351644 307148 351696 307154
rect 351644 307090 351696 307096
rect 351460 305448 351512 305454
rect 351460 305390 351512 305396
rect 352024 302802 352052 310420
rect 352472 308712 352524 308718
rect 352472 308654 352524 308660
rect 352484 308514 352512 308654
rect 352472 308508 352524 308514
rect 352472 308450 352524 308456
rect 352012 302796 352064 302802
rect 352012 302738 352064 302744
rect 350816 299940 350868 299946
rect 350816 299882 350868 299888
rect 352576 246362 352604 434454
rect 352840 432268 352892 432274
rect 352840 432210 352892 432216
rect 352748 432200 352800 432206
rect 352748 432142 352800 432148
rect 352656 432064 352708 432070
rect 352656 432006 352708 432012
rect 352668 299470 352696 432006
rect 352760 353258 352788 432142
rect 352852 405686 352880 432210
rect 352840 405680 352892 405686
rect 352840 405622 352892 405628
rect 352748 353252 352800 353258
rect 352748 353194 352800 353200
rect 352748 308712 352800 308718
rect 352748 308654 352800 308660
rect 352760 307970 352788 308654
rect 352748 307964 352800 307970
rect 352748 307906 352800 307912
rect 352656 299464 352708 299470
rect 352656 299406 352708 299412
rect 353956 259418 353984 436358
rect 355324 436348 355376 436354
rect 355324 436290 355376 436296
rect 355336 273222 355364 436290
rect 356704 435056 356756 435062
rect 356704 434998 356756 435004
rect 355416 430636 355468 430642
rect 355416 430578 355468 430584
rect 355428 419490 355456 430578
rect 355416 419484 355468 419490
rect 355416 419426 355468 419432
rect 356716 325650 356744 434998
rect 580908 434920 580960 434926
rect 580908 434862 580960 434868
rect 580540 434852 580592 434858
rect 580540 434794 580592 434800
rect 577504 434784 577556 434790
rect 577504 434726 577556 434732
rect 357898 433800 357954 433809
rect 357898 433735 357954 433744
rect 356704 325644 356756 325650
rect 356704 325586 356756 325592
rect 356796 309596 356848 309602
rect 356796 309538 356848 309544
rect 356704 309460 356756 309466
rect 356704 309402 356756 309408
rect 355414 308680 355470 308689
rect 355414 308615 355470 308624
rect 355324 273216 355376 273222
rect 355324 273158 355376 273164
rect 353944 259412 353996 259418
rect 353944 259354 353996 259360
rect 352564 246356 352616 246362
rect 352564 246298 352616 246304
rect 336740 245200 336792 245206
rect 336740 245142 336792 245148
rect 349896 245200 349948 245206
rect 349896 245142 349948 245148
rect 314660 244870 314712 244876
rect 332598 244896 332654 244905
rect 332598 244831 332654 244840
rect 302332 244792 302384 244798
rect 302332 244734 302384 244740
rect 355428 244526 355456 308615
rect 355416 244520 355468 244526
rect 355416 244462 355468 244468
rect 295708 243772 295760 243778
rect 295708 243714 295760 243720
rect 295616 243704 295668 243710
rect 295616 243646 295668 243652
rect 295524 243636 295576 243642
rect 295524 243578 295576 243584
rect 295340 243510 295392 243516
rect 295430 243536 295486 243545
rect 295430 243471 295486 243480
rect 256700 159928 256752 159934
rect 238206 159896 238262 159905
rect 238206 159831 238262 159840
rect 239586 159896 239642 159905
rect 239586 159831 239642 159840
rect 241702 159896 241758 159905
rect 256700 159870 256752 159876
rect 273626 159896 273682 159905
rect 241702 159831 241758 159840
rect 238220 158982 238248 159831
rect 238208 158976 238260 158982
rect 238208 158918 238260 158924
rect 239600 158914 239628 159831
rect 239588 158908 239640 158914
rect 239588 158850 239640 158856
rect 241716 158846 241744 159831
rect 255962 159624 256018 159633
rect 255962 159559 256018 159568
rect 241704 158840 241756 158846
rect 241704 158782 241756 158788
rect 240508 158772 240560 158778
rect 240508 158714 240560 158720
rect 234620 158704 234672 158710
rect 220818 158672 220874 158681
rect 240520 158681 240548 158714
rect 248328 158704 248380 158710
rect 234620 158646 234672 158652
rect 240506 158672 240562 158681
rect 220818 158607 220874 158616
rect 233240 158636 233292 158642
rect 219438 157856 219494 157865
rect 219438 157791 219494 157800
rect 219452 16574 219480 157791
rect 220832 16574 220860 158607
rect 233240 158578 233292 158584
rect 224958 158536 225014 158545
rect 224958 158471 225014 158480
rect 223578 158400 223634 158409
rect 223578 158335 223634 158344
rect 219452 16546 220032 16574
rect 220832 16546 221136 16574
rect 219348 4072 219400 4078
rect 219348 4014 219400 4020
rect 219254 3768 219310 3777
rect 219310 3726 219388 3754
rect 219254 3703 219310 3712
rect 219360 3641 219388 3726
rect 219346 3632 219402 3641
rect 219346 3567 219402 3576
rect 219254 3496 219310 3505
rect 219164 3460 219216 3466
rect 219254 3431 219310 3440
rect 219164 3402 219216 3408
rect 219268 480 219296 3431
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 16546
rect 222750 3904 222806 3913
rect 222750 3839 222806 3848
rect 222764 480 222792 3839
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 158335
rect 224972 16574 225000 158471
rect 231858 158264 231914 158273
rect 231858 158199 231914 158208
rect 230480 157956 230532 157962
rect 230480 157898 230532 157904
rect 229100 157888 229152 157894
rect 229100 157830 229152 157836
rect 227720 157820 227772 157826
rect 227720 157762 227772 157768
rect 227732 16574 227760 157762
rect 229112 16574 229140 157830
rect 230492 16574 230520 157898
rect 224972 16546 225184 16574
rect 227732 16546 228312 16574
rect 229112 16546 229416 16574
rect 230492 16546 231072 16574
rect 225156 480 225184 16546
rect 226338 3632 226394 3641
rect 226338 3567 226394 3576
rect 226352 480 226380 3567
rect 227534 3224 227590 3233
rect 227534 3159 227590 3168
rect 227548 480 227576 3159
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 16546
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 16546
rect 231044 480 231072 16546
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 231872 354 231900 158199
rect 233252 16574 233280 158578
rect 233252 16546 233464 16574
rect 233436 480 233464 16546
rect 234632 11762 234660 158646
rect 240506 158607 240562 158616
rect 248326 158672 248328 158681
rect 248380 158672 248382 158681
rect 248326 158607 248382 158616
rect 250166 158672 250222 158681
rect 250166 158607 250222 158616
rect 251454 158672 251510 158681
rect 251454 158607 251510 158616
rect 254582 158672 254638 158681
rect 254582 158607 254638 158616
rect 236000 158568 236052 158574
rect 236000 158510 236052 158516
rect 234712 158500 234764 158506
rect 234712 158442 234764 158448
rect 234620 11756 234672 11762
rect 234620 11698 234672 11704
rect 234724 6914 234752 158442
rect 236012 16574 236040 158510
rect 242992 158432 243044 158438
rect 242992 158374 243044 158380
rect 242900 158364 242952 158370
rect 242900 158306 242952 158312
rect 238758 158128 238814 158137
rect 238758 158063 238814 158072
rect 237380 155780 237432 155786
rect 237380 155722 237432 155728
rect 237392 16574 237420 155722
rect 238772 16574 238800 158063
rect 241520 155712 241572 155718
rect 241520 155654 241572 155660
rect 241532 16574 241560 155654
rect 236012 16546 236592 16574
rect 237392 16546 237696 16574
rect 238772 16546 239352 16574
rect 241532 16546 241744 16574
rect 235816 11756 235868 11762
rect 235816 11698 235868 11704
rect 234632 6886 234752 6914
rect 234632 480 234660 6886
rect 235828 480 235856 11698
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 16546
rect 239324 480 239352 16546
rect 240506 3360 240562 3369
rect 240506 3295 240562 3304
rect 240520 480 240548 3295
rect 241716 480 241744 16546
rect 242912 11762 242940 158306
rect 242900 11756 242952 11762
rect 242900 11698 242952 11704
rect 243004 6914 243032 158374
rect 245660 158296 245712 158302
rect 245660 158238 245712 158244
rect 245672 16574 245700 158238
rect 247040 158228 247092 158234
rect 247040 158170 247092 158176
rect 247052 16574 247080 158170
rect 249800 158160 249852 158166
rect 249800 158102 249852 158108
rect 248420 155644 248472 155650
rect 248420 155586 248472 155592
rect 245672 16546 245976 16574
rect 247052 16546 247632 16574
rect 244096 11756 244148 11762
rect 244096 11698 244148 11704
rect 242912 6886 243032 6914
rect 242912 480 242940 6886
rect 244108 480 244136 11698
rect 245200 3256 245252 3262
rect 245200 3198 245252 3204
rect 245212 480 245240 3198
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 16546
rect 247604 480 247632 16546
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248432 354 248460 155586
rect 249812 16574 249840 158102
rect 250180 157350 250208 158607
rect 251086 158128 251142 158137
rect 251086 158063 251142 158072
rect 250168 157344 250220 157350
rect 250168 157286 250220 157292
rect 251100 155854 251128 158063
rect 251178 157992 251234 158001
rect 251178 157927 251234 157936
rect 251088 155848 251140 155854
rect 251088 155790 251140 155796
rect 249812 16546 250024 16574
rect 249996 480 250024 16546
rect 251192 480 251220 157927
rect 251468 157282 251496 158607
rect 254596 158370 254624 158607
rect 255976 158506 256004 159559
rect 256054 158672 256110 158681
rect 256054 158607 256056 158616
rect 256108 158607 256110 158616
rect 256056 158578 256108 158584
rect 255964 158500 256016 158506
rect 255964 158442 256016 158448
rect 254584 158364 254636 158370
rect 254584 158306 254636 158312
rect 252560 158092 252612 158098
rect 252560 158034 252612 158040
rect 252374 157992 252430 158001
rect 252374 157927 252430 157936
rect 251456 157276 251508 157282
rect 251456 157218 251508 157224
rect 252388 155922 252416 157927
rect 252376 155916 252428 155922
rect 252376 155858 252428 155864
rect 251270 155272 251326 155281
rect 251270 155207 251326 155216
rect 251284 16574 251312 155207
rect 252572 16574 252600 158034
rect 253570 157992 253626 158001
rect 253570 157927 253626 157936
rect 253584 155786 253612 157927
rect 253662 157448 253718 157457
rect 253662 157383 253718 157392
rect 253572 155780 253624 155786
rect 253572 155722 253624 155728
rect 253676 154562 253704 157383
rect 255320 155576 255372 155582
rect 255320 155518 255372 155524
rect 253664 154556 253716 154562
rect 253664 154498 253716 154504
rect 255332 16574 255360 155518
rect 251284 16546 252416 16574
rect 252572 16546 253520 16574
rect 255332 16546 255912 16574
rect 252388 480 252416 16546
rect 253492 480 253520 16546
rect 254676 3324 254728 3330
rect 254676 3266 254728 3272
rect 254688 480 254716 3266
rect 255884 480 255912 16546
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 256712 354 256740 159870
rect 264980 159860 265032 159866
rect 273626 159831 273682 159840
rect 276110 159896 276166 159905
rect 276110 159831 276166 159840
rect 278502 159896 278558 159905
rect 278502 159831 278558 159840
rect 293498 159896 293554 159905
rect 293498 159831 293554 159840
rect 295890 159896 295946 159905
rect 295890 159831 295946 159840
rect 303526 159896 303582 159905
rect 303526 159831 303582 159840
rect 310978 159896 311034 159905
rect 310978 159831 311034 159840
rect 313462 159896 313518 159905
rect 313462 159831 313518 159840
rect 264980 159802 265032 159808
rect 263600 159792 263652 159798
rect 263600 159734 263652 159740
rect 260840 159724 260892 159730
rect 260840 159666 260892 159672
rect 259552 158772 259604 158778
rect 259552 158714 259604 158720
rect 259564 158681 259592 158714
rect 257158 158672 257214 158681
rect 257158 158607 257214 158616
rect 258262 158672 258318 158681
rect 258262 158607 258318 158616
rect 258630 158672 258686 158681
rect 258630 158607 258686 158616
rect 259550 158672 259606 158681
rect 259550 158607 259606 158616
rect 257172 158438 257200 158607
rect 257160 158432 257212 158438
rect 257160 158374 257212 158380
rect 258276 158302 258304 158607
rect 258264 158296 258316 158302
rect 258264 158238 258316 158244
rect 258644 154494 258672 158607
rect 259552 155508 259604 155514
rect 259552 155450 259604 155456
rect 258632 154488 258684 154494
rect 258632 154430 258684 154436
rect 259564 6914 259592 155450
rect 260852 16574 260880 159666
rect 262864 158840 262916 158846
rect 262864 158782 262916 158788
rect 262876 158681 262904 158782
rect 261206 158672 261262 158681
rect 261206 158607 261262 158616
rect 262862 158672 262918 158681
rect 262862 158607 262918 158616
rect 261220 158574 261248 158607
rect 261208 158568 261260 158574
rect 261208 158510 261260 158516
rect 263612 16574 263640 159734
rect 263968 158908 264020 158914
rect 263968 158850 264020 158856
rect 263980 158681 264008 158850
rect 263966 158672 264022 158681
rect 263966 158607 264022 158616
rect 263966 157448 264022 157457
rect 263966 157383 264022 157392
rect 263980 154426 264008 157383
rect 263968 154420 264020 154426
rect 263968 154362 264020 154368
rect 260852 16546 261800 16574
rect 263612 16546 264192 16574
rect 259472 6886 259592 6914
rect 258264 3392 258316 3398
rect 258264 3334 258316 3340
rect 258276 480 258304 3334
rect 259472 480 259500 6886
rect 260656 4140 260708 4146
rect 260656 4082 260708 4088
rect 260668 480 260696 4082
rect 261772 480 261800 16546
rect 262956 3936 263008 3942
rect 262956 3878 263008 3884
rect 262968 480 262996 3878
rect 264164 480 264192 16546
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 264992 354 265020 159802
rect 269120 159656 269172 159662
rect 265346 159624 265402 159633
rect 269120 159598 269172 159604
rect 271050 159624 271106 159633
rect 265346 159559 265402 159568
rect 265360 158982 265388 159559
rect 265348 158976 265400 158982
rect 265348 158918 265400 158924
rect 265990 158672 266046 158681
rect 265990 158607 266046 158616
rect 266818 158672 266874 158681
rect 266818 158607 266874 158616
rect 267646 158672 267702 158681
rect 267646 158607 267702 158616
rect 268750 158672 268806 158681
rect 268750 158607 268806 158616
rect 266004 158234 266032 158607
rect 265992 158228 266044 158234
rect 265992 158170 266044 158176
rect 266832 157010 266860 158607
rect 267660 157214 267688 158607
rect 267648 157208 267700 157214
rect 267648 157150 267700 157156
rect 268764 157146 268792 158607
rect 268934 157992 268990 158001
rect 268934 157927 268990 157936
rect 268752 157140 268804 157146
rect 268752 157082 268804 157088
rect 266820 157004 266872 157010
rect 266820 156946 266872 156952
rect 268948 155718 268976 157927
rect 268936 155712 268988 155718
rect 268936 155654 268988 155660
rect 269132 16574 269160 159598
rect 271050 159559 271106 159568
rect 269854 158672 269910 158681
rect 269854 158607 269910 158616
rect 269868 156942 269896 158607
rect 269856 156936 269908 156942
rect 269856 156878 269908 156884
rect 271064 154358 271092 159559
rect 273640 159050 273668 159831
rect 276020 159520 276072 159526
rect 276020 159462 276072 159468
rect 273628 159044 273680 159050
rect 273628 158986 273680 158992
rect 271142 158672 271198 158681
rect 271142 158607 271198 158616
rect 272246 158672 272302 158681
rect 272246 158607 272302 158616
rect 274178 158672 274234 158681
rect 274178 158607 274234 158616
rect 274454 158672 274510 158681
rect 274454 158607 274510 158616
rect 275926 158672 275982 158681
rect 275926 158607 275982 158616
rect 271156 157078 271184 158607
rect 271144 157072 271196 157078
rect 271144 157014 271196 157020
rect 272260 156874 272288 158607
rect 273260 158024 273312 158030
rect 273260 157966 273312 157972
rect 272248 156868 272300 156874
rect 272248 156810 272300 156816
rect 271052 154352 271104 154358
rect 271052 154294 271104 154300
rect 269132 16546 270080 16574
rect 266544 4072 266596 4078
rect 266544 4014 266596 4020
rect 266556 480 266584 4014
rect 267740 4004 267792 4010
rect 267740 3946 267792 3952
rect 267752 480 267780 3946
rect 268844 3868 268896 3874
rect 268844 3810 268896 3816
rect 268856 480 268884 3810
rect 270052 480 270080 16546
rect 271236 3800 271288 3806
rect 271236 3742 271288 3748
rect 271248 480 271276 3742
rect 272432 3664 272484 3670
rect 272432 3606 272484 3612
rect 272444 480 272472 3606
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273272 354 273300 157966
rect 274192 156806 274220 158607
rect 274180 156800 274232 156806
rect 274180 156742 274232 156748
rect 274468 156738 274496 158607
rect 274456 156732 274508 156738
rect 274456 156674 274508 156680
rect 275940 156670 275968 158607
rect 275928 156664 275980 156670
rect 275928 156606 275980 156612
rect 274824 3596 274876 3602
rect 274824 3538 274876 3544
rect 274836 480 274864 3538
rect 276032 480 276060 159462
rect 276124 159186 276152 159831
rect 276204 159588 276256 159594
rect 276204 159530 276256 159536
rect 276112 159180 276164 159186
rect 276112 159122 276164 159128
rect 276216 142154 276244 159530
rect 278516 159118 278544 159831
rect 278780 159452 278832 159458
rect 278780 159394 278832 159400
rect 278504 159112 278556 159118
rect 278504 159054 278556 159060
rect 277122 158128 277178 158137
rect 277122 158063 277178 158072
rect 278134 158128 278190 158137
rect 278134 158063 278190 158072
rect 277136 156602 277164 158063
rect 277124 156596 277176 156602
rect 277124 156538 277176 156544
rect 278148 156466 278176 158063
rect 278136 156460 278188 156466
rect 278136 156402 278188 156408
rect 276124 142126 276244 142154
rect 276124 16574 276152 142126
rect 278792 16574 278820 159394
rect 282920 159384 282972 159390
rect 282920 159326 282972 159332
rect 281078 158672 281134 158681
rect 281078 158607 281134 158616
rect 279974 158128 280030 158137
rect 279974 158063 280030 158072
rect 279988 156534 280016 158063
rect 279976 156528 280028 156534
rect 279976 156470 280028 156476
rect 281092 155650 281120 158607
rect 281080 155644 281132 155650
rect 281080 155586 281132 155592
rect 280160 155440 280212 155446
rect 280160 155382 280212 155388
rect 280172 16574 280200 155382
rect 282932 16574 282960 159326
rect 293512 159254 293540 159831
rect 295904 159322 295932 159831
rect 298466 159760 298522 159769
rect 298466 159695 298522 159704
rect 298480 159526 298508 159695
rect 298468 159520 298520 159526
rect 298468 159462 298520 159468
rect 303540 159390 303568 159831
rect 310992 159458 311020 159831
rect 313476 159594 313504 159831
rect 313464 159588 313516 159594
rect 313464 159530 313516 159536
rect 310980 159452 311032 159458
rect 310980 159394 311032 159400
rect 303528 159384 303580 159390
rect 303528 159326 303580 159332
rect 295892 159316 295944 159322
rect 295892 159258 295944 159264
rect 293500 159248 293552 159254
rect 293500 159190 293552 159196
rect 291014 158672 291070 158681
rect 291014 158607 291070 158616
rect 300950 158672 301006 158681
rect 300950 158607 301006 158616
rect 308678 158672 308734 158681
rect 308678 158607 308734 158616
rect 321098 158672 321154 158681
rect 321098 158607 321154 158616
rect 323398 158672 323454 158681
rect 323398 158607 323454 158616
rect 325974 158672 326030 158681
rect 325974 158607 326030 158616
rect 291028 158166 291056 158607
rect 291016 158160 291068 158166
rect 291016 158102 291068 158108
rect 300964 158098 300992 158607
rect 300952 158092 301004 158098
rect 300952 158034 301004 158040
rect 308692 158030 308720 158607
rect 308680 158024 308732 158030
rect 308680 157966 308732 157972
rect 321112 157962 321140 158607
rect 321100 157956 321152 157962
rect 321100 157898 321152 157904
rect 323412 157894 323440 158607
rect 323400 157888 323452 157894
rect 283746 157856 283802 157865
rect 283746 157791 283802 157800
rect 286506 157856 286562 157865
rect 323400 157830 323452 157836
rect 325988 157826 326016 158607
rect 353942 158128 353998 158137
rect 353942 158063 353998 158072
rect 286506 157791 286562 157800
rect 325976 157820 326028 157826
rect 283760 155582 283788 157791
rect 283748 155576 283800 155582
rect 283748 155518 283800 155524
rect 286520 155514 286548 157791
rect 325976 157762 326028 157768
rect 288254 157448 288310 157457
rect 288254 157383 288310 157392
rect 306102 157448 306158 157457
rect 306102 157383 306158 157392
rect 315854 157448 315910 157457
rect 315854 157383 315910 157392
rect 318614 157448 318670 157457
rect 318614 157383 318670 157392
rect 286508 155508 286560 155514
rect 286508 155450 286560 155456
rect 284392 155372 284444 155378
rect 284392 155314 284444 155320
rect 284300 155236 284352 155242
rect 284300 155178 284352 155184
rect 276124 16546 276704 16574
rect 278792 16546 279096 16574
rect 280172 16546 280752 16574
rect 282932 16546 283144 16574
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276676 354 276704 16546
rect 278320 3732 278372 3738
rect 278320 3674 278372 3680
rect 278332 480 278360 3674
rect 277094 354 277206 480
rect 276676 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 280724 480 280752 16546
rect 281908 3528 281960 3534
rect 281908 3470 281960 3476
rect 281920 480 281948 3470
rect 283116 480 283144 16546
rect 284312 480 284340 155178
rect 284404 16574 284432 155314
rect 285680 155304 285732 155310
rect 285680 155246 285732 155252
rect 285692 16574 285720 155246
rect 288268 154290 288296 157383
rect 292580 155372 292632 155378
rect 292580 155314 292632 155320
rect 289820 155236 289872 155242
rect 289820 155178 289872 155184
rect 288256 154284 288308 154290
rect 288256 154226 288308 154232
rect 284404 16546 284984 16574
rect 285692 16546 286640 16574
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 284956 354 284984 16546
rect 286612 480 286640 16546
rect 287796 3460 287848 3466
rect 287796 3402 287848 3408
rect 288992 3460 289044 3466
rect 288992 3402 289044 3408
rect 287808 480 287836 3402
rect 289004 480 289032 3402
rect 285374 354 285486 480
rect 284956 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 289832 354 289860 155178
rect 291384 3664 291436 3670
rect 291384 3606 291436 3612
rect 291396 480 291424 3606
rect 292592 3602 292620 155314
rect 292672 155304 292724 155310
rect 292672 155246 292724 155252
rect 292580 3596 292632 3602
rect 292580 3538 292632 3544
rect 292684 3482 292712 155246
rect 306116 154222 306144 157383
rect 306104 154216 306156 154222
rect 306104 154158 306156 154164
rect 315868 154154 315896 157383
rect 315856 154148 315908 154154
rect 315856 154090 315908 154096
rect 318628 154086 318656 157383
rect 348516 155440 348568 155446
rect 348516 155382 348568 155388
rect 348424 155168 348476 155174
rect 348424 155110 348476 155116
rect 318616 154080 318668 154086
rect 318616 154022 318668 154028
rect 316224 9376 316276 9382
rect 316224 9318 316276 9324
rect 312636 9308 312688 9314
rect 312636 9250 312688 9256
rect 298468 9240 298520 9246
rect 298468 9182 298520 9188
rect 297272 8968 297324 8974
rect 297272 8910 297324 8916
rect 294880 3732 294932 3738
rect 294880 3674 294932 3680
rect 293316 3596 293368 3602
rect 293316 3538 293368 3544
rect 292592 3454 292712 3482
rect 292592 480 292620 3454
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293328 354 293356 3538
rect 294892 480 294920 3674
rect 296076 3596 296128 3602
rect 296076 3538 296128 3544
rect 296088 480 296116 3538
rect 297284 480 297312 8910
rect 298480 480 298508 9182
rect 301964 9172 302016 9178
rect 301964 9114 302016 9120
rect 300768 9104 300820 9110
rect 300768 9046 300820 9052
rect 299664 3528 299716 3534
rect 299664 3470 299716 3476
rect 299676 480 299704 3470
rect 300780 480 300808 9046
rect 301976 480 302004 9114
rect 304356 9036 304408 9042
rect 304356 8978 304408 8984
rect 303160 6180 303212 6186
rect 303160 6122 303212 6128
rect 303172 480 303200 6122
rect 304368 480 304396 8978
rect 305550 8936 305606 8945
rect 305550 8871 305606 8880
rect 305564 480 305592 8871
rect 310244 6452 310296 6458
rect 310244 6394 310296 6400
rect 307944 6316 307996 6322
rect 307944 6258 307996 6264
rect 306748 6248 306800 6254
rect 306748 6190 306800 6196
rect 306760 480 306788 6190
rect 307956 480 307984 6258
rect 309048 3800 309100 3806
rect 309048 3742 309100 3748
rect 309060 480 309088 3742
rect 310256 480 310284 6394
rect 311440 6384 311492 6390
rect 311440 6326 311492 6332
rect 311452 480 311480 6326
rect 312648 480 312676 9250
rect 315028 6656 315080 6662
rect 315028 6598 315080 6604
rect 313832 6588 313884 6594
rect 313832 6530 313884 6536
rect 313844 480 313872 6530
rect 315040 480 315068 6598
rect 316236 480 316264 9318
rect 319718 9072 319774 9081
rect 319718 9007 319774 9016
rect 317328 6860 317380 6866
rect 317328 6802 317380 6808
rect 317340 480 317368 6802
rect 318524 6520 318576 6526
rect 318524 6462 318576 6468
rect 318536 480 318564 6462
rect 319732 480 319760 9007
rect 322112 6792 322164 6798
rect 322112 6734 322164 6740
rect 348054 6760 348110 6769
rect 320916 6724 320968 6730
rect 320916 6666 320968 6672
rect 320928 480 320956 6666
rect 322124 480 322152 6734
rect 348054 6695 348110 6704
rect 344558 6624 344614 6633
rect 344558 6559 344614 6568
rect 340970 6488 341026 6497
rect 340970 6423 341026 6432
rect 337474 6352 337530 6361
rect 337474 6287 337530 6296
rect 333886 6216 333942 6225
rect 333886 6151 333942 6160
rect 326804 6112 326856 6118
rect 326804 6054 326856 6060
rect 323308 6044 323360 6050
rect 323308 5986 323360 5992
rect 323320 480 323348 5986
rect 324412 4004 324464 4010
rect 324412 3946 324464 3952
rect 324424 480 324452 3946
rect 325608 3868 325660 3874
rect 325608 3810 325660 3816
rect 325620 480 325648 3810
rect 326816 480 326844 6054
rect 330392 5976 330444 5982
rect 330392 5918 330444 5924
rect 328000 4072 328052 4078
rect 328000 4014 328052 4020
rect 328012 480 328040 4014
rect 329196 3936 329248 3942
rect 329196 3878 329248 3884
rect 329208 480 329236 3878
rect 330404 480 330432 5918
rect 332692 4140 332744 4146
rect 332692 4082 332744 4088
rect 331588 3392 331640 3398
rect 331588 3334 331640 3340
rect 331600 480 331628 3334
rect 332704 480 332732 4082
rect 333900 480 333928 6151
rect 336280 3324 336332 3330
rect 336280 3266 336332 3272
rect 335084 3256 335136 3262
rect 335084 3198 335136 3204
rect 335096 480 335124 3198
rect 336292 480 336320 3266
rect 337488 480 337516 6287
rect 338670 3496 338726 3505
rect 338670 3431 338726 3440
rect 338684 480 338712 3431
rect 339866 3360 339922 3369
rect 339866 3295 339922 3304
rect 339880 480 339908 3295
rect 340984 480 341012 6423
rect 342166 3768 342222 3777
rect 342166 3703 342222 3712
rect 342180 480 342208 3703
rect 343362 3632 343418 3641
rect 343362 3567 343418 3576
rect 343376 480 343404 3567
rect 344572 480 344600 6559
rect 346950 4040 347006 4049
rect 346950 3975 347006 3984
rect 345754 3904 345810 3913
rect 345754 3839 345810 3848
rect 345768 480 345796 3839
rect 346964 480 346992 3975
rect 348068 480 348096 6695
rect 348436 3670 348464 155110
rect 348528 3738 348556 155382
rect 351642 6896 351698 6905
rect 351642 6831 351698 6840
rect 348516 3732 348568 3738
rect 348516 3674 348568 3680
rect 349252 3732 349304 3738
rect 349252 3674 349304 3680
rect 348424 3664 348476 3670
rect 348424 3606 348476 3612
rect 349264 480 349292 3674
rect 350448 3664 350500 3670
rect 350448 3606 350500 3612
rect 350460 480 350488 3606
rect 351656 480 351684 6831
rect 353956 3602 353984 158063
rect 354126 157992 354182 158001
rect 354126 157927 354182 157936
rect 353944 3596 353996 3602
rect 353944 3538 353996 3544
rect 354140 3466 354168 157927
rect 356716 3806 356744 309402
rect 356808 6322 356836 309538
rect 357530 308544 357586 308553
rect 357530 308479 357586 308488
rect 357440 279744 357492 279750
rect 357440 279686 357492 279692
rect 356796 6316 356848 6322
rect 356796 6258 356848 6264
rect 356704 3800 356756 3806
rect 356704 3742 356756 3748
rect 357348 3800 357400 3806
rect 357348 3742 357400 3748
rect 356702 3632 356758 3641
rect 356702 3567 356758 3576
rect 354128 3460 354180 3466
rect 354128 3402 354180 3408
rect 356336 3460 356388 3466
rect 356336 3402 356388 3408
rect 356152 3324 356204 3330
rect 356152 3266 356204 3272
rect 352838 3224 352894 3233
rect 352838 3159 352894 3168
rect 354036 3188 354088 3194
rect 352852 480 352880 3159
rect 354036 3130 354088 3136
rect 354048 480 354076 3130
rect 356164 3126 356192 3266
rect 356152 3120 356204 3126
rect 356152 3062 356204 3068
rect 355232 3052 355284 3058
rect 355232 2994 355284 3000
rect 355244 480 355272 2994
rect 356348 480 356376 3402
rect 356716 3097 356744 3567
rect 357360 3534 357388 3742
rect 357452 3534 357480 279686
rect 357544 4010 357572 308479
rect 357716 247648 357768 247654
rect 357716 247590 357768 247596
rect 357624 244792 357676 244798
rect 357624 244734 357676 244740
rect 357532 4004 357584 4010
rect 357532 3946 357584 3952
rect 357636 3738 357664 244734
rect 357728 6050 357756 247590
rect 357808 245336 357860 245342
rect 357808 245278 357860 245284
rect 357820 6458 357848 245278
rect 357912 244361 357940 433735
rect 480904 433492 480956 433498
rect 480904 433434 480956 433440
rect 358084 432132 358136 432138
rect 358084 432074 358136 432080
rect 357990 305688 358046 305697
rect 357990 305623 358046 305632
rect 357898 244352 357954 244361
rect 357898 244287 357954 244296
rect 357900 243772 357952 243778
rect 357900 243714 357952 243720
rect 357912 9246 357940 243714
rect 358004 155378 358032 305623
rect 358096 206990 358124 432074
rect 358820 309392 358872 309398
rect 358820 309334 358872 309340
rect 358176 302728 358228 302734
rect 358176 302670 358228 302676
rect 358084 206984 358136 206990
rect 358084 206926 358136 206932
rect 358082 205592 358138 205601
rect 358082 205527 358138 205536
rect 358096 158137 358124 205527
rect 358188 159526 358216 302670
rect 358266 300520 358322 300529
rect 358266 300455 358322 300464
rect 358280 204746 358308 300455
rect 358360 204876 358412 204882
rect 358360 204818 358412 204824
rect 358268 204740 358320 204746
rect 358268 204682 358320 204688
rect 358176 159520 358228 159526
rect 358176 159462 358228 159468
rect 358082 158128 358138 158137
rect 358082 158063 358138 158072
rect 358372 158001 358400 204818
rect 358358 157992 358414 158001
rect 358358 157927 358414 157936
rect 357992 155372 358044 155378
rect 357992 155314 358044 155320
rect 357900 9240 357952 9246
rect 357900 9182 357952 9188
rect 358832 6866 358860 309334
rect 361580 309324 361632 309330
rect 361580 309266 361632 309272
rect 360292 309256 360344 309262
rect 360292 309198 360344 309204
rect 360198 308816 360254 308825
rect 360198 308751 360254 308760
rect 359554 308272 359610 308281
rect 359554 308207 359610 308216
rect 359280 245608 359332 245614
rect 359280 245550 359332 245556
rect 359004 245540 359056 245546
rect 359004 245482 359056 245488
rect 358912 245472 358964 245478
rect 358912 245414 358964 245420
rect 358820 6860 358872 6866
rect 358820 6802 358872 6808
rect 357808 6452 357860 6458
rect 357808 6394 357860 6400
rect 357716 6044 357768 6050
rect 357716 5986 357768 5992
rect 357624 3732 357676 3738
rect 357624 3674 357676 3680
rect 357532 3596 357584 3602
rect 357532 3538 357584 3544
rect 357348 3528 357400 3534
rect 357348 3470 357400 3476
rect 357440 3528 357492 3534
rect 357440 3470 357492 3476
rect 356702 3088 356758 3097
rect 356702 3023 356758 3032
rect 357544 480 357572 3538
rect 358728 3528 358780 3534
rect 358728 3470 358780 3476
rect 358740 480 358768 3470
rect 358924 3398 358952 245414
rect 359016 3874 359044 245482
rect 359188 245404 359240 245410
rect 359188 245346 359240 245352
rect 359096 244860 359148 244866
rect 359096 244802 359148 244808
rect 359004 3868 359056 3874
rect 359004 3810 359056 3816
rect 359108 3641 359136 244802
rect 359200 4078 359228 245346
rect 359188 4072 359240 4078
rect 359188 4014 359240 4020
rect 359094 3632 359150 3641
rect 359094 3567 359150 3576
rect 358912 3392 358964 3398
rect 358912 3334 358964 3340
rect 359292 3262 359320 245550
rect 359372 245268 359424 245274
rect 359372 245210 359424 245216
rect 359384 6390 359412 245210
rect 359464 243704 359516 243710
rect 359464 243646 359516 243652
rect 359476 8974 359504 243646
rect 359568 158545 359596 308207
rect 359648 307896 359700 307902
rect 359648 307838 359700 307844
rect 359660 158982 359688 307838
rect 359648 158976 359700 158982
rect 359648 158918 359700 158924
rect 359554 158536 359610 158545
rect 359554 158471 359610 158480
rect 359464 8968 359516 8974
rect 359464 8910 359516 8916
rect 359372 6384 359424 6390
rect 359372 6326 359424 6332
rect 359922 3496 359978 3505
rect 359922 3431 359978 3440
rect 359280 3256 359332 3262
rect 359280 3198 359332 3204
rect 359936 480 359964 3431
rect 360212 3233 360240 308751
rect 360304 9314 360332 309198
rect 360936 308372 360988 308378
rect 360936 308314 360988 308320
rect 360660 250980 360712 250986
rect 360660 250922 360712 250928
rect 360568 248260 360620 248266
rect 360568 248202 360620 248208
rect 360476 248192 360528 248198
rect 360476 248134 360528 248140
rect 360384 247580 360436 247586
rect 360384 247522 360436 247528
rect 360292 9308 360344 9314
rect 360292 9250 360344 9256
rect 360396 4049 360424 247522
rect 360488 4146 360516 248134
rect 360476 4140 360528 4146
rect 360476 4082 360528 4088
rect 360382 4040 360438 4049
rect 360382 3975 360438 3984
rect 360580 3369 360608 248202
rect 360672 6594 360700 250922
rect 360752 248056 360804 248062
rect 360752 247998 360804 248004
rect 360660 6588 360712 6594
rect 360660 6530 360712 6536
rect 360764 6118 360792 247998
rect 360844 243636 360896 243642
rect 360844 243578 360896 243584
rect 360856 9110 360884 243578
rect 360948 158370 360976 308314
rect 361028 305448 361080 305454
rect 361028 305390 361080 305396
rect 361040 171134 361068 305390
rect 361040 171106 361160 171134
rect 360936 158364 360988 158370
rect 360936 158306 360988 158312
rect 360934 157448 360990 157457
rect 360934 157383 360990 157392
rect 360844 9104 360896 9110
rect 360844 9046 360896 9052
rect 360752 6112 360804 6118
rect 360752 6054 360804 6060
rect 360566 3360 360622 3369
rect 360566 3295 360622 3304
rect 360198 3224 360254 3233
rect 360948 3194 360976 157383
rect 361132 156466 361160 171106
rect 361120 156460 361172 156466
rect 361120 156402 361172 156408
rect 361592 6662 361620 309266
rect 367100 309188 367152 309194
rect 367100 309130 367152 309136
rect 363604 309120 363656 309126
rect 362222 309088 362278 309097
rect 363604 309062 363656 309068
rect 362222 309023 362278 309032
rect 361948 248396 362000 248402
rect 361948 248338 362000 248344
rect 361764 248328 361816 248334
rect 361764 248270 361816 248276
rect 361672 248124 361724 248130
rect 361672 248066 361724 248072
rect 361580 6656 361632 6662
rect 361580 6598 361632 6604
rect 361118 3496 361174 3505
rect 361118 3431 361174 3440
rect 360198 3159 360254 3168
rect 360936 3188 360988 3194
rect 360936 3130 360988 3136
rect 361132 480 361160 3431
rect 361684 3126 361712 248066
rect 361672 3120 361724 3126
rect 361776 3097 361804 248270
rect 361856 247988 361908 247994
rect 361856 247930 361908 247936
rect 361868 3942 361896 247930
rect 361856 3936 361908 3942
rect 361856 3878 361908 3884
rect 361960 3670 361988 248338
rect 362040 245200 362092 245206
rect 362040 245142 362092 245148
rect 362052 3806 362080 245142
rect 362132 243568 362184 243574
rect 362132 243510 362184 243516
rect 362144 9178 362172 243510
rect 362236 158273 362264 309023
rect 362314 308952 362370 308961
rect 362314 308887 362370 308896
rect 362222 158264 362278 158273
rect 362222 158199 362278 158208
rect 362328 157593 362356 308887
rect 362498 308408 362554 308417
rect 362498 308343 362554 308352
rect 362406 306368 362462 306377
rect 362406 306303 362462 306312
rect 362420 171134 362448 306303
rect 362512 245614 362540 308343
rect 363512 308304 363564 308310
rect 363512 308246 363564 308252
rect 363052 251184 363104 251190
rect 363052 251126 363104 251132
rect 362960 251116 363012 251122
rect 362960 251058 363012 251064
rect 362500 245608 362552 245614
rect 362500 245550 362552 245556
rect 362420 171106 362540 171134
rect 362314 157584 362370 157593
rect 362314 157519 362370 157528
rect 362222 157448 362278 157457
rect 362222 157383 362278 157392
rect 362132 9172 362184 9178
rect 362132 9114 362184 9120
rect 362040 3800 362092 3806
rect 362040 3742 362092 3748
rect 361948 3664 362000 3670
rect 361948 3606 362000 3612
rect 361672 3062 361724 3068
rect 361762 3088 361818 3097
rect 362236 3058 362264 157383
rect 362512 157049 362540 171106
rect 362498 157040 362554 157049
rect 362498 156975 362554 156984
rect 362972 6225 363000 251058
rect 363064 6361 363092 251126
rect 363236 251048 363288 251054
rect 363236 250990 363288 250996
rect 363144 250912 363196 250918
rect 363144 250854 363196 250860
rect 363050 6352 363106 6361
rect 363050 6287 363106 6296
rect 362958 6216 363014 6225
rect 362958 6151 363014 6160
rect 363156 5982 363184 250854
rect 363248 6497 363276 250990
rect 363328 245132 363380 245138
rect 363328 245074 363380 245080
rect 363234 6488 363290 6497
rect 363234 6423 363290 6432
rect 363340 6186 363368 245074
rect 363420 244520 363472 244526
rect 363420 244462 363472 244468
rect 363432 9382 363460 244462
rect 363524 157010 363552 308246
rect 363616 158914 363644 309062
rect 364616 309052 364668 309058
rect 364616 308994 364668 309000
rect 364340 308916 364392 308922
rect 364340 308858 364392 308864
rect 363694 303512 363750 303521
rect 363694 303447 363750 303456
rect 363708 159186 363736 303447
rect 363786 302832 363842 302841
rect 363786 302767 363842 302776
rect 363800 204882 363828 302767
rect 363788 204876 363840 204882
rect 363788 204818 363840 204824
rect 363788 204740 363840 204746
rect 363788 204682 363840 204688
rect 363696 159180 363748 159186
rect 363696 159122 363748 159128
rect 363604 158908 363656 158914
rect 363604 158850 363656 158856
rect 363512 157004 363564 157010
rect 363512 156946 363564 156952
rect 363800 155310 363828 204682
rect 364352 158438 364380 308858
rect 364524 308848 364576 308854
rect 364524 308790 364576 308796
rect 364432 308644 364484 308650
rect 364432 308586 364484 308592
rect 364444 158506 364472 308586
rect 364432 158500 364484 158506
rect 364432 158442 364484 158448
rect 364340 158432 364392 158438
rect 364340 158374 364392 158380
rect 364536 158302 364564 308790
rect 364628 158846 364656 308994
rect 364984 308984 365036 308990
rect 364984 308926 365036 308932
rect 364892 308780 364944 308786
rect 364892 308722 364944 308728
rect 364708 308712 364760 308718
rect 364708 308654 364760 308660
rect 364616 158840 364668 158846
rect 364616 158782 364668 158788
rect 364720 158778 364748 308654
rect 364800 308576 364852 308582
rect 364800 308518 364852 308524
rect 364812 158817 364840 308518
rect 364904 158953 364932 308722
rect 364996 159089 365024 308926
rect 366272 306332 366324 306338
rect 366272 306274 366324 306280
rect 365904 306128 365956 306134
rect 365904 306070 365956 306076
rect 365994 306096 366050 306105
rect 365166 303104 365222 303113
rect 365166 303039 365222 303048
rect 365076 300824 365128 300830
rect 365076 300766 365128 300772
rect 364982 159080 365038 159089
rect 364982 159015 365038 159024
rect 364890 158944 364946 158953
rect 364890 158879 364946 158888
rect 364798 158808 364854 158817
rect 364708 158772 364760 158778
rect 364798 158743 364854 158752
rect 364708 158714 364760 158720
rect 364524 158296 364576 158302
rect 364524 158238 364576 158244
rect 365088 155718 365116 300766
rect 365180 158710 365208 303039
rect 365812 247920 365864 247926
rect 365812 247862 365864 247868
rect 365720 245608 365772 245614
rect 365720 245550 365772 245556
rect 365168 158704 365220 158710
rect 365168 158646 365220 158652
rect 365076 155712 365128 155718
rect 365076 155654 365128 155660
rect 363788 155304 363840 155310
rect 363788 155246 363840 155252
rect 363420 9376 363472 9382
rect 363420 9318 363472 9324
rect 365732 6526 365760 245550
rect 365824 9042 365852 247862
rect 365916 156942 365944 306070
rect 365994 306031 366050 306040
rect 366008 157185 366036 306031
rect 366180 305584 366232 305590
rect 366180 305526 366232 305532
rect 366088 305516 366140 305522
rect 366088 305458 366140 305464
rect 365994 157176 366050 157185
rect 365994 157111 366050 157120
rect 365904 156936 365956 156942
rect 365904 156878 365956 156884
rect 366100 156602 366128 305458
rect 366088 156596 366140 156602
rect 366088 156538 366140 156544
rect 366192 156534 366220 305526
rect 366284 156874 366312 306274
rect 366364 306264 366416 306270
rect 366364 306206 366416 306212
rect 366272 156868 366324 156874
rect 366272 156810 366324 156816
rect 366376 156738 366404 306206
rect 366454 303240 366510 303249
rect 366454 303175 366510 303184
rect 366364 156732 366416 156738
rect 366364 156674 366416 156680
rect 366180 156528 366232 156534
rect 366180 156470 366232 156476
rect 366468 155854 366496 303175
rect 366546 300384 366602 300393
rect 366546 300319 366602 300328
rect 366456 155848 366508 155854
rect 366456 155790 366508 155796
rect 366560 155174 366588 300319
rect 366548 155168 366600 155174
rect 366548 155110 366600 155116
rect 365812 9036 365864 9042
rect 365812 8978 365864 8984
rect 367112 6730 367140 309130
rect 367376 308508 367428 308514
rect 367376 308450 367428 308456
rect 367284 308440 367336 308446
rect 367284 308382 367336 308388
rect 367192 244996 367244 245002
rect 367192 244938 367244 244944
rect 367100 6724 367152 6730
rect 367100 6666 367152 6672
rect 365720 6520 365772 6526
rect 365720 6462 365772 6468
rect 367204 6254 367232 244938
rect 367296 156670 367324 308382
rect 367388 157214 367416 308450
rect 437480 307216 437532 307222
rect 437480 307158 437532 307164
rect 368662 306232 368718 306241
rect 367560 306196 367612 306202
rect 368662 306167 368718 306176
rect 367560 306138 367612 306144
rect 367468 305924 367520 305930
rect 367468 305866 367520 305872
rect 367376 157208 367428 157214
rect 367376 157150 367428 157156
rect 367284 156664 367336 156670
rect 367284 156606 367336 156612
rect 367480 155786 367508 305866
rect 367572 156806 367600 306138
rect 367744 306060 367796 306066
rect 367744 306002 367796 306008
rect 367652 305992 367704 305998
rect 367652 305934 367704 305940
rect 367664 157146 367692 305934
rect 367652 157140 367704 157146
rect 367652 157082 367704 157088
rect 367756 157078 367784 306002
rect 367836 305856 367888 305862
rect 367836 305798 367888 305804
rect 367848 159050 367876 305798
rect 368572 305788 368624 305794
rect 368572 305730 368624 305736
rect 367926 303376 367982 303385
rect 367926 303311 367982 303320
rect 367940 159118 367968 303311
rect 368480 245064 368532 245070
rect 368480 245006 368532 245012
rect 367928 159112 367980 159118
rect 367928 159054 367980 159060
rect 367836 159044 367888 159050
rect 367836 158986 367888 158992
rect 367744 157072 367796 157078
rect 367744 157014 367796 157020
rect 367560 156800 367612 156806
rect 367560 156742 367612 156748
rect 367468 155780 367520 155786
rect 367468 155722 367520 155728
rect 368492 6798 368520 245006
rect 368584 157350 368612 305730
rect 368572 157344 368624 157350
rect 368572 157286 368624 157292
rect 368676 155922 368704 306167
rect 368754 305960 368810 305969
rect 368754 305895 368810 305904
rect 368768 157321 368796 305895
rect 378782 305824 378838 305833
rect 378782 305759 378838 305768
rect 368848 305720 368900 305726
rect 368848 305662 368900 305668
rect 368754 157312 368810 157321
rect 368860 157282 368888 305662
rect 368940 305652 368992 305658
rect 368940 305594 368992 305600
rect 368952 158409 368980 305594
rect 371332 303612 371384 303618
rect 371332 303554 371384 303560
rect 370504 303476 370556 303482
rect 370504 303418 370556 303424
rect 369124 303408 369176 303414
rect 369124 303350 369176 303356
rect 369032 300144 369084 300150
rect 369032 300086 369084 300092
rect 368938 158400 368994 158409
rect 368938 158335 368994 158344
rect 368754 157247 368810 157256
rect 368848 157276 368900 157282
rect 368848 157218 368900 157224
rect 368664 155916 368716 155922
rect 368664 155858 368716 155864
rect 369044 155446 369072 300086
rect 369136 159322 369164 303350
rect 369952 303340 370004 303346
rect 369952 303282 370004 303288
rect 369216 302864 369268 302870
rect 369216 302806 369268 302812
rect 369228 159390 369256 302806
rect 369308 300620 369360 300626
rect 369308 300562 369360 300568
rect 369216 159384 369268 159390
rect 369216 159326 369268 159332
rect 369124 159316 369176 159322
rect 369124 159258 369176 159264
rect 369320 158234 369348 300562
rect 369860 247512 369912 247518
rect 369860 247454 369912 247460
rect 369398 158808 369454 158817
rect 369398 158743 369454 158752
rect 369308 158228 369360 158234
rect 369308 158170 369360 158176
rect 369032 155440 369084 155446
rect 369032 155382 369084 155388
rect 369412 6914 369440 158743
rect 369320 6886 369440 6914
rect 368480 6792 368532 6798
rect 368480 6734 368532 6740
rect 367192 6248 367244 6254
rect 367192 6190 367244 6196
rect 363328 6180 363380 6186
rect 363328 6122 363380 6128
rect 363144 5976 363196 5982
rect 363144 5918 363196 5924
rect 367006 3904 367062 3913
rect 367006 3839 367062 3848
rect 362314 3496 362370 3505
rect 362314 3431 362370 3440
rect 363510 3496 363566 3505
rect 363510 3431 363566 3440
rect 364614 3496 364670 3505
rect 364614 3431 364670 3440
rect 365810 3496 365866 3505
rect 365810 3431 365866 3440
rect 361762 3023 361818 3032
rect 362224 3052 362276 3058
rect 362224 2994 362276 3000
rect 362328 480 362356 3431
rect 363524 480 363552 3431
rect 364628 480 364656 3431
rect 365824 480 365852 3431
rect 367020 480 367048 3839
rect 369320 3602 369348 6886
rect 369308 3596 369360 3602
rect 369308 3538 369360 3544
rect 368202 3496 368258 3505
rect 368202 3431 368258 3440
rect 369398 3496 369454 3505
rect 369872 3466 369900 247454
rect 369964 154290 369992 303282
rect 370136 303068 370188 303074
rect 370136 303010 370188 303016
rect 370044 303000 370096 303006
rect 370044 302942 370096 302948
rect 370056 155582 370084 302942
rect 370044 155576 370096 155582
rect 370044 155518 370096 155524
rect 370148 155514 370176 303010
rect 370228 302932 370280 302938
rect 370228 302874 370280 302880
rect 370240 155650 370268 302874
rect 370320 300484 370372 300490
rect 370320 300426 370372 300432
rect 370228 155644 370280 155650
rect 370228 155586 370280 155592
rect 370136 155508 370188 155514
rect 370136 155450 370188 155456
rect 370332 154494 370360 300426
rect 370410 300248 370466 300257
rect 370410 300183 370466 300192
rect 370424 155242 370452 300183
rect 370516 158098 370544 303418
rect 370688 303204 370740 303210
rect 370688 303146 370740 303152
rect 370596 303136 370648 303142
rect 370596 303078 370648 303084
rect 370608 158166 370636 303078
rect 370700 159254 370728 303146
rect 371240 282600 371292 282606
rect 371240 282542 371292 282548
rect 370688 159248 370740 159254
rect 370688 159190 370740 159196
rect 370596 158160 370648 158166
rect 370596 158102 370648 158108
rect 370504 158092 370556 158098
rect 370504 158034 370556 158040
rect 370412 155236 370464 155242
rect 370412 155178 370464 155184
rect 370320 154488 370372 154494
rect 370320 154430 370372 154436
rect 369952 154284 370004 154290
rect 369952 154226 370004 154232
rect 370594 3496 370650 3505
rect 369398 3431 369454 3440
rect 369860 3460 369912 3466
rect 368216 480 368244 3431
rect 369412 480 369440 3431
rect 370594 3431 370650 3440
rect 369860 3402 369912 3408
rect 370608 480 370636 3431
rect 293654 354 293766 480
rect 293328 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371252 354 371280 282542
rect 371344 154222 371372 303554
rect 371608 303544 371660 303550
rect 371608 303486 371660 303492
rect 371424 300552 371476 300558
rect 371424 300494 371476 300500
rect 371436 154426 371464 300494
rect 371516 299940 371568 299946
rect 371516 299882 371568 299888
rect 371424 154420 371476 154426
rect 371424 154362 371476 154368
rect 371332 154216 371384 154222
rect 371332 154158 371384 154164
rect 371528 154154 371556 299882
rect 371620 159458 371648 303486
rect 372988 303272 373040 303278
rect 372988 303214 373040 303220
rect 372712 300756 372764 300762
rect 372712 300698 372764 300704
rect 371792 300280 371844 300286
rect 371792 300222 371844 300228
rect 371700 300008 371752 300014
rect 371700 299950 371752 299956
rect 371608 159452 371660 159458
rect 371608 159394 371660 159400
rect 371712 157962 371740 299950
rect 371804 158642 371832 300222
rect 371884 300076 371936 300082
rect 371884 300018 371936 300024
rect 371792 158636 371844 158642
rect 371792 158578 371844 158584
rect 371700 157956 371752 157962
rect 371700 157898 371752 157904
rect 371896 157894 371924 300018
rect 372620 285252 372672 285258
rect 372620 285194 372672 285200
rect 371884 157888 371936 157894
rect 371884 157830 371936 157836
rect 371516 154148 371568 154154
rect 371516 154090 371568 154096
rect 372632 16574 372660 285194
rect 372724 154086 372752 300698
rect 372804 300416 372856 300422
rect 372804 300358 372856 300364
rect 372816 154358 372844 300358
rect 372896 300212 372948 300218
rect 372896 300154 372948 300160
rect 372908 154562 372936 300154
rect 373000 158030 373028 303214
rect 373080 302796 373132 302802
rect 373080 302738 373132 302744
rect 372988 158024 373040 158030
rect 372988 157966 373040 157972
rect 373092 157826 373120 302738
rect 373264 300688 373316 300694
rect 373264 300630 373316 300636
rect 373172 300348 373224 300354
rect 373172 300290 373224 300296
rect 373184 158574 373212 300290
rect 373276 159594 373304 300630
rect 375380 286680 375432 286686
rect 375380 286622 375432 286628
rect 374000 282532 374052 282538
rect 374000 282474 374052 282480
rect 373264 159588 373316 159594
rect 373264 159530 373316 159536
rect 373172 158568 373224 158574
rect 373172 158510 373224 158516
rect 373080 157820 373132 157826
rect 373080 157762 373132 157768
rect 372896 154556 372948 154562
rect 372896 154498 372948 154504
rect 372804 154352 372856 154358
rect 372804 154294 372856 154300
rect 372712 154080 372764 154086
rect 372712 154022 372764 154028
rect 372632 16546 372936 16574
rect 372908 480 372936 16546
rect 374012 3534 374040 282474
rect 374092 263152 374144 263158
rect 374092 263094 374144 263100
rect 374000 3528 374052 3534
rect 374000 3470 374052 3476
rect 374104 480 374132 263094
rect 375392 16574 375420 286622
rect 378140 283756 378192 283762
rect 378140 283698 378192 283704
rect 376760 264580 376812 264586
rect 376760 264522 376812 264528
rect 376772 16574 376800 264522
rect 378152 16574 378180 283698
rect 375392 16546 376064 16574
rect 376772 16546 377720 16574
rect 378152 16546 378456 16574
rect 375288 3528 375340 3534
rect 375288 3470 375340 3476
rect 375300 480 375328 3470
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 16546
rect 377692 480 377720 16546
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378428 354 378456 16546
rect 378796 3466 378824 305759
rect 422944 291916 422996 291922
rect 422944 291858 422996 291864
rect 407120 289468 407172 289474
rect 407120 289410 407172 289416
rect 382280 288040 382332 288046
rect 382280 287982 382332 287988
rect 380900 264512 380952 264518
rect 380900 264454 380952 264460
rect 379520 254924 379572 254930
rect 379520 254866 379572 254872
rect 378784 3460 378836 3466
rect 378784 3402 378836 3408
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 379532 354 379560 254866
rect 380912 16574 380940 264454
rect 380912 16546 381216 16574
rect 381188 480 381216 16546
rect 382292 1970 382320 287982
rect 386420 287972 386472 287978
rect 386420 287914 386472 287920
rect 385040 283688 385092 283694
rect 385040 283630 385092 283636
rect 382372 278248 382424 278254
rect 382372 278190 382424 278196
rect 382280 1964 382332 1970
rect 382280 1906 382332 1912
rect 382384 480 382412 278190
rect 383660 265940 383712 265946
rect 383660 265882 383712 265888
rect 383672 16574 383700 265882
rect 385052 16574 385080 283630
rect 386432 16574 386460 287914
rect 400220 287904 400272 287910
rect 400220 287846 400272 287852
rect 397460 286612 397512 286618
rect 397460 286554 397512 286560
rect 391940 285184 391992 285190
rect 391940 285126 391992 285132
rect 389180 283620 389232 283626
rect 389180 283562 389232 283568
rect 387800 265872 387852 265878
rect 387800 265814 387852 265820
rect 383672 16546 384344 16574
rect 385052 16546 386000 16574
rect 386432 16546 386736 16574
rect 383568 1964 383620 1970
rect 383568 1906 383620 1912
rect 383580 480 383608 1906
rect 379950 354 380062 480
rect 379532 326 380062 354
rect 378846 -960 378958 326
rect 379950 -960 380062 326
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 354 384344 16546
rect 385972 480 386000 16546
rect 384734 354 384846 480
rect 384316 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 386708 354 386736 16546
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387812 354 387840 265814
rect 389192 16574 389220 283562
rect 390560 267300 390612 267306
rect 390560 267242 390612 267248
rect 389192 16546 389496 16574
rect 389468 480 389496 16546
rect 390572 3534 390600 267242
rect 390652 254856 390704 254862
rect 390652 254798 390704 254804
rect 390560 3528 390612 3534
rect 390560 3470 390612 3476
rect 390664 480 390692 254798
rect 391952 16574 391980 285126
rect 396080 285116 396132 285122
rect 396080 285058 396132 285064
rect 393320 275664 393372 275670
rect 393320 275606 393372 275612
rect 393332 16574 393360 275606
rect 394700 267232 394752 267238
rect 394700 267174 394752 267180
rect 394712 16574 394740 267174
rect 391952 16546 392624 16574
rect 393332 16546 394280 16574
rect 394712 16546 395384 16574
rect 391848 3528 391900 3534
rect 391848 3470 391900 3476
rect 391860 480 391888 3470
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 387126 -960 387238 326
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 394252 480 394280 16546
rect 395356 480 395384 16546
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 285058
rect 397472 16574 397500 286554
rect 398840 285048 398892 285054
rect 398840 284990 398892 284996
rect 397472 16546 397776 16574
rect 397748 480 397776 16546
rect 398852 2242 398880 284990
rect 398932 268728 398984 268734
rect 398932 268670 398984 268676
rect 398840 2236 398892 2242
rect 398840 2178 398892 2184
rect 398944 480 398972 268670
rect 400232 16574 400260 287846
rect 404360 287836 404412 287842
rect 404360 287778 404412 287784
rect 402980 282464 403032 282470
rect 402980 282406 403032 282412
rect 401600 270156 401652 270162
rect 401600 270098 401652 270104
rect 401612 16574 401640 270098
rect 402992 16574 403020 282406
rect 400232 16546 400904 16574
rect 401612 16546 402560 16574
rect 402992 16546 403664 16574
rect 400128 2236 400180 2242
rect 400128 2178 400180 2184
rect 400140 480 400168 2178
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 16546
rect 402532 480 402560 16546
rect 403636 480 403664 16546
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 287778
rect 405740 265804 405792 265810
rect 405740 265746 405792 265752
rect 405752 16574 405780 265746
rect 405752 16546 406056 16574
rect 406028 480 406056 16546
rect 407132 2242 407160 289410
rect 413284 289400 413336 289406
rect 413284 289342 413336 289348
rect 411260 289332 411312 289338
rect 411260 289274 411312 289280
rect 407212 272740 407264 272746
rect 407212 272682 407264 272688
rect 407120 2236 407172 2242
rect 407120 2178 407172 2184
rect 407224 480 407252 272682
rect 408500 271448 408552 271454
rect 408500 271390 408552 271396
rect 408512 16574 408540 271390
rect 409880 250844 409932 250850
rect 409880 250786 409932 250792
rect 409892 16574 409920 250786
rect 411272 16574 411300 289274
rect 412640 272672 412692 272678
rect 412640 272614 412692 272620
rect 408512 16546 409184 16574
rect 409892 16546 410840 16574
rect 411272 16546 411944 16574
rect 408408 2236 408460 2242
rect 408408 2178 408460 2184
rect 408420 480 408448 2178
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 410812 480 410840 16546
rect 411916 480 411944 16546
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 272614
rect 413296 3602 413324 289342
rect 415400 289264 415452 289270
rect 415400 289206 415452 289212
rect 414020 284980 414072 284986
rect 414020 284922 414072 284928
rect 414032 16574 414060 284922
rect 414032 16546 414336 16574
rect 413284 3596 413336 3602
rect 413284 3538 413336 3544
rect 414308 480 414336 16546
rect 415412 3346 415440 289206
rect 418160 289196 418212 289202
rect 418160 289138 418212 289144
rect 416780 286544 416832 286550
rect 416780 286486 416832 286492
rect 415492 274304 415544 274310
rect 415492 274246 415544 274252
rect 415504 3534 415532 274246
rect 416792 16574 416820 286486
rect 418172 16574 418200 289138
rect 419540 275596 419592 275602
rect 419540 275538 419592 275544
rect 419552 16574 419580 275538
rect 422300 256420 422352 256426
rect 422300 256362 422352 256368
rect 420920 252136 420972 252142
rect 420920 252078 420972 252084
rect 416792 16546 417464 16574
rect 418172 16546 418568 16574
rect 419552 16546 420224 16574
rect 415492 3528 415544 3534
rect 415492 3470 415544 3476
rect 416688 3528 416740 3534
rect 416688 3470 416740 3476
rect 415412 3318 415532 3346
rect 415504 480 415532 3318
rect 416700 480 416728 3470
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16546
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 418540 354 418568 16546
rect 420196 480 420224 16546
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 252078
rect 422312 16574 422340 256362
rect 422312 16546 422616 16574
rect 422588 480 422616 16546
rect 422956 3534 422984 291858
rect 431960 290488 432012 290494
rect 431960 290430 432012 290436
rect 426440 281036 426492 281042
rect 426440 280978 426492 280984
rect 423772 275528 423824 275534
rect 423772 275470 423824 275476
rect 422944 3528 422996 3534
rect 422944 3470 422996 3476
rect 423784 480 423812 275470
rect 426452 16574 426480 280978
rect 430580 279676 430632 279682
rect 430580 279618 430632 279624
rect 427820 267164 427872 267170
rect 427820 267106 427872 267112
rect 426452 16546 426848 16574
rect 426164 3596 426216 3602
rect 426164 3538 426216 3544
rect 424968 3528 425020 3534
rect 424968 3470 425020 3476
rect 424980 480 425008 3470
rect 426176 480 426204 3538
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 426820 354 426848 16546
rect 427832 6914 427860 267106
rect 428464 256284 428516 256290
rect 428464 256226 428516 256232
rect 428476 16574 428504 256226
rect 430592 16574 430620 279618
rect 428476 16546 428596 16574
rect 430592 16546 430896 16574
rect 427832 6886 428504 6914
rect 428476 480 428504 6886
rect 428568 3534 428596 16546
rect 428556 3528 428608 3534
rect 428556 3470 428608 3476
rect 429660 3528 429712 3534
rect 429660 3470 429712 3476
rect 429672 480 429700 3470
rect 430868 480 430896 16546
rect 431972 3534 432000 290430
rect 433340 277024 433392 277030
rect 433340 276966 433392 276972
rect 432052 244928 432104 244934
rect 432052 244870 432104 244876
rect 431960 3528 432012 3534
rect 431960 3470 432012 3476
rect 432064 480 432092 244870
rect 433352 16574 433380 276966
rect 434720 275460 434772 275466
rect 434720 275402 434772 275408
rect 434732 16574 434760 275402
rect 436100 256216 436152 256222
rect 436100 256158 436152 256164
rect 436112 16574 436140 256158
rect 433352 16546 434024 16574
rect 434732 16546 435128 16574
rect 436112 16546 436784 16574
rect 433248 3528 433300 3534
rect 433248 3470 433300 3476
rect 433260 480 433288 3470
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 16546
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 16546
rect 436756 480 436784 16546
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437492 354 437520 307158
rect 467102 300112 467158 300121
rect 467102 300047 467158 300056
rect 440240 280900 440292 280906
rect 440240 280842 440292 280848
rect 438860 265736 438912 265742
rect 438860 265678 438912 265684
rect 438872 16574 438900 265678
rect 438872 16546 439176 16574
rect 439148 480 439176 16546
rect 440252 3346 440280 280842
rect 440332 278180 440384 278186
rect 440332 278122 440384 278128
rect 440344 3534 440372 278122
rect 449900 272604 449952 272610
rect 449900 272546 449952 272552
rect 447140 268660 447192 268666
rect 447140 268602 447192 268608
rect 441620 263084 441672 263090
rect 441620 263026 441672 263032
rect 441632 16574 441660 263026
rect 444380 263016 444432 263022
rect 444380 262958 444432 262964
rect 443000 256148 443052 256154
rect 443000 256090 443052 256096
rect 443012 16574 443040 256090
rect 444392 16574 444420 262958
rect 445760 250776 445812 250782
rect 445760 250718 445812 250724
rect 441632 16546 442672 16574
rect 443012 16546 443408 16574
rect 444392 16546 445064 16574
rect 440332 3528 440384 3534
rect 440332 3470 440384 3476
rect 441528 3528 441580 3534
rect 441528 3470 441580 3476
rect 440252 3318 440372 3346
rect 440344 480 440372 3318
rect 441540 480 441568 3470
rect 442644 480 442672 16546
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 354 443408 16546
rect 445036 480 445064 16546
rect 443798 354 443910 480
rect 443380 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 445772 354 445800 250718
rect 447152 16574 447180 268602
rect 448520 264444 448572 264450
rect 448520 264386 448572 264392
rect 447152 16546 447456 16574
rect 447428 480 447456 16546
rect 448532 3346 448560 264386
rect 448612 247852 448664 247858
rect 448612 247794 448664 247800
rect 448624 3534 448652 247794
rect 449912 16574 449940 272546
rect 465080 271380 465132 271386
rect 465080 271322 465132 271328
rect 458180 270088 458232 270094
rect 458180 270030 458232 270036
rect 455420 268592 455472 268598
rect 455420 268534 455472 268540
rect 451280 267096 451332 267102
rect 451280 267038 451332 267044
rect 451292 16574 451320 267038
rect 452660 249348 452712 249354
rect 452660 249290 452712 249296
rect 452672 16574 452700 249290
rect 454040 247784 454092 247790
rect 454040 247726 454092 247732
rect 449912 16546 450952 16574
rect 451292 16546 451688 16574
rect 452672 16546 453344 16574
rect 448612 3528 448664 3534
rect 448612 3470 448664 3476
rect 449808 3528 449860 3534
rect 449808 3470 449860 3476
rect 448532 3318 448652 3346
rect 448624 480 448652 3318
rect 449820 480 449848 3470
rect 450924 480 450952 16546
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 453316 480 453344 16546
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454052 354 454080 247726
rect 455432 16574 455460 268534
rect 456800 253564 456852 253570
rect 456800 253506 456852 253512
rect 455432 16546 455736 16574
rect 455708 480 455736 16546
rect 456812 2242 456840 253506
rect 456892 249280 456944 249286
rect 456892 249222 456944 249228
rect 456800 2236 456852 2242
rect 456800 2178 456852 2184
rect 456904 480 456932 249222
rect 458192 16574 458220 270030
rect 462320 261724 462372 261730
rect 462320 261666 462372 261672
rect 460940 254788 460992 254794
rect 460940 254730 460992 254736
rect 459560 252068 459612 252074
rect 459560 252010 459612 252016
rect 459572 16574 459600 252010
rect 460952 16574 460980 254730
rect 458192 16546 459232 16574
rect 459572 16546 459968 16574
rect 460952 16546 461624 16574
rect 458088 2236 458140 2242
rect 458088 2178 458140 2184
rect 458100 480 458128 2178
rect 459204 480 459232 16546
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 461596 480 461624 16546
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462332 354 462360 261666
rect 463700 261656 463752 261662
rect 463700 261598 463752 261604
rect 463712 16574 463740 261598
rect 463712 16546 464016 16574
rect 463988 480 464016 16546
rect 465092 3534 465120 271322
rect 465172 270020 465224 270026
rect 465172 269962 465224 269968
rect 465080 3528 465132 3534
rect 465080 3470 465132 3476
rect 465184 480 465212 269962
rect 466460 262948 466512 262954
rect 466460 262890 466512 262896
rect 466472 16574 466500 262890
rect 466472 16546 467052 16574
rect 465908 3528 465960 3534
rect 465908 3470 465960 3476
rect 467024 3482 467052 16546
rect 467116 4146 467144 300047
rect 471244 294636 471296 294642
rect 471244 294578 471296 294584
rect 469220 274236 469272 274242
rect 469220 274178 469272 274184
rect 467838 245304 467894 245313
rect 467838 245239 467894 245248
rect 467852 16574 467880 245239
rect 469232 16574 469260 274178
rect 467852 16546 468248 16574
rect 469232 16546 469904 16574
rect 467104 4140 467156 4146
rect 467104 4082 467156 4088
rect 467656 4140 467708 4146
rect 467656 4082 467708 4088
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465920 354 465948 3470
rect 467024 3454 467512 3482
rect 467484 480 467512 3454
rect 467668 3058 467696 4082
rect 467656 3052 467708 3058
rect 467656 2994 467708 3000
rect 466246 354 466358 480
rect 465920 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468220 354 468248 16546
rect 469876 480 469904 16546
rect 471256 3534 471284 294578
rect 471980 287768 472032 287774
rect 471980 287710 472032 287716
rect 471992 16574 472020 287710
rect 475384 282328 475436 282334
rect 475384 282270 475436 282276
rect 473452 274168 473504 274174
rect 473452 274110 473504 274116
rect 473464 16574 473492 274110
rect 474740 261588 474792 261594
rect 474740 261530 474792 261536
rect 474752 16574 474780 261530
rect 471992 16546 472296 16574
rect 473464 16546 474136 16574
rect 474752 16546 475332 16574
rect 471244 3528 471296 3534
rect 471244 3470 471296 3476
rect 471060 3052 471112 3058
rect 471060 2994 471112 3000
rect 471072 480 471100 2994
rect 472268 480 472296 16546
rect 473452 3528 473504 3534
rect 473452 3470 473504 3476
rect 473464 480 473492 3470
rect 468638 354 468750 480
rect 468220 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 16546
rect 475304 3482 475332 16546
rect 475396 3602 475424 282270
rect 476764 274100 476816 274106
rect 476764 274042 476816 274048
rect 475384 3596 475436 3602
rect 475384 3538 475436 3544
rect 475304 3454 475792 3482
rect 475764 480 475792 3454
rect 476776 3126 476804 274042
rect 477500 247716 477552 247722
rect 477500 247658 477552 247664
rect 477512 16574 477540 247658
rect 480258 245168 480314 245177
rect 480258 245103 480314 245112
rect 480272 16574 480300 245103
rect 477512 16546 478184 16574
rect 480272 16546 480576 16574
rect 476948 3596 477000 3602
rect 476948 3538 477000 3544
rect 476764 3120 476816 3126
rect 476764 3062 476816 3068
rect 476960 480 476988 3538
rect 478156 480 478184 16546
rect 479340 3120 479392 3126
rect 479340 3062 479392 3068
rect 479352 480 479380 3062
rect 480548 480 480576 16546
rect 480916 3534 480944 433434
rect 500960 307080 501012 307086
rect 500960 307022 501012 307028
rect 488540 287700 488592 287706
rect 488540 287642 488592 287648
rect 481640 280832 481692 280838
rect 481640 280774 481692 280780
rect 481652 6914 481680 280774
rect 484400 271312 484452 271318
rect 484400 271254 484452 271260
rect 483018 247888 483074 247897
rect 483018 247823 483074 247832
rect 481730 245032 481786 245041
rect 481730 244967 481786 244976
rect 481744 16574 481772 244967
rect 483032 16574 483060 247823
rect 484412 16574 484440 271254
rect 485780 253496 485832 253502
rect 485780 253438 485832 253444
rect 485792 16574 485820 253438
rect 487160 250708 487212 250714
rect 487160 250650 487212 250656
rect 481744 16546 482416 16574
rect 483032 16546 484072 16574
rect 484412 16546 484808 16574
rect 485792 16546 486464 16574
rect 481652 6886 481772 6914
rect 480904 3528 480956 3534
rect 480904 3470 480956 3476
rect 481744 480 481772 6886
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 354 482416 16546
rect 484044 480 484072 16546
rect 482806 354 482918 480
rect 482388 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 486436 480 486464 16546
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487172 354 487200 250650
rect 488552 16574 488580 287642
rect 492680 286408 492732 286414
rect 492680 286350 492732 286356
rect 491300 279608 491352 279614
rect 491300 279550 491352 279556
rect 489920 253428 489972 253434
rect 489920 253370 489972 253376
rect 488552 16546 488856 16574
rect 488828 480 488856 16546
rect 489932 480 489960 253370
rect 490012 249212 490064 249218
rect 490012 249154 490064 249160
rect 490024 16574 490052 249154
rect 491312 16574 491340 279550
rect 492692 16574 492720 286350
rect 498200 275392 498252 275398
rect 498200 275334 498252 275340
rect 495440 269952 495492 269958
rect 495440 269894 495492 269900
rect 494060 250640 494112 250646
rect 494060 250582 494112 250588
rect 494072 16574 494100 250582
rect 490024 16546 490696 16574
rect 491312 16546 492352 16574
rect 492692 16546 493088 16574
rect 494072 16546 494744 16574
rect 487590 354 487702 480
rect 487172 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490668 354 490696 16546
rect 492324 480 492352 16546
rect 491086 354 491198 480
rect 490668 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 494716 480 494744 16546
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 269894
rect 496084 261520 496136 261526
rect 496084 261462 496136 261468
rect 496096 3602 496124 261462
rect 498212 3602 498240 275334
rect 499580 264376 499632 264382
rect 499580 264318 499632 264324
rect 498292 254720 498344 254726
rect 498292 254662 498344 254668
rect 496084 3596 496136 3602
rect 496084 3538 496136 3544
rect 497096 3596 497148 3602
rect 497096 3538 497148 3544
rect 498200 3596 498252 3602
rect 498200 3538 498252 3544
rect 497108 480 497136 3538
rect 498304 3482 498332 254662
rect 499592 16574 499620 264318
rect 500972 16574 501000 307022
rect 538864 298784 538916 298790
rect 538864 298726 538916 298732
rect 509240 286340 509292 286346
rect 509240 286282 509292 286288
rect 506572 276956 506624 276962
rect 506572 276898 506624 276904
rect 504364 269884 504416 269890
rect 504364 269826 504416 269832
rect 502340 268524 502392 268530
rect 502340 268466 502392 268472
rect 502352 16574 502380 268466
rect 503720 268456 503772 268462
rect 503720 268398 503772 268404
rect 499592 16546 500632 16574
rect 500972 16546 501368 16574
rect 502352 16546 503024 16574
rect 499028 3596 499080 3602
rect 499028 3538 499080 3544
rect 498212 3454 498332 3482
rect 498212 480 498240 3454
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499040 354 499068 3538
rect 500604 480 500632 16546
rect 499366 354 499478 480
rect 499040 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501340 354 501368 16546
rect 502996 480 503024 16546
rect 501758 354 501870 480
rect 501340 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 503732 354 503760 268398
rect 504376 3602 504404 269826
rect 505100 256080 505152 256086
rect 505100 256022 505152 256028
rect 505112 16574 505140 256022
rect 505112 16546 505416 16574
rect 504364 3596 504416 3602
rect 504364 3538 504416 3544
rect 505388 480 505416 16546
rect 506584 6914 506612 276898
rect 507860 253360 507912 253366
rect 507860 253302 507912 253308
rect 507872 16574 507900 253302
rect 509252 16574 509280 286282
rect 524420 282260 524472 282266
rect 524420 282202 524472 282208
rect 511264 276888 511316 276894
rect 511264 276830 511316 276836
rect 510620 246628 510672 246634
rect 510620 246570 510672 246576
rect 510632 16574 510660 246570
rect 507872 16546 508912 16574
rect 509252 16546 509648 16574
rect 510632 16546 511212 16574
rect 506492 6886 506612 6914
rect 506492 480 506520 6886
rect 507676 3596 507728 3602
rect 507676 3538 507728 3544
rect 507688 480 507716 3538
rect 508884 480 508912 16546
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 511184 3482 511212 16546
rect 511276 3602 511304 276830
rect 516140 274032 516192 274038
rect 516140 273974 516192 273980
rect 514024 267028 514076 267034
rect 514024 266970 514076 266976
rect 512000 256012 512052 256018
rect 512000 255954 512052 255960
rect 511264 3596 511316 3602
rect 511264 3538 511316 3544
rect 511184 3454 511304 3482
rect 511276 480 511304 3454
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 255954
rect 514036 3602 514064 266970
rect 514852 257508 514904 257514
rect 514852 257450 514904 257456
rect 514864 16574 514892 257450
rect 516152 16574 516180 273974
rect 521660 264308 521712 264314
rect 521660 264250 521712 264256
rect 518900 252000 518952 252006
rect 518900 251942 518952 251948
rect 517520 250572 517572 250578
rect 517520 250514 517572 250520
rect 517532 16574 517560 250514
rect 518912 16574 518940 251942
rect 520278 247752 520334 247761
rect 520278 247687 520334 247696
rect 514864 16546 515536 16574
rect 516152 16546 517192 16574
rect 517532 16546 517928 16574
rect 518912 16546 519584 16574
rect 513564 3596 513616 3602
rect 513564 3538 513616 3544
rect 514024 3596 514076 3602
rect 514024 3538 514076 3544
rect 514760 3596 514812 3602
rect 514760 3538 514812 3544
rect 513576 480 513604 3538
rect 514772 480 514800 3538
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 512430 -960 512542 326
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515508 354 515536 16546
rect 517164 480 517192 16546
rect 515926 354 516038 480
rect 515508 326 516038 354
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 519556 480 519584 16546
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 247687
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 264250
rect 523040 257440 523092 257446
rect 523040 257382 523092 257388
rect 523052 480 523080 257382
rect 523132 249144 523184 249150
rect 523132 249086 523184 249092
rect 523144 16574 523172 249086
rect 524432 16574 524460 282202
rect 534080 278112 534132 278118
rect 534080 278054 534132 278060
rect 531320 276820 531372 276826
rect 531320 276762 531372 276768
rect 527180 275324 527232 275330
rect 527180 275266 527232 275272
rect 525800 258800 525852 258806
rect 525800 258742 525852 258748
rect 525812 16574 525840 258742
rect 527192 16574 527220 275266
rect 528560 271244 528612 271250
rect 528560 271186 528612 271192
rect 523144 16546 523816 16574
rect 524432 16546 525472 16574
rect 525812 16546 526208 16574
rect 527192 16546 527864 16574
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523788 354 523816 16546
rect 525444 480 525472 16546
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527836 480 527864 16546
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 271186
rect 529940 258732 529992 258738
rect 529940 258674 529992 258680
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 258674
rect 531332 480 531360 276762
rect 531412 265668 531464 265674
rect 531412 265610 531464 265616
rect 531424 16574 531452 265610
rect 532700 260364 532752 260370
rect 532700 260306 532752 260312
rect 532712 16574 532740 260306
rect 534092 16574 534120 278054
rect 538220 273964 538272 273970
rect 538220 273906 538272 273912
rect 536840 260296 536892 260302
rect 536840 260238 536892 260244
rect 535460 253292 535512 253298
rect 535460 253234 535512 253240
rect 535472 16574 535500 253234
rect 536852 16574 536880 260238
rect 531424 16546 532096 16574
rect 532712 16546 533752 16574
rect 534092 16546 534488 16574
rect 535472 16546 536144 16574
rect 536852 16546 537248 16574
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532068 354 532096 16546
rect 533724 480 533752 16546
rect 532486 354 532598 480
rect 532068 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 536116 480 536144 16546
rect 537220 480 537248 16546
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 273906
rect 538876 3602 538904 298726
rect 567844 297424 567896 297430
rect 567844 297366 567896 297372
rect 543740 293344 543792 293350
rect 543740 293286 543792 293292
rect 540980 278044 541032 278050
rect 540980 277986 541032 277992
rect 539600 264240 539652 264246
rect 539600 264182 539652 264188
rect 538864 3596 538916 3602
rect 538864 3538 538916 3544
rect 539612 480 539640 264182
rect 539692 260228 539744 260234
rect 539692 260170 539744 260176
rect 539704 16574 539732 260170
rect 540992 16574 541020 277986
rect 542360 276752 542412 276758
rect 542360 276694 542412 276700
rect 542372 16574 542400 276694
rect 543752 16574 543780 293286
rect 547880 291848 547932 291854
rect 547880 291790 547932 291796
rect 546500 276684 546552 276690
rect 546500 276626 546552 276632
rect 545118 244896 545174 244905
rect 545118 244831 545174 244840
rect 545132 16574 545160 244831
rect 539704 16546 540376 16574
rect 540992 16546 542032 16574
rect 542372 16546 542768 16574
rect 543752 16546 544424 16574
rect 545132 16546 545528 16574
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540348 354 540376 16546
rect 542004 480 542032 16546
rect 540766 354 540878 480
rect 540348 326 540878 354
rect 540766 -960 540878 326
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 544396 480 544424 16546
rect 545500 480 545528 16546
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 276626
rect 547892 480 547920 291790
rect 547972 279540 548024 279546
rect 547972 279482 548024 279488
rect 547984 16574 548012 279482
rect 556160 279472 556212 279478
rect 556160 279414 556212 279420
rect 552020 271176 552072 271182
rect 552020 271118 552072 271124
rect 549260 251932 549312 251938
rect 549260 251874 549312 251880
rect 549272 16574 549300 251874
rect 552032 16574 552060 271118
rect 553400 246560 553452 246566
rect 553400 246502 553452 246508
rect 553412 16574 553440 246502
rect 554780 246492 554832 246498
rect 554780 246434 554832 246440
rect 547984 16546 548656 16574
rect 549272 16546 550312 16574
rect 552032 16546 552704 16574
rect 553412 16546 553808 16574
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 548628 354 548656 16546
rect 550284 480 550312 16546
rect 551468 3596 551520 3602
rect 551468 3538 551520 3544
rect 551480 480 551508 3538
rect 552676 480 552704 16546
rect 553780 480 553808 16546
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 246434
rect 556172 480 556200 279414
rect 558920 269816 558972 269822
rect 558920 269758 558972 269764
rect 556252 254652 556304 254658
rect 556252 254594 556304 254600
rect 556264 16574 556292 254594
rect 557538 247616 557594 247625
rect 557538 247551 557594 247560
rect 557552 16574 557580 247551
rect 558932 16574 558960 269758
rect 565820 268388 565872 268394
rect 565820 268330 565872 268336
rect 564440 257372 564492 257378
rect 564440 257314 564492 257320
rect 560300 254584 560352 254590
rect 560300 254526 560352 254532
rect 560312 16574 560340 254526
rect 561680 253224 561732 253230
rect 561680 253166 561732 253172
rect 561692 16574 561720 253166
rect 563060 246424 563112 246430
rect 563060 246366 563112 246372
rect 556264 16546 556936 16574
rect 557552 16546 558592 16574
rect 558932 16546 559328 16574
rect 560312 16546 560432 16574
rect 561692 16546 562088 16574
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 556908 354 556936 16546
rect 558564 480 558592 16546
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 16546
rect 562060 480 562088 16546
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563072 354 563100 246366
rect 564452 3602 564480 257314
rect 564532 251864 564584 251870
rect 564532 251806 564584 251812
rect 564440 3596 564492 3602
rect 564440 3538 564492 3544
rect 564544 3482 564572 251806
rect 565832 16574 565860 268330
rect 567200 249076 567252 249082
rect 567200 249018 567252 249024
rect 567212 16574 567240 249018
rect 565832 16546 566872 16574
rect 567212 16546 567608 16574
rect 565268 3596 565320 3602
rect 565268 3538 565320 3544
rect 564452 3454 564572 3482
rect 564452 480 564480 3454
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565280 354 565308 3538
rect 566844 480 566872 16546
rect 565606 354 565718 480
rect 565280 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 567856 3262 567884 297366
rect 571984 293276 572036 293282
rect 571984 293218 572036 293224
rect 569960 272536 570012 272542
rect 569960 272478 570012 272484
rect 568580 260160 568632 260166
rect 568580 260102 568632 260108
rect 568592 16574 568620 260102
rect 569972 16574 570000 272478
rect 568592 16546 568712 16574
rect 569972 16546 570368 16574
rect 567844 3256 567896 3262
rect 567844 3198 567896 3204
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 568684 354 568712 16546
rect 570340 480 570368 16546
rect 571524 3256 571576 3262
rect 571524 3198 571576 3204
rect 571536 480 571564 3198
rect 571996 3058 572024 293218
rect 575480 289128 575532 289134
rect 575480 289070 575532 289076
rect 574100 282192 574152 282198
rect 574100 282134 574152 282140
rect 574112 16574 574140 282134
rect 575492 16574 575520 289070
rect 576860 250504 576912 250510
rect 576860 250446 576912 250452
rect 576872 16574 576900 250446
rect 577516 179382 577544 434726
rect 579986 433664 580042 433673
rect 579986 433599 580042 433608
rect 579896 431928 579948 431934
rect 579896 431870 579948 431876
rect 579908 431633 579936 431870
rect 579894 431624 579950 431633
rect 579894 431559 579950 431568
rect 577594 430672 577650 430681
rect 577594 430607 577650 430616
rect 577608 219230 577636 430607
rect 580000 427174 580028 433599
rect 580446 433528 580502 433537
rect 580446 433463 580502 433472
rect 580262 433392 580318 433401
rect 580262 433327 580318 433336
rect 580172 432812 580224 432818
rect 580172 432754 580224 432760
rect 580080 432608 580132 432614
rect 580080 432550 580132 432556
rect 579988 427168 580040 427174
rect 579988 427110 580040 427116
rect 579988 419484 580040 419490
rect 579988 419426 580040 419432
rect 580000 418305 580028 419426
rect 579986 418296 580042 418305
rect 579986 418231 580042 418240
rect 579988 405680 580040 405686
rect 579988 405622 580040 405628
rect 580000 404977 580028 405622
rect 579986 404968 580042 404977
rect 579986 404903 580042 404912
rect 580092 378457 580120 432550
rect 580078 378448 580134 378457
rect 580078 378383 580134 378392
rect 580184 365129 580212 432754
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 580172 325644 580224 325650
rect 580172 325586 580224 325592
rect 580184 325281 580212 325586
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 579988 273216 580040 273222
rect 579988 273158 580040 273164
rect 580000 272241 580028 273158
rect 579986 272232 580042 272241
rect 579986 272167 580042 272176
rect 578240 262880 578292 262886
rect 578240 262822 578292 262828
rect 577596 219224 577648 219230
rect 577596 219166 577648 219172
rect 577504 179376 577556 179382
rect 577504 179318 577556 179324
rect 578252 16574 578280 262822
rect 579804 259412 579856 259418
rect 579804 259354 579856 259360
rect 579816 258913 579844 259354
rect 579802 258904 579858 258913
rect 579802 258839 579858 258848
rect 580172 246356 580224 246362
rect 580172 246298 580224 246304
rect 580184 245585 580212 246298
rect 580170 245576 580226 245585
rect 580170 245511 580226 245520
rect 579712 219224 579764 219230
rect 579712 219166 579764 219172
rect 579724 219065 579752 219166
rect 579710 219056 579766 219065
rect 579710 218991 579766 219000
rect 579620 206984 579672 206990
rect 579620 206926 579672 206932
rect 579632 205737 579660 206926
rect 579618 205728 579674 205737
rect 579618 205663 579674 205672
rect 579712 179376 579764 179382
rect 579712 179318 579764 179324
rect 579724 179217 579752 179318
rect 579710 179208 579766 179217
rect 579710 179143 579766 179152
rect 574112 16546 575152 16574
rect 575492 16546 575888 16574
rect 576872 16546 576992 16574
rect 578252 16546 578648 16574
rect 572720 3460 572772 3466
rect 572720 3402 572772 3408
rect 571984 3052 572036 3058
rect 571984 2994 572036 3000
rect 572732 480 572760 3402
rect 573916 3052 573968 3058
rect 573916 2994 573968 3000
rect 573928 480 573956 2994
rect 575124 480 575152 16546
rect 569102 354 569214 480
rect 568684 326 569214 354
rect 567998 -960 568110 326
rect 569102 -960 569214 326
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 575860 354 575888 16546
rect 576278 354 576390 480
rect 575860 326 576390 354
rect 576964 354 576992 16546
rect 578620 480 578648 16546
rect 580276 6633 580304 433327
rect 580356 431996 580408 432002
rect 580356 431938 580408 431944
rect 580368 33153 580396 431938
rect 580460 126041 580488 433463
rect 580552 152697 580580 434794
rect 580632 432744 580684 432750
rect 580632 432686 580684 432692
rect 580644 427258 580672 432686
rect 580724 432676 580776 432682
rect 580724 432618 580776 432624
rect 580736 427378 580764 432618
rect 580724 427372 580776 427378
rect 580724 427314 580776 427320
rect 580644 427230 580856 427258
rect 580632 427168 580684 427174
rect 580632 427110 580684 427116
rect 580724 427168 580776 427174
rect 580724 427110 580776 427116
rect 580538 152688 580594 152697
rect 580538 152623 580594 152632
rect 580644 139369 580672 427110
rect 580736 192545 580764 427110
rect 580828 232393 580856 427230
rect 580920 312089 580948 434862
rect 581092 433424 581144 433430
rect 581092 433366 581144 433372
rect 580906 312080 580962 312089
rect 580906 312015 580962 312024
rect 580814 232384 580870 232393
rect 580814 232319 580870 232328
rect 580722 192536 580778 192545
rect 580722 192471 580778 192480
rect 580630 139360 580686 139369
rect 580630 139295 580686 139304
rect 580446 126032 580502 126041
rect 580446 125967 580502 125976
rect 580354 33144 580410 33153
rect 580354 33079 580410 33088
rect 581104 16574 581132 433366
rect 582380 433356 582432 433362
rect 582380 433298 582432 433304
rect 582392 16574 582420 433298
rect 581104 16546 581776 16574
rect 582392 16546 583432 16574
rect 580262 6624 580318 6633
rect 580262 6559 580318 6568
rect 581000 3528 581052 3534
rect 581000 3470 581052 3476
rect 581012 480 581040 3470
rect 577382 354 577494 480
rect 576964 326 577494 354
rect 576278 -960 576390 326
rect 577382 -960 577494 326
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 581748 354 581776 16546
rect 583404 480 583432 16546
rect 582166 354 582278 480
rect 581748 326 582278 354
rect 582166 -960 582278 326
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3422 606076 3478 606112
rect 3422 606056 3424 606076
rect 3424 606056 3476 606076
rect 3476 606056 3478 606076
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3422 553832 3478 553888
rect 2778 527856 2834 527912
rect 3422 514800 3478 514856
rect 3054 501744 3110 501800
rect 3422 475632 3478 475688
rect 3238 462576 3294 462632
rect 3146 449520 3202 449576
rect 217782 516840 217838 516896
rect 217690 515888 217746 515944
rect 217598 513712 217654 513768
rect 217414 489912 217470 489968
rect 217322 488008 217378 488064
rect 217506 488280 217562 488336
rect 3330 423580 3332 423600
rect 3332 423580 3384 423600
rect 3384 423580 3386 423600
rect 3330 423544 3386 423580
rect 3330 410488 3386 410544
rect 3330 397432 3386 397488
rect 3330 371320 3386 371376
rect 3330 319232 3386 319288
rect 3330 306176 3386 306232
rect 3330 214920 3386 214976
rect 3054 201864 3110 201920
rect 3698 358400 3754 358456
rect 3606 345344 3662 345400
rect 3514 293120 3570 293176
rect 3514 267144 3570 267200
rect 3514 254088 3570 254144
rect 3514 241032 3570 241088
rect 3514 188808 3570 188864
rect 3514 149776 3570 149832
rect 3514 136720 3570 136776
rect 3514 97552 3570 97608
rect 3514 84632 3570 84688
rect 3514 71576 3570 71632
rect 3514 58520 3570 58576
rect 3422 45464 3478 45520
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 25502 430752 25558 430808
rect 32402 300056 32458 300112
rect 97814 364656 97870 364712
rect 97722 361936 97778 361992
rect 97814 356496 97870 356552
rect 97722 345616 97778 345672
rect 97630 340176 97686 340232
rect 97538 332016 97594 332072
rect 97446 326576 97502 326632
rect 97354 315696 97410 315752
rect 97262 310256 97318 310312
rect 97170 299376 97226 299432
rect 97906 351056 97962 351112
rect 97906 348336 97962 348392
rect 98550 321136 98606 321192
rect 97906 304816 97962 304872
rect 97538 299240 97594 299296
rect 134154 372680 134210 372736
rect 159914 374040 159970 374096
rect 118330 371612 118386 371648
rect 118330 371592 118332 371612
rect 118332 371592 118384 371612
rect 118384 371592 118386 371612
rect 119066 371612 119122 371648
rect 119066 371592 119068 371612
rect 119068 371592 119120 371612
rect 119120 371592 119122 371612
rect 99838 367920 99894 367976
rect 99286 359216 99342 359272
rect 99194 353776 99250 353832
rect 99102 342896 99158 342952
rect 99010 337456 99066 337512
rect 98918 329296 98974 329352
rect 98826 323856 98882 323912
rect 98734 318416 98790 318472
rect 98642 307536 98698 307592
rect 99378 334736 99434 334792
rect 99286 300736 99342 300792
rect 99470 312976 99526 313032
rect 170770 309712 170826 309768
rect 171782 350376 171838 350432
rect 171322 323176 171378 323232
rect 171506 320456 171562 320512
rect 171506 317736 171562 317792
rect 170954 309304 171010 309360
rect 99838 302096 99894 302152
rect 166630 300600 166686 300656
rect 169758 301688 169814 301744
rect 169850 300600 169906 300656
rect 168378 300328 168434 300384
rect 160098 300192 160154 300248
rect 150898 297880 150954 297936
rect 170402 305632 170458 305688
rect 172334 369416 172390 369472
rect 171966 366696 172022 366752
rect 172334 363976 172390 364032
rect 172058 361256 172114 361312
rect 172426 358536 172482 358592
rect 172426 355816 172482 355872
rect 172426 353096 172482 353152
rect 172426 347656 172482 347712
rect 172150 344936 172206 344992
rect 172426 342252 172428 342272
rect 172428 342252 172480 342272
rect 172480 342252 172482 342272
rect 172426 342216 172482 342252
rect 172426 339516 172482 339552
rect 172426 339496 172428 339516
rect 172428 339496 172480 339516
rect 172480 339496 172482 339516
rect 172426 336796 172482 336832
rect 172426 336776 172428 336796
rect 172428 336776 172480 336796
rect 172480 336776 172482 336796
rect 172242 334056 172298 334112
rect 172426 331336 172482 331392
rect 172426 328616 172482 328672
rect 172334 325896 172390 325952
rect 172426 315016 172482 315072
rect 172426 312296 172482 312352
rect 172426 309576 172482 309632
rect 173254 309440 173310 309496
rect 173438 308896 173494 308952
rect 173622 308760 173678 308816
rect 174634 309168 174690 309224
rect 174542 308488 174598 308544
rect 172426 306856 172482 306912
rect 172334 304136 172390 304192
rect 172426 301416 172482 301472
rect 219162 512760 219218 512816
rect 219070 510992 219126 511048
rect 218886 509904 218942 509960
rect 218978 508136 219034 508192
rect 238482 477264 238538 477320
rect 242806 477128 242862 477184
rect 240046 476856 240102 476912
rect 241426 476856 241482 476912
rect 237378 476312 237434 476368
rect 237286 476176 237342 476232
rect 249062 476584 249118 476640
rect 259274 476584 259330 476640
rect 264886 476604 264942 476640
rect 264886 476584 264888 476604
rect 264888 476584 264940 476604
rect 264940 476584 264942 476604
rect 245474 476312 245530 476368
rect 247682 476312 247738 476368
rect 244186 476176 244242 476232
rect 246302 476176 246358 476232
rect 248234 476176 248290 476232
rect 253846 476448 253902 476504
rect 251086 476312 251142 476368
rect 252374 476312 252430 476368
rect 256606 476312 256662 476368
rect 249706 476176 249762 476232
rect 250994 476176 251050 476232
rect 252466 476176 252522 476232
rect 253754 476176 253810 476232
rect 255226 476176 255282 476232
rect 256514 476176 256570 476232
rect 211894 300464 211950 300520
rect 211802 297608 211858 297664
rect 211066 297336 211122 297392
rect 212354 297744 212410 297800
rect 212170 297472 212226 297528
rect 212170 3440 212226 3496
rect 213366 3440 213422 3496
rect 214562 297880 214618 297936
rect 214470 3440 214526 3496
rect 215666 3440 215722 3496
rect 215114 3168 215170 3224
rect 216678 188128 216734 188184
rect 217138 196832 217194 196888
rect 217046 192752 217102 192808
rect 217414 195880 217470 195936
rect 217230 168272 217286 168328
rect 216494 3304 216550 3360
rect 217690 193704 217746 193760
rect 217598 169904 217654 169960
rect 217782 168000 217838 168056
rect 218426 243480 218482 243536
rect 218518 190984 218574 191040
rect 218702 189896 218758 189952
rect 218058 3576 218114 3632
rect 237470 436192 237526 436248
rect 235722 436056 235778 436112
rect 234434 434696 234490 434752
rect 233882 433744 233938 433800
rect 232686 433336 232742 433392
rect 236274 434832 236330 434888
rect 238114 433472 238170 433528
rect 239310 433608 239366 433664
rect 240046 432248 240102 432304
rect 253202 433880 253258 433936
rect 257986 476176 258042 476232
rect 259366 476468 259422 476504
rect 259366 476448 259368 476468
rect 259368 476448 259420 476468
rect 259420 476448 259422 476468
rect 260654 476312 260710 476368
rect 262034 476312 262090 476368
rect 260746 476176 260802 476232
rect 262126 476176 262182 476232
rect 263506 476176 263562 476232
rect 264794 476176 264850 476232
rect 266266 476312 266322 476368
rect 266174 476176 266230 476232
rect 267554 476312 267610 476368
rect 267646 476176 267702 476232
rect 269026 477264 269082 477320
rect 281446 476856 281502 476912
rect 274546 476448 274602 476504
rect 271694 476312 271750 476368
rect 274454 476312 274510 476368
rect 268934 476176 268990 476232
rect 270406 476176 270462 476232
rect 271786 476176 271842 476232
rect 273166 476176 273222 476232
rect 274362 476176 274418 476232
rect 237286 432112 237342 432168
rect 235446 431976 235502 432032
rect 277306 476312 277362 476368
rect 278594 476312 278650 476368
rect 275926 476176 275982 476232
rect 277214 476176 277270 476232
rect 278686 476176 278742 476232
rect 280066 476176 280122 476232
rect 284206 476176 284262 476232
rect 286966 476176 287022 476232
rect 288346 476176 288402 476232
rect 291106 476176 291162 476232
rect 293866 476176 293922 476232
rect 296626 476176 296682 476232
rect 299386 476176 299442 476232
rect 302146 476176 302202 476232
rect 294694 435240 294750 435296
rect 296442 434968 296498 435024
rect 300122 435104 300178 435160
rect 298926 433880 298982 433936
rect 306102 476992 306158 477048
rect 309046 476720 309102 476776
rect 303526 476332 303582 476368
rect 303526 476312 303528 476332
rect 303528 476312 303580 476332
rect 303580 476312 303582 476332
rect 321466 476992 321522 477048
rect 311806 476176 311862 476232
rect 314566 476584 314622 476640
rect 315946 476176 316002 476232
rect 318706 476448 318762 476504
rect 324226 476312 324282 476368
rect 326986 476176 327042 476232
rect 580170 697176 580226 697232
rect 580262 683848 580318 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 579986 630808 580042 630864
rect 580170 617480 580226 617536
rect 580170 590960 580226 591016
rect 580170 577632 580226 577688
rect 580170 564304 580226 564360
rect 579894 537784 579950 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 578882 511264 578938 511320
rect 580170 484608 580226 484664
rect 580170 471416 580226 471472
rect 580170 458088 580226 458144
rect 243358 431704 243414 431760
rect 299478 431704 299534 431760
rect 226982 310528 227038 310584
rect 230018 309712 230074 309768
rect 229926 309032 229982 309088
rect 231214 310256 231270 310312
rect 231490 370232 231546 370288
rect 231858 310392 231914 310448
rect 231490 308624 231546 308680
rect 231306 308352 231362 308408
rect 232778 310528 232834 310584
rect 232226 310412 232282 310448
rect 232226 310392 232228 310412
rect 232228 310392 232280 310412
rect 232280 310392 232282 310412
rect 234342 309032 234398 309088
rect 233330 299240 233386 299296
rect 234986 310256 235042 310312
rect 235354 309032 235410 309088
rect 236458 299376 236514 299432
rect 239034 301144 239090 301200
rect 239402 308624 239458 308680
rect 239402 308352 239458 308408
rect 240506 309576 240562 309632
rect 242438 308216 242494 308272
rect 243358 308760 243414 308816
rect 245290 309440 245346 309496
rect 245474 309304 245530 309360
rect 246210 309848 246266 309904
rect 244646 300736 244702 300792
rect 246854 309712 246910 309768
rect 247038 308896 247094 308952
rect 250258 309168 250314 309224
rect 249982 301552 250038 301608
rect 250810 308488 250866 308544
rect 251178 308624 251234 308680
rect 253478 305632 253534 305688
rect 255870 300056 255926 300112
rect 270038 300192 270094 300248
rect 276478 300328 276534 300384
rect 281998 265512 282054 265568
rect 284298 306040 284354 306096
rect 284114 303184 284170 303240
rect 284850 306176 284906 306232
rect 285034 303320 285090 303376
rect 284666 303048 284722 303104
rect 284482 302912 284538 302968
rect 285862 305768 285918 305824
rect 283378 301688 283434 301744
rect 286966 305904 287022 305960
rect 286138 300464 286194 300520
rect 288714 302776 288770 302832
rect 288622 301416 288678 301472
rect 287610 297880 287666 297936
rect 287518 297744 287574 297800
rect 287426 297608 287482 297664
rect 289266 297472 289322 297528
rect 288898 297336 288954 297392
rect 283194 293120 283250 293176
rect 283102 284824 283158 284880
rect 282918 262792 282974 262848
rect 294326 302776 294382 302832
rect 294234 300464 294290 300520
rect 294694 300328 294750 300384
rect 295062 305632 295118 305688
rect 294786 300192 294842 300248
rect 298466 308624 298522 308680
rect 298834 308352 298890 308408
rect 296994 247968 297050 248024
rect 299662 308488 299718 308544
rect 298190 248104 298246 248160
rect 302238 245384 302294 245440
rect 303986 308760 304042 308816
rect 302698 250552 302754 250608
rect 302882 250416 302938 250472
rect 303894 250824 303950 250880
rect 305642 302912 305698 302968
rect 305550 300600 305606 300656
rect 305458 295976 305514 296032
rect 305366 294480 305422 294536
rect 305274 283464 305330 283520
rect 305182 280744 305238 280800
rect 305090 267008 305146 267064
rect 304998 265512 305054 265568
rect 306654 306312 306710 306368
rect 306470 306040 306526 306096
rect 306654 272448 306710 272504
rect 306470 262792 306526 262848
rect 304078 250688 304134 250744
rect 303710 248240 303766 248296
rect 303618 246200 303674 246256
rect 302422 245520 302478 245576
rect 322110 300056 322166 300112
rect 320178 245248 320234 245304
rect 323030 247832 323086 247888
rect 322938 245112 322994 245168
rect 328458 247696 328514 247752
rect 323122 244976 323178 245032
rect 333150 306448 333206 306504
rect 333058 306176 333114 306232
rect 334162 247560 334218 247616
rect 336922 306312 336978 306368
rect 338670 309032 338726 309088
rect 338486 308216 338542 308272
rect 338854 303048 338910 303104
rect 339222 308896 339278 308952
rect 340142 306312 340198 306368
rect 339498 303184 339554 303240
rect 340786 306040 340842 306096
rect 341522 305904 341578 305960
rect 343730 306176 343786 306232
rect 344926 303456 344982 303512
rect 345202 303320 345258 303376
rect 357898 433744 357954 433800
rect 355414 308624 355470 308680
rect 332598 244840 332654 244896
rect 295430 243480 295486 243536
rect 238206 159840 238262 159896
rect 239586 159840 239642 159896
rect 241702 159840 241758 159896
rect 255962 159568 256018 159624
rect 220818 158616 220874 158672
rect 219438 157800 219494 157856
rect 224958 158480 225014 158536
rect 223578 158344 223634 158400
rect 219254 3712 219310 3768
rect 219346 3576 219402 3632
rect 219254 3440 219310 3496
rect 222750 3848 222806 3904
rect 231858 158208 231914 158264
rect 226338 3576 226394 3632
rect 227534 3168 227590 3224
rect 240506 158616 240562 158672
rect 248326 158652 248328 158672
rect 248328 158652 248380 158672
rect 248380 158652 248382 158672
rect 248326 158616 248382 158652
rect 250166 158616 250222 158672
rect 251454 158616 251510 158672
rect 254582 158616 254638 158672
rect 238758 158072 238814 158128
rect 240506 3304 240562 3360
rect 251086 158072 251142 158128
rect 251178 157936 251234 157992
rect 256054 158636 256110 158672
rect 256054 158616 256056 158636
rect 256056 158616 256108 158636
rect 256108 158616 256110 158636
rect 252374 157936 252430 157992
rect 251270 155216 251326 155272
rect 253570 157936 253626 157992
rect 253662 157392 253718 157448
rect 273626 159840 273682 159896
rect 276110 159840 276166 159896
rect 278502 159840 278558 159896
rect 293498 159840 293554 159896
rect 295890 159840 295946 159896
rect 303526 159840 303582 159896
rect 310978 159840 311034 159896
rect 313462 159840 313518 159896
rect 257158 158616 257214 158672
rect 258262 158616 258318 158672
rect 258630 158616 258686 158672
rect 259550 158616 259606 158672
rect 261206 158616 261262 158672
rect 262862 158616 262918 158672
rect 263966 158616 264022 158672
rect 263966 157392 264022 157448
rect 265346 159568 265402 159624
rect 265990 158616 266046 158672
rect 266818 158616 266874 158672
rect 267646 158616 267702 158672
rect 268750 158616 268806 158672
rect 268934 157936 268990 157992
rect 271050 159568 271106 159624
rect 269854 158616 269910 158672
rect 271142 158616 271198 158672
rect 272246 158616 272302 158672
rect 274178 158616 274234 158672
rect 274454 158616 274510 158672
rect 275926 158616 275982 158672
rect 277122 158072 277178 158128
rect 278134 158072 278190 158128
rect 281078 158616 281134 158672
rect 279974 158072 280030 158128
rect 298466 159704 298522 159760
rect 291014 158616 291070 158672
rect 300950 158616 301006 158672
rect 308678 158616 308734 158672
rect 321098 158616 321154 158672
rect 323398 158616 323454 158672
rect 325974 158616 326030 158672
rect 283746 157800 283802 157856
rect 286506 157800 286562 157856
rect 353942 158072 353998 158128
rect 288254 157392 288310 157448
rect 306102 157392 306158 157448
rect 315854 157392 315910 157448
rect 318614 157392 318670 157448
rect 305550 8880 305606 8936
rect 319718 9016 319774 9072
rect 348054 6704 348110 6760
rect 344558 6568 344614 6624
rect 340970 6432 341026 6488
rect 337474 6296 337530 6352
rect 333886 6160 333942 6216
rect 338670 3440 338726 3496
rect 339866 3304 339922 3360
rect 342166 3712 342222 3768
rect 343362 3576 343418 3632
rect 346950 3984 347006 4040
rect 345754 3848 345810 3904
rect 351642 6840 351698 6896
rect 354126 157936 354182 157992
rect 357530 308488 357586 308544
rect 356702 3576 356758 3632
rect 352838 3168 352894 3224
rect 357990 305632 358046 305688
rect 357898 244296 357954 244352
rect 358082 205536 358138 205592
rect 358266 300464 358322 300520
rect 358082 158072 358138 158128
rect 358358 157936 358414 157992
rect 360198 308760 360254 308816
rect 359554 308216 359610 308272
rect 356702 3032 356758 3088
rect 359094 3576 359150 3632
rect 359554 158480 359610 158536
rect 359922 3440 359978 3496
rect 360382 3984 360438 4040
rect 360934 157392 360990 157448
rect 360566 3304 360622 3360
rect 360198 3168 360254 3224
rect 362222 309032 362278 309088
rect 361118 3440 361174 3496
rect 362314 308896 362370 308952
rect 362222 158208 362278 158264
rect 362498 308352 362554 308408
rect 362406 306312 362462 306368
rect 362314 157528 362370 157584
rect 362222 157392 362278 157448
rect 361762 3032 361818 3088
rect 362498 156984 362554 157040
rect 363050 6296 363106 6352
rect 362958 6160 363014 6216
rect 363234 6432 363290 6488
rect 363694 303456 363750 303512
rect 363786 302776 363842 302832
rect 365166 303048 365222 303104
rect 364982 159024 365038 159080
rect 364890 158888 364946 158944
rect 364798 158752 364854 158808
rect 365994 306040 366050 306096
rect 365994 157120 366050 157176
rect 366454 303184 366510 303240
rect 366546 300328 366602 300384
rect 368662 306176 368718 306232
rect 367926 303320 367982 303376
rect 368754 305904 368810 305960
rect 378782 305768 378838 305824
rect 368754 157256 368810 157312
rect 368938 158344 368994 158400
rect 369398 158752 369454 158808
rect 367006 3848 367062 3904
rect 362314 3440 362370 3496
rect 363510 3440 363566 3496
rect 364614 3440 364670 3496
rect 365810 3440 365866 3496
rect 368202 3440 368258 3496
rect 369398 3440 369454 3496
rect 370410 300192 370466 300248
rect 370594 3440 370650 3496
rect 467102 300056 467158 300112
rect 467838 245248 467894 245304
rect 480258 245112 480314 245168
rect 483018 247832 483074 247888
rect 481730 244976 481786 245032
rect 520278 247696 520334 247752
rect 545118 244840 545174 244896
rect 557538 247560 557594 247616
rect 579986 433608 580042 433664
rect 579894 431568 579950 431624
rect 577594 430616 577650 430672
rect 580446 433472 580502 433528
rect 580262 433336 580318 433392
rect 579986 418240 580042 418296
rect 579986 404912 580042 404968
rect 580078 378392 580134 378448
rect 580170 365064 580226 365120
rect 580170 351872 580226 351928
rect 580170 325216 580226 325272
rect 580170 298696 580226 298752
rect 579986 272176 580042 272232
rect 579802 258848 579858 258904
rect 580170 245520 580226 245576
rect 579710 219000 579766 219056
rect 579618 205672 579674 205728
rect 579710 179152 579766 179208
rect 580538 152632 580594 152688
rect 580906 312024 580962 312080
rect 580814 232328 580870 232384
rect 580722 192480 580778 192536
rect 580630 139304 580686 139360
rect 580446 125976 580502 126032
rect 580354 33088 580410 33144
rect 580262 6568 580318 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580257 683906 580323 683909
rect 583520 683906 584960 683996
rect 580257 683904 584960 683906
rect 580257 683848 580262 683904
rect 580318 683848 584960 683904
rect 580257 683846 584960 683848
rect 580257 683843 580323 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 579981 630866 580047 630869
rect 583520 630866 584960 630956
rect 579981 630864 584960 630866
rect 579981 630808 579986 630864
rect 580042 630808 584960 630864
rect 579981 630806 584960 630808
rect 579981 630803 580047 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3417 606114 3483 606117
rect -960 606112 3483 606114
rect -960 606056 3422 606112
rect 3478 606056 3483 606112
rect -960 606054 3483 606056
rect -960 605964 480 606054
rect 3417 606051 3483 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 579889 537842 579955 537845
rect 583520 537842 584960 537932
rect 579889 537840 584960 537842
rect 579889 537784 579894 537840
rect 579950 537784 584960 537840
rect 579889 537782 584960 537784
rect 579889 537779 579955 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 2773 527914 2839 527917
rect -960 527912 2839 527914
rect -960 527856 2778 527912
rect 2834 527856 2839 527912
rect -960 527854 2839 527856
rect -960 527764 480 527854
rect 2773 527851 2839 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect 217777 516898 217843 516901
rect 219390 516898 220064 516924
rect 217777 516896 220064 516898
rect 217777 516840 217782 516896
rect 217838 516864 220064 516896
rect 217838 516840 219450 516864
rect 217777 516838 219450 516840
rect 217777 516835 217843 516838
rect 217685 515946 217751 515949
rect 219390 515946 220064 515972
rect 217685 515944 220064 515946
rect 217685 515888 217690 515944
rect 217746 515912 220064 515944
rect 217746 515888 219450 515912
rect 217685 515886 219450 515888
rect 217685 515883 217751 515886
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 217593 513770 217659 513773
rect 219390 513770 220064 513796
rect 217593 513768 220064 513770
rect 217593 513712 217598 513768
rect 217654 513736 220064 513768
rect 217654 513712 219450 513736
rect 217593 513710 219450 513712
rect 217593 513707 217659 513710
rect 219157 512818 219223 512821
rect 219390 512818 220064 512844
rect 219157 512816 220064 512818
rect 219157 512760 219162 512816
rect 219218 512784 220064 512816
rect 219218 512760 219450 512784
rect 219157 512758 219450 512760
rect 219157 512755 219223 512758
rect 578877 511322 578943 511325
rect 583520 511322 584960 511412
rect 578877 511320 584960 511322
rect 578877 511264 578882 511320
rect 578938 511264 584960 511320
rect 578877 511262 584960 511264
rect 578877 511259 578943 511262
rect 583520 511172 584960 511262
rect 219065 511050 219131 511053
rect 219390 511050 220064 511076
rect 219065 511048 220064 511050
rect 219065 510992 219070 511048
rect 219126 511016 220064 511048
rect 219126 510992 219450 511016
rect 219065 510990 219450 510992
rect 219065 510987 219131 510990
rect 218881 509962 218947 509965
rect 219390 509962 220064 509988
rect 218881 509960 220064 509962
rect 218881 509904 218886 509960
rect 218942 509928 220064 509960
rect 218942 509904 219450 509928
rect 218881 509902 219450 509904
rect 218881 509899 218947 509902
rect 218973 508194 219039 508197
rect 219390 508194 220064 508220
rect 218973 508192 220064 508194
rect 218973 508136 218978 508192
rect 219034 508160 220064 508192
rect 219034 508136 219450 508160
rect 218973 508134 219450 508136
rect 218973 508131 219039 508134
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 583520 497844 584960 498084
rect 217409 489970 217475 489973
rect 219390 489970 220064 489996
rect 217409 489968 220064 489970
rect 217409 489912 217414 489968
rect 217470 489936 220064 489968
rect 217470 489912 219450 489936
rect 217409 489910 219450 489912
rect 217409 489907 217475 489910
rect -960 488596 480 488836
rect 217501 488338 217567 488341
rect 219390 488338 220064 488364
rect 217501 488336 220064 488338
rect 217501 488280 217506 488336
rect 217562 488304 220064 488336
rect 217562 488280 219450 488304
rect 217501 488278 219450 488280
rect 217501 488275 217567 488278
rect 217317 488066 217383 488069
rect 219390 488066 220064 488092
rect 217317 488064 220064 488066
rect 217317 488008 217322 488064
rect 217378 488032 220064 488064
rect 217378 488008 219450 488032
rect 217317 488006 219450 488008
rect 217317 488003 217383 488006
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect 238334 477260 238340 477324
rect 238404 477322 238410 477324
rect 238477 477322 238543 477325
rect 238404 477320 238543 477322
rect 238404 477264 238482 477320
rect 238538 477264 238543 477320
rect 238404 477262 238543 477264
rect 238404 477260 238410 477262
rect 238477 477259 238543 477262
rect 268326 477260 268332 477324
rect 268396 477322 268402 477324
rect 269021 477322 269087 477325
rect 268396 477320 269087 477322
rect 268396 477264 269026 477320
rect 269082 477264 269087 477320
rect 268396 477262 269087 477264
rect 268396 477260 268402 477262
rect 269021 477259 269087 477262
rect 241830 477124 241836 477188
rect 241900 477186 241906 477188
rect 242801 477186 242867 477189
rect 241900 477184 242867 477186
rect 241900 477128 242806 477184
rect 242862 477128 242867 477184
rect 241900 477126 242867 477128
rect 241900 477124 241906 477126
rect 242801 477123 242867 477126
rect 306097 477052 306163 477053
rect 306046 476988 306052 477052
rect 306116 477050 306163 477052
rect 306116 477048 306208 477050
rect 306158 476992 306208 477048
rect 306116 476990 306208 476992
rect 306116 476988 306163 476990
rect 320950 476988 320956 477052
rect 321020 477050 321026 477052
rect 321461 477050 321527 477053
rect 321020 477048 321527 477050
rect 321020 476992 321466 477048
rect 321522 476992 321527 477048
rect 321020 476990 321527 476992
rect 321020 476988 321026 476990
rect 306097 476987 306163 476988
rect 321461 476987 321527 476990
rect 239622 476852 239628 476916
rect 239692 476914 239698 476916
rect 240041 476914 240107 476917
rect 239692 476912 240107 476914
rect 239692 476856 240046 476912
rect 240102 476856 240107 476912
rect 239692 476854 240107 476856
rect 239692 476852 239698 476854
rect 240041 476851 240107 476854
rect 240542 476852 240548 476916
rect 240612 476914 240618 476916
rect 241421 476914 241487 476917
rect 240612 476912 241487 476914
rect 240612 476856 241426 476912
rect 241482 476856 241487 476912
rect 240612 476854 241487 476856
rect 240612 476852 240618 476854
rect 241421 476851 241487 476854
rect 281022 476852 281028 476916
rect 281092 476914 281098 476916
rect 281441 476914 281507 476917
rect 281092 476912 281507 476914
rect 281092 476856 281446 476912
rect 281502 476856 281507 476912
rect 281092 476854 281507 476856
rect 281092 476852 281098 476854
rect 281441 476851 281507 476854
rect 308622 476716 308628 476780
rect 308692 476778 308698 476780
rect 309041 476778 309107 476781
rect 308692 476776 309107 476778
rect 308692 476720 309046 476776
rect 309102 476720 309107 476776
rect 308692 476718 309107 476720
rect 308692 476716 308698 476718
rect 309041 476715 309107 476718
rect 248270 476580 248276 476644
rect 248340 476642 248346 476644
rect 249057 476642 249123 476645
rect 248340 476640 249123 476642
rect 248340 476584 249062 476640
rect 249118 476584 249123 476640
rect 248340 476582 249123 476584
rect 248340 476580 248346 476582
rect 249057 476579 249123 476582
rect 258022 476580 258028 476644
rect 258092 476642 258098 476644
rect 259269 476642 259335 476645
rect 258092 476640 259335 476642
rect 258092 476584 259274 476640
rect 259330 476584 259335 476640
rect 258092 476582 259335 476584
rect 258092 476580 258098 476582
rect 259269 476579 259335 476582
rect 263542 476580 263548 476644
rect 263612 476642 263618 476644
rect 264881 476642 264947 476645
rect 263612 476640 264947 476642
rect 263612 476584 264886 476640
rect 264942 476584 264947 476640
rect 263612 476582 264947 476584
rect 263612 476580 263618 476582
rect 264881 476579 264947 476582
rect 313406 476580 313412 476644
rect 313476 476642 313482 476644
rect 314561 476642 314627 476645
rect 313476 476640 314627 476642
rect 313476 476584 314566 476640
rect 314622 476584 314627 476640
rect 313476 476582 314627 476584
rect 313476 476580 313482 476582
rect 314561 476579 314627 476582
rect 253606 476444 253612 476508
rect 253676 476506 253682 476508
rect 253841 476506 253907 476509
rect 253676 476504 253907 476506
rect 253676 476448 253846 476504
rect 253902 476448 253907 476504
rect 253676 476446 253907 476448
rect 253676 476444 253682 476446
rect 253841 476443 253907 476446
rect 259126 476444 259132 476508
rect 259196 476506 259202 476508
rect 259361 476506 259427 476509
rect 259196 476504 259427 476506
rect 259196 476448 259366 476504
rect 259422 476448 259427 476504
rect 259196 476446 259427 476448
rect 259196 476444 259202 476446
rect 259361 476443 259427 476446
rect 273662 476444 273668 476508
rect 273732 476506 273738 476508
rect 274541 476506 274607 476509
rect 273732 476504 274607 476506
rect 273732 476448 274546 476504
rect 274602 476448 274607 476504
rect 273732 476446 274607 476448
rect 273732 476444 273738 476446
rect 274541 476443 274607 476446
rect 318558 476444 318564 476508
rect 318628 476506 318634 476508
rect 318701 476506 318767 476509
rect 318628 476504 318767 476506
rect 318628 476448 318706 476504
rect 318762 476448 318767 476504
rect 318628 476446 318767 476448
rect 318628 476444 318634 476446
rect 318701 476443 318767 476446
rect 236126 476308 236132 476372
rect 236196 476370 236202 476372
rect 237373 476370 237439 476373
rect 236196 476368 237439 476370
rect 236196 476312 237378 476368
rect 237434 476312 237439 476368
rect 236196 476310 237439 476312
rect 236196 476308 236202 476310
rect 237373 476307 237439 476310
rect 244222 476308 244228 476372
rect 244292 476370 244298 476372
rect 245469 476370 245535 476373
rect 244292 476368 245535 476370
rect 244292 476312 245474 476368
rect 245530 476312 245535 476368
rect 244292 476310 245535 476312
rect 244292 476308 244298 476310
rect 245469 476307 245535 476310
rect 246614 476308 246620 476372
rect 246684 476370 246690 476372
rect 247677 476370 247743 476373
rect 246684 476368 247743 476370
rect 246684 476312 247682 476368
rect 247738 476312 247743 476368
rect 246684 476310 247743 476312
rect 246684 476308 246690 476310
rect 247677 476307 247743 476310
rect 250110 476308 250116 476372
rect 250180 476370 250186 476372
rect 251081 476370 251147 476373
rect 250180 476368 251147 476370
rect 250180 476312 251086 476368
rect 251142 476312 251147 476368
rect 250180 476310 251147 476312
rect 250180 476308 250186 476310
rect 251081 476307 251147 476310
rect 251398 476308 251404 476372
rect 251468 476370 251474 476372
rect 252369 476370 252435 476373
rect 251468 476368 252435 476370
rect 251468 476312 252374 476368
rect 252430 476312 252435 476368
rect 251468 476310 252435 476312
rect 251468 476308 251474 476310
rect 252369 476307 252435 476310
rect 255814 476308 255820 476372
rect 255884 476370 255890 476372
rect 256601 476370 256667 476373
rect 255884 476368 256667 476370
rect 255884 476312 256606 476368
rect 256662 476312 256667 476368
rect 255884 476310 256667 476312
rect 255884 476308 255890 476310
rect 256601 476307 256667 476310
rect 259494 476308 259500 476372
rect 259564 476370 259570 476372
rect 260649 476370 260715 476373
rect 259564 476368 260715 476370
rect 259564 476312 260654 476368
rect 260710 476312 260715 476368
rect 259564 476310 260715 476312
rect 259564 476308 259570 476310
rect 260649 476307 260715 476310
rect 261150 476308 261156 476372
rect 261220 476370 261226 476372
rect 262029 476370 262095 476373
rect 261220 476368 262095 476370
rect 261220 476312 262034 476368
rect 262090 476312 262095 476368
rect 261220 476310 262095 476312
rect 261220 476308 261226 476310
rect 262029 476307 262095 476310
rect 265382 476308 265388 476372
rect 265452 476370 265458 476372
rect 266261 476370 266327 476373
rect 265452 476368 266327 476370
rect 265452 476312 266266 476368
rect 266322 476312 266327 476368
rect 265452 476310 266327 476312
rect 265452 476308 265458 476310
rect 266261 476307 266327 476310
rect 266486 476308 266492 476372
rect 266556 476370 266562 476372
rect 267549 476370 267615 476373
rect 266556 476368 267615 476370
rect 266556 476312 267554 476368
rect 267610 476312 267615 476368
rect 266556 476310 267615 476312
rect 266556 476308 266562 476310
rect 267549 476307 267615 476310
rect 270902 476308 270908 476372
rect 270972 476370 270978 476372
rect 271689 476370 271755 476373
rect 270972 476368 271755 476370
rect 270972 476312 271694 476368
rect 271750 476312 271755 476368
rect 270972 476310 271755 476312
rect 270972 476308 270978 476310
rect 271689 476307 271755 476310
rect 273294 476308 273300 476372
rect 273364 476370 273370 476372
rect 274449 476370 274515 476373
rect 273364 476368 274515 476370
rect 273364 476312 274454 476368
rect 274510 476312 274515 476368
rect 273364 476310 274515 476312
rect 273364 476308 273370 476310
rect 274449 476307 274515 476310
rect 276054 476308 276060 476372
rect 276124 476370 276130 476372
rect 277301 476370 277367 476373
rect 276124 476368 277367 476370
rect 276124 476312 277306 476368
rect 277362 476312 277367 476368
rect 276124 476310 277367 476312
rect 276124 476308 276130 476310
rect 277301 476307 277367 476310
rect 278078 476308 278084 476372
rect 278148 476370 278154 476372
rect 278589 476370 278655 476373
rect 303521 476372 303587 476373
rect 278148 476368 278655 476370
rect 278148 476312 278594 476368
rect 278650 476312 278655 476368
rect 278148 476310 278655 476312
rect 278148 476308 278154 476310
rect 278589 476307 278655 476310
rect 303470 476308 303476 476372
rect 303540 476370 303587 476372
rect 303540 476368 303632 476370
rect 303582 476312 303632 476368
rect 303540 476310 303632 476312
rect 303540 476308 303587 476310
rect 323342 476308 323348 476372
rect 323412 476370 323418 476372
rect 324221 476370 324287 476373
rect 323412 476368 324287 476370
rect 323412 476312 324226 476368
rect 324282 476312 324287 476368
rect 323412 476310 324287 476312
rect 323412 476308 323418 476310
rect 303521 476307 303587 476308
rect 324221 476307 324287 476310
rect 237281 476236 237347 476237
rect 237230 476172 237236 476236
rect 237300 476234 237347 476236
rect 237300 476232 237392 476234
rect 237342 476176 237392 476232
rect 237300 476174 237392 476176
rect 237300 476172 237347 476174
rect 243118 476172 243124 476236
rect 243188 476234 243194 476236
rect 244181 476234 244247 476237
rect 243188 476232 244247 476234
rect 243188 476176 244186 476232
rect 244242 476176 244247 476232
rect 243188 476174 244247 476176
rect 243188 476172 243194 476174
rect 237281 476171 237347 476172
rect 244181 476171 244247 476174
rect 245510 476172 245516 476236
rect 245580 476234 245586 476236
rect 246297 476234 246363 476237
rect 245580 476232 246363 476234
rect 245580 476176 246302 476232
rect 246358 476176 246363 476232
rect 245580 476174 246363 476176
rect 245580 476172 245586 476174
rect 246297 476171 246363 476174
rect 247718 476172 247724 476236
rect 247788 476234 247794 476236
rect 248229 476234 248295 476237
rect 247788 476232 248295 476234
rect 247788 476176 248234 476232
rect 248290 476176 248295 476232
rect 247788 476174 248295 476176
rect 247788 476172 247794 476174
rect 248229 476171 248295 476174
rect 248638 476172 248644 476236
rect 248708 476234 248714 476236
rect 249701 476234 249767 476237
rect 248708 476232 249767 476234
rect 248708 476176 249706 476232
rect 249762 476176 249767 476232
rect 248708 476174 249767 476176
rect 248708 476172 248714 476174
rect 249701 476171 249767 476174
rect 250846 476172 250852 476236
rect 250916 476234 250922 476236
rect 250989 476234 251055 476237
rect 250916 476232 251055 476234
rect 250916 476176 250994 476232
rect 251050 476176 251055 476232
rect 250916 476174 251055 476176
rect 250916 476172 250922 476174
rect 250989 476171 251055 476174
rect 252318 476172 252324 476236
rect 252388 476234 252394 476236
rect 252461 476234 252527 476237
rect 252388 476232 252527 476234
rect 252388 476176 252466 476232
rect 252522 476176 252527 476232
rect 252388 476174 252527 476176
rect 252388 476172 252394 476174
rect 252461 476171 252527 476174
rect 253422 476172 253428 476236
rect 253492 476234 253498 476236
rect 253749 476234 253815 476237
rect 253492 476232 253815 476234
rect 253492 476176 253754 476232
rect 253810 476176 253815 476232
rect 253492 476174 253815 476176
rect 253492 476172 253498 476174
rect 253749 476171 253815 476174
rect 254526 476172 254532 476236
rect 254596 476234 254602 476236
rect 255221 476234 255287 476237
rect 254596 476232 255287 476234
rect 254596 476176 255226 476232
rect 255282 476176 255287 476232
rect 254596 476174 255287 476176
rect 254596 476172 254602 476174
rect 255221 476171 255287 476174
rect 256182 476172 256188 476236
rect 256252 476234 256258 476236
rect 256509 476234 256575 476237
rect 256252 476232 256575 476234
rect 256252 476176 256514 476232
rect 256570 476176 256575 476232
rect 256252 476174 256575 476176
rect 256252 476172 256258 476174
rect 256509 476171 256575 476174
rect 257102 476172 257108 476236
rect 257172 476234 257178 476236
rect 257981 476234 258047 476237
rect 257172 476232 258047 476234
rect 257172 476176 257986 476232
rect 258042 476176 258047 476232
rect 257172 476174 258047 476176
rect 257172 476172 257178 476174
rect 257981 476171 258047 476174
rect 260598 476172 260604 476236
rect 260668 476234 260674 476236
rect 260741 476234 260807 476237
rect 260668 476232 260807 476234
rect 260668 476176 260746 476232
rect 260802 476176 260807 476232
rect 260668 476174 260807 476176
rect 260668 476172 260674 476174
rect 260741 476171 260807 476174
rect 261702 476172 261708 476236
rect 261772 476234 261778 476236
rect 262121 476234 262187 476237
rect 261772 476232 262187 476234
rect 261772 476176 262126 476232
rect 262182 476176 262187 476232
rect 261772 476174 262187 476176
rect 261772 476172 261778 476174
rect 262121 476171 262187 476174
rect 262806 476172 262812 476236
rect 262876 476234 262882 476236
rect 263501 476234 263567 476237
rect 262876 476232 263567 476234
rect 262876 476176 263506 476232
rect 263562 476176 263567 476232
rect 262876 476174 263567 476176
rect 262876 476172 262882 476174
rect 263501 476171 263567 476174
rect 263910 476172 263916 476236
rect 263980 476234 263986 476236
rect 264789 476234 264855 476237
rect 263980 476232 264855 476234
rect 263980 476176 264794 476232
rect 264850 476176 264855 476232
rect 263980 476174 264855 476176
rect 263980 476172 263986 476174
rect 264789 476171 264855 476174
rect 265934 476172 265940 476236
rect 266004 476234 266010 476236
rect 266169 476234 266235 476237
rect 267641 476236 267707 476237
rect 267590 476234 267596 476236
rect 266004 476232 266235 476234
rect 266004 476176 266174 476232
rect 266230 476176 266235 476232
rect 266004 476174 266235 476176
rect 267550 476174 267596 476234
rect 267660 476232 267707 476236
rect 267702 476176 267707 476232
rect 266004 476172 266010 476174
rect 266169 476171 266235 476174
rect 267590 476172 267596 476174
rect 267660 476172 267707 476176
rect 268694 476172 268700 476236
rect 268764 476234 268770 476236
rect 268929 476234 268995 476237
rect 268764 476232 268995 476234
rect 268764 476176 268934 476232
rect 268990 476176 268995 476232
rect 268764 476174 268995 476176
rect 268764 476172 268770 476174
rect 267641 476171 267707 476172
rect 268929 476171 268995 476174
rect 269798 476172 269804 476236
rect 269868 476234 269874 476236
rect 270401 476234 270467 476237
rect 269868 476232 270467 476234
rect 269868 476176 270406 476232
rect 270462 476176 270467 476232
rect 269868 476174 270467 476176
rect 269868 476172 269874 476174
rect 270401 476171 270467 476174
rect 271270 476172 271276 476236
rect 271340 476234 271346 476236
rect 271781 476234 271847 476237
rect 271340 476232 271847 476234
rect 271340 476176 271786 476232
rect 271842 476176 271847 476232
rect 271340 476174 271847 476176
rect 271340 476172 271346 476174
rect 271781 476171 271847 476174
rect 272190 476172 272196 476236
rect 272260 476234 272266 476236
rect 273161 476234 273227 476237
rect 274357 476236 274423 476237
rect 275921 476236 275987 476237
rect 274357 476234 274404 476236
rect 272260 476232 273227 476234
rect 272260 476176 273166 476232
rect 273222 476176 273227 476232
rect 272260 476174 273227 476176
rect 274312 476232 274404 476234
rect 274312 476176 274362 476232
rect 274312 476174 274404 476176
rect 272260 476172 272266 476174
rect 273161 476171 273227 476174
rect 274357 476172 274404 476174
rect 274468 476172 274474 476236
rect 275870 476172 275876 476236
rect 275940 476234 275987 476236
rect 275940 476232 276032 476234
rect 275982 476176 276032 476232
rect 275940 476174 276032 476176
rect 275940 476172 275987 476174
rect 276974 476172 276980 476236
rect 277044 476234 277050 476236
rect 277209 476234 277275 476237
rect 277044 476232 277275 476234
rect 277044 476176 277214 476232
rect 277270 476176 277275 476232
rect 277044 476174 277275 476176
rect 277044 476172 277050 476174
rect 274357 476171 274423 476172
rect 275921 476171 275987 476172
rect 277209 476171 277275 476174
rect 278446 476172 278452 476236
rect 278516 476234 278522 476236
rect 278681 476234 278747 476237
rect 278516 476232 278747 476234
rect 278516 476176 278686 476232
rect 278742 476176 278747 476232
rect 278516 476174 278747 476176
rect 278516 476172 278522 476174
rect 278681 476171 278747 476174
rect 279182 476172 279188 476236
rect 279252 476234 279258 476236
rect 280061 476234 280127 476237
rect 279252 476232 280127 476234
rect 279252 476176 280066 476232
rect 280122 476176 280127 476232
rect 279252 476174 280127 476176
rect 279252 476172 279258 476174
rect 280061 476171 280127 476174
rect 283598 476172 283604 476236
rect 283668 476234 283674 476236
rect 284201 476234 284267 476237
rect 283668 476232 284267 476234
rect 283668 476176 284206 476232
rect 284262 476176 284267 476232
rect 283668 476174 284267 476176
rect 283668 476172 283674 476174
rect 284201 476171 284267 476174
rect 285990 476172 285996 476236
rect 286060 476234 286066 476236
rect 286961 476234 287027 476237
rect 286060 476232 287027 476234
rect 286060 476176 286966 476232
rect 287022 476176 287027 476232
rect 286060 476174 287027 476176
rect 286060 476172 286066 476174
rect 286961 476171 287027 476174
rect 288198 476172 288204 476236
rect 288268 476234 288274 476236
rect 288341 476234 288407 476237
rect 288268 476232 288407 476234
rect 288268 476176 288346 476232
rect 288402 476176 288407 476232
rect 288268 476174 288407 476176
rect 288268 476172 288274 476174
rect 288341 476171 288407 476174
rect 290958 476172 290964 476236
rect 291028 476234 291034 476236
rect 291101 476234 291167 476237
rect 291028 476232 291167 476234
rect 291028 476176 291106 476232
rect 291162 476176 291167 476232
rect 291028 476174 291167 476176
rect 291028 476172 291034 476174
rect 291101 476171 291167 476174
rect 293534 476172 293540 476236
rect 293604 476234 293610 476236
rect 293861 476234 293927 476237
rect 293604 476232 293927 476234
rect 293604 476176 293866 476232
rect 293922 476176 293927 476232
rect 293604 476174 293927 476176
rect 293604 476172 293610 476174
rect 293861 476171 293927 476174
rect 295926 476172 295932 476236
rect 295996 476234 296002 476236
rect 296621 476234 296687 476237
rect 295996 476232 296687 476234
rect 295996 476176 296626 476232
rect 296682 476176 296687 476232
rect 295996 476174 296687 476176
rect 295996 476172 296002 476174
rect 296621 476171 296687 476174
rect 298502 476172 298508 476236
rect 298572 476234 298578 476236
rect 299381 476234 299447 476237
rect 298572 476232 299447 476234
rect 298572 476176 299386 476232
rect 299442 476176 299447 476232
rect 298572 476174 299447 476176
rect 298572 476172 298578 476174
rect 299381 476171 299447 476174
rect 300894 476172 300900 476236
rect 300964 476234 300970 476236
rect 302141 476234 302207 476237
rect 300964 476232 302207 476234
rect 300964 476176 302146 476232
rect 302202 476176 302207 476232
rect 300964 476174 302207 476176
rect 300964 476172 300970 476174
rect 302141 476171 302207 476174
rect 311014 476172 311020 476236
rect 311084 476234 311090 476236
rect 311801 476234 311867 476237
rect 311084 476232 311867 476234
rect 311084 476176 311806 476232
rect 311862 476176 311867 476232
rect 311084 476174 311867 476176
rect 311084 476172 311090 476174
rect 311801 476171 311867 476174
rect 315798 476172 315804 476236
rect 315868 476234 315874 476236
rect 315941 476234 316007 476237
rect 315868 476232 316007 476234
rect 315868 476176 315946 476232
rect 316002 476176 316007 476232
rect 315868 476174 316007 476176
rect 315868 476172 315874 476174
rect 315941 476171 316007 476174
rect 326654 476172 326660 476236
rect 326724 476234 326730 476236
rect 326981 476234 327047 476237
rect 326724 476232 327047 476234
rect 326724 476176 326986 476232
rect 327042 476176 327047 476232
rect 326724 476174 327047 476176
rect 326724 476172 326730 476174
rect 326981 476171 327047 476174
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3233 462634 3299 462637
rect -960 462632 3299 462634
rect -960 462576 3238 462632
rect 3294 462576 3299 462632
rect -960 462574 3299 462576
rect -960 462484 480 462574
rect 3233 462571 3299 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 237465 436250 237531 436253
rect 368974 436250 368980 436252
rect 237465 436248 368980 436250
rect 237465 436192 237470 436248
rect 237526 436192 368980 436248
rect 237465 436190 368980 436192
rect 237465 436187 237531 436190
rect 368974 436188 368980 436190
rect 369044 436188 369050 436252
rect 235717 436114 235783 436117
rect 367686 436114 367692 436116
rect 235717 436112 367692 436114
rect 235717 436056 235722 436112
rect 235778 436056 367692 436112
rect 235717 436054 367692 436056
rect 235717 436051 235783 436054
rect 367686 436052 367692 436054
rect 367756 436052 367762 436116
rect 214414 435236 214420 435300
rect 214484 435298 214490 435300
rect 294689 435298 294755 435301
rect 214484 435296 294755 435298
rect 214484 435240 294694 435296
rect 294750 435240 294755 435296
rect 214484 435238 294755 435240
rect 214484 435236 214490 435238
rect 294689 435235 294755 435238
rect 215886 435100 215892 435164
rect 215956 435162 215962 435164
rect 300117 435162 300183 435165
rect 215956 435160 300183 435162
rect 215956 435104 300122 435160
rect 300178 435104 300183 435160
rect 215956 435102 300183 435104
rect 215956 435100 215962 435102
rect 300117 435099 300183 435102
rect 211654 434964 211660 435028
rect 211724 435026 211730 435028
rect 296437 435026 296503 435029
rect 211724 435024 296503 435026
rect 211724 434968 296442 435024
rect 296498 434968 296503 435024
rect 211724 434966 296503 434968
rect 211724 434964 211730 434966
rect 296437 434963 296503 434966
rect 236269 434890 236335 434893
rect 360694 434890 360700 434892
rect 236269 434888 360700 434890
rect 236269 434832 236274 434888
rect 236330 434832 360700 434888
rect 236269 434830 360700 434832
rect 236269 434827 236335 434830
rect 360694 434828 360700 434830
rect 360764 434828 360770 434892
rect 234429 434754 234495 434757
rect 359406 434754 359412 434756
rect 234429 434752 359412 434754
rect 234429 434696 234434 434752
rect 234490 434696 359412 434752
rect 234429 434694 359412 434696
rect 234429 434691 234495 434694
rect 359406 434692 359412 434694
rect 359476 434692 359482 434756
rect 253197 433938 253263 433941
rect 298921 433938 298987 433941
rect 253197 433936 298987 433938
rect 253197 433880 253202 433936
rect 253258 433880 298926 433936
rect 298982 433880 298987 433936
rect 253197 433878 298987 433880
rect 253197 433875 253263 433878
rect 298921 433875 298987 433878
rect 233877 433802 233943 433805
rect 357893 433802 357959 433805
rect 233877 433800 357959 433802
rect 233877 433744 233882 433800
rect 233938 433744 357898 433800
rect 357954 433744 357959 433800
rect 233877 433742 357959 433744
rect 233877 433739 233943 433742
rect 357893 433739 357959 433742
rect 239305 433666 239371 433669
rect 579981 433666 580047 433669
rect 239305 433664 580047 433666
rect 239305 433608 239310 433664
rect 239366 433608 579986 433664
rect 580042 433608 580047 433664
rect 239305 433606 580047 433608
rect 239305 433603 239371 433606
rect 579981 433603 580047 433606
rect 238109 433530 238175 433533
rect 580441 433530 580507 433533
rect 238109 433528 580507 433530
rect 238109 433472 238114 433528
rect 238170 433472 580446 433528
rect 580502 433472 580507 433528
rect 238109 433470 580507 433472
rect 238109 433467 238175 433470
rect 580441 433467 580507 433470
rect 232681 433394 232747 433397
rect 580257 433394 580323 433397
rect 232681 433392 580323 433394
rect 232681 433336 232686 433392
rect 232742 433336 580262 433392
rect 580318 433336 580323 433392
rect 232681 433334 580323 433336
rect 232681 433331 232747 433334
rect 580257 433331 580323 433334
rect 240041 432306 240107 432309
rect 358486 432306 358492 432308
rect 240041 432304 358492 432306
rect 240041 432248 240046 432304
rect 240102 432248 358492 432304
rect 240041 432246 358492 432248
rect 240041 432243 240107 432246
rect 358486 432244 358492 432246
rect 358556 432244 358562 432308
rect 237281 432170 237347 432173
rect 358302 432170 358308 432172
rect 237281 432168 358308 432170
rect 237281 432112 237286 432168
rect 237342 432112 358308 432168
rect 237281 432110 358308 432112
rect 237281 432107 237347 432110
rect 358302 432108 358308 432110
rect 358372 432108 358378 432172
rect 235441 432034 235507 432037
rect 358118 432034 358124 432036
rect 235441 432032 358124 432034
rect 235441 431976 235446 432032
rect 235502 431976 358124 432032
rect 235441 431974 358124 431976
rect 235441 431971 235507 431974
rect 358118 431972 358124 431974
rect 358188 431972 358194 432036
rect 243353 431762 243419 431765
rect 245694 431762 245700 431764
rect 243353 431760 245700 431762
rect 243353 431704 243358 431760
rect 243414 431704 245700 431760
rect 243353 431702 245700 431704
rect 243353 431699 243419 431702
rect 245694 431700 245700 431702
rect 245764 431700 245770 431764
rect 299473 431762 299539 431765
rect 296670 431760 299539 431762
rect 296670 431704 299478 431760
rect 299534 431704 299539 431760
rect 296670 431702 299539 431704
rect 25497 430810 25563 430813
rect 296670 430810 296730 431702
rect 299473 431699 299539 431702
rect 579889 431626 579955 431629
rect 583520 431626 584960 431716
rect 579889 431624 584960 431626
rect 579889 431568 579894 431624
rect 579950 431568 584960 431624
rect 579889 431566 584960 431568
rect 579889 431563 579955 431566
rect 583520 431476 584960 431566
rect 25497 430808 296730 430810
rect 25497 430752 25502 430808
rect 25558 430752 296730 430808
rect 25497 430750 296730 430752
rect 25497 430747 25563 430750
rect 245694 430612 245700 430676
rect 245764 430674 245770 430676
rect 577589 430674 577655 430677
rect 245764 430672 577655 430674
rect 245764 430616 577594 430672
rect 577650 430616 577655 430672
rect 245764 430614 577655 430616
rect 245764 430612 245770 430614
rect 577589 430611 577655 430614
rect -960 423602 480 423692
rect 3325 423602 3391 423605
rect -960 423600 3391 423602
rect -960 423544 3330 423600
rect 3386 423544 3391 423600
rect -960 423542 3391 423544
rect -960 423452 480 423542
rect 3325 423539 3391 423542
rect 579981 418298 580047 418301
rect 583520 418298 584960 418388
rect 579981 418296 584960 418298
rect 579981 418240 579986 418296
rect 580042 418240 584960 418296
rect 579981 418238 584960 418240
rect 579981 418235 580047 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 579981 404970 580047 404973
rect 583520 404970 584960 405060
rect 579981 404968 584960 404970
rect 579981 404912 579986 404968
rect 580042 404912 584960 404968
rect 579981 404910 584960 404912
rect 579981 404907 580047 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580073 378450 580139 378453
rect 583520 378450 584960 378540
rect 580073 378448 584960 378450
rect 580073 378392 580078 378448
rect 580134 378392 584960 378448
rect 580073 378390 584960 378392
rect 580073 378387 580139 378390
rect 583520 378300 584960 378390
rect 159909 374098 159975 374101
rect 232078 374098 232084 374100
rect 159909 374096 232084 374098
rect 159909 374040 159914 374096
rect 159970 374040 232084 374096
rect 159909 374038 232084 374040
rect 159909 374035 159975 374038
rect 232078 374036 232084 374038
rect 232148 374036 232154 374100
rect 134149 372738 134215 372741
rect 232078 372738 232084 372740
rect 134149 372736 232084 372738
rect 134149 372680 134154 372736
rect 134210 372680 232084 372736
rect 134149 372678 232084 372680
rect 134149 372675 134215 372678
rect 232078 372676 232084 372678
rect 232148 372676 232154 372740
rect 118325 371650 118391 371653
rect 119061 371650 119127 371653
rect 118325 371648 119127 371650
rect 118325 371592 118330 371648
rect 118386 371592 119066 371648
rect 119122 371592 119127 371648
rect 118325 371590 119127 371592
rect 118325 371587 118391 371590
rect 119061 371587 119127 371590
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 231485 370290 231551 370293
rect 100710 370288 231551 370290
rect 100710 370232 231490 370288
rect 231546 370232 231551 370288
rect 100710 370230 231551 370232
rect 100710 370124 100770 370230
rect 231485 370227 231551 370230
rect 172329 369474 172395 369477
rect 169924 369472 172395 369474
rect 169924 369416 172334 369472
rect 172390 369416 172395 369472
rect 169924 369414 172395 369416
rect 172329 369411 172395 369414
rect 99833 367978 99899 367981
rect 99833 367976 100218 367978
rect 99833 367920 99838 367976
rect 99894 367920 100218 367976
rect 99833 367918 100218 367920
rect 99833 367915 99899 367918
rect 100158 367404 100218 367918
rect 171961 366754 172027 366757
rect 169924 366752 172027 366754
rect 169924 366696 171966 366752
rect 172022 366696 172027 366752
rect 169924 366694 172027 366696
rect 171961 366691 172027 366694
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect 97809 364714 97875 364717
rect 97809 364712 100188 364714
rect 97809 364656 97814 364712
rect 97870 364656 100188 364712
rect 97809 364654 100188 364656
rect 97809 364651 97875 364654
rect 172329 364034 172395 364037
rect 169924 364032 172395 364034
rect 169924 363976 172334 364032
rect 172390 363976 172395 364032
rect 169924 363974 172395 363976
rect 172329 363971 172395 363974
rect 97717 361994 97783 361997
rect 97717 361992 100188 361994
rect 97717 361936 97722 361992
rect 97778 361936 100188 361992
rect 97717 361934 100188 361936
rect 97717 361931 97783 361934
rect 172053 361314 172119 361317
rect 169924 361312 172119 361314
rect 169924 361256 172058 361312
rect 172114 361256 172119 361312
rect 169924 361254 172119 361256
rect 172053 361251 172119 361254
rect 99281 359274 99347 359277
rect 99281 359272 100188 359274
rect 99281 359216 99286 359272
rect 99342 359216 100188 359272
rect 99281 359214 100188 359216
rect 99281 359211 99347 359214
rect 172421 358594 172487 358597
rect 169924 358592 172487 358594
rect -960 358458 480 358548
rect 169924 358536 172426 358592
rect 172482 358536 172487 358592
rect 169924 358534 172487 358536
rect 172421 358531 172487 358534
rect 3693 358458 3759 358461
rect -960 358456 3759 358458
rect -960 358400 3698 358456
rect 3754 358400 3759 358456
rect -960 358398 3759 358400
rect -960 358308 480 358398
rect 3693 358395 3759 358398
rect 97809 356554 97875 356557
rect 97809 356552 100188 356554
rect 97809 356496 97814 356552
rect 97870 356496 100188 356552
rect 97809 356494 100188 356496
rect 97809 356491 97875 356494
rect 172421 355874 172487 355877
rect 169924 355872 172487 355874
rect 169924 355816 172426 355872
rect 172482 355816 172487 355872
rect 169924 355814 172487 355816
rect 172421 355811 172487 355814
rect 99189 353834 99255 353837
rect 99189 353832 100188 353834
rect 99189 353776 99194 353832
rect 99250 353776 100188 353832
rect 99189 353774 100188 353776
rect 99189 353771 99255 353774
rect 172421 353154 172487 353157
rect 169924 353152 172487 353154
rect 169924 353096 172426 353152
rect 172482 353096 172487 353152
rect 169924 353094 172487 353096
rect 172421 353091 172487 353094
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect 97901 351114 97967 351117
rect 97901 351112 100188 351114
rect 97901 351056 97906 351112
rect 97962 351056 100188 351112
rect 97901 351054 100188 351056
rect 97901 351051 97967 351054
rect 171777 350434 171843 350437
rect 169924 350432 171843 350434
rect 169924 350376 171782 350432
rect 171838 350376 171843 350432
rect 169924 350374 171843 350376
rect 171777 350371 171843 350374
rect 97901 348394 97967 348397
rect 97901 348392 100188 348394
rect 97901 348336 97906 348392
rect 97962 348336 100188 348392
rect 97901 348334 100188 348336
rect 97901 348331 97967 348334
rect 172421 347714 172487 347717
rect 169924 347712 172487 347714
rect 169924 347656 172426 347712
rect 172482 347656 172487 347712
rect 169924 347654 172487 347656
rect 172421 347651 172487 347654
rect 97717 345674 97783 345677
rect 97717 345672 100188 345674
rect 97717 345616 97722 345672
rect 97778 345616 100188 345672
rect 97717 345614 100188 345616
rect 97717 345611 97783 345614
rect -960 345402 480 345492
rect 3601 345402 3667 345405
rect -960 345400 3667 345402
rect -960 345344 3606 345400
rect 3662 345344 3667 345400
rect -960 345342 3667 345344
rect -960 345252 480 345342
rect 3601 345339 3667 345342
rect 172145 344994 172211 344997
rect 169924 344992 172211 344994
rect 169924 344936 172150 344992
rect 172206 344936 172211 344992
rect 169924 344934 172211 344936
rect 172145 344931 172211 344934
rect 99097 342954 99163 342957
rect 99097 342952 100188 342954
rect 99097 342896 99102 342952
rect 99158 342896 100188 342952
rect 99097 342894 100188 342896
rect 99097 342891 99163 342894
rect 172421 342274 172487 342277
rect 169924 342272 172487 342274
rect 169924 342216 172426 342272
rect 172482 342216 172487 342272
rect 169924 342214 172487 342216
rect 172421 342211 172487 342214
rect 97625 340234 97691 340237
rect 97625 340232 100188 340234
rect 97625 340176 97630 340232
rect 97686 340176 100188 340232
rect 97625 340174 100188 340176
rect 97625 340171 97691 340174
rect 172421 339554 172487 339557
rect 169924 339552 172487 339554
rect 169924 339496 172426 339552
rect 172482 339496 172487 339552
rect 169924 339494 172487 339496
rect 172421 339491 172487 339494
rect 583520 338452 584960 338692
rect 99005 337514 99071 337517
rect 99005 337512 100188 337514
rect 99005 337456 99010 337512
rect 99066 337456 100188 337512
rect 99005 337454 100188 337456
rect 99005 337451 99071 337454
rect 172421 336834 172487 336837
rect 169924 336832 172487 336834
rect 169924 336776 172426 336832
rect 172482 336776 172487 336832
rect 169924 336774 172487 336776
rect 172421 336771 172487 336774
rect 99373 334794 99439 334797
rect 99373 334792 100188 334794
rect 99373 334736 99378 334792
rect 99434 334736 100188 334792
rect 99373 334734 100188 334736
rect 99373 334731 99439 334734
rect 172237 334114 172303 334117
rect 169924 334112 172303 334114
rect 169924 334056 172242 334112
rect 172298 334056 172303 334112
rect 169924 334054 172303 334056
rect 172237 334051 172303 334054
rect -960 332196 480 332436
rect 97533 332074 97599 332077
rect 97533 332072 100188 332074
rect 97533 332016 97538 332072
rect 97594 332016 100188 332072
rect 97533 332014 100188 332016
rect 97533 332011 97599 332014
rect 172421 331394 172487 331397
rect 169924 331392 172487 331394
rect 169924 331336 172426 331392
rect 172482 331336 172487 331392
rect 169924 331334 172487 331336
rect 172421 331331 172487 331334
rect 98913 329354 98979 329357
rect 98913 329352 100188 329354
rect 98913 329296 98918 329352
rect 98974 329296 100188 329352
rect 98913 329294 100188 329296
rect 98913 329291 98979 329294
rect 172421 328674 172487 328677
rect 169924 328672 172487 328674
rect 169924 328616 172426 328672
rect 172482 328616 172487 328672
rect 169924 328614 172487 328616
rect 172421 328611 172487 328614
rect 97441 326634 97507 326637
rect 97441 326632 100188 326634
rect 97441 326576 97446 326632
rect 97502 326576 100188 326632
rect 97441 326574 100188 326576
rect 97441 326571 97507 326574
rect 172329 325954 172395 325957
rect 169924 325952 172395 325954
rect 169924 325896 172334 325952
rect 172390 325896 172395 325952
rect 169924 325894 172395 325896
rect 172329 325891 172395 325894
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 98821 323914 98887 323917
rect 98821 323912 100188 323914
rect 98821 323856 98826 323912
rect 98882 323856 100188 323912
rect 98821 323854 100188 323856
rect 98821 323851 98887 323854
rect 171317 323234 171383 323237
rect 169924 323232 171383 323234
rect 169924 323176 171322 323232
rect 171378 323176 171383 323232
rect 169924 323174 171383 323176
rect 171317 323171 171383 323174
rect 98545 321194 98611 321197
rect 98545 321192 100188 321194
rect 98545 321136 98550 321192
rect 98606 321136 100188 321192
rect 98545 321134 100188 321136
rect 98545 321131 98611 321134
rect 171501 320514 171567 320517
rect 169924 320512 171567 320514
rect 169924 320456 171506 320512
rect 171562 320456 171567 320512
rect 169924 320454 171567 320456
rect 171501 320451 171567 320454
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 98729 318474 98795 318477
rect 98729 318472 100188 318474
rect 98729 318416 98734 318472
rect 98790 318416 100188 318472
rect 98729 318414 100188 318416
rect 98729 318411 98795 318414
rect 171501 317794 171567 317797
rect 169924 317792 171567 317794
rect 169924 317736 171506 317792
rect 171562 317736 171567 317792
rect 169924 317734 171567 317736
rect 171501 317731 171567 317734
rect 97349 315754 97415 315757
rect 97349 315752 100188 315754
rect 97349 315696 97354 315752
rect 97410 315696 100188 315752
rect 97349 315694 100188 315696
rect 97349 315691 97415 315694
rect 172421 315074 172487 315077
rect 169924 315072 172487 315074
rect 169924 315016 172426 315072
rect 172482 315016 172487 315072
rect 169924 315014 172487 315016
rect 172421 315011 172487 315014
rect 99465 313034 99531 313037
rect 99465 313032 100188 313034
rect 99465 312976 99470 313032
rect 99526 312976 100188 313032
rect 99465 312974 100188 312976
rect 99465 312971 99531 312974
rect 172421 312354 172487 312357
rect 169924 312352 172487 312354
rect 169924 312296 172426 312352
rect 172482 312296 172487 312352
rect 169924 312294 172487 312296
rect 172421 312291 172487 312294
rect 580901 312082 580967 312085
rect 583520 312082 584960 312172
rect 580901 312080 584960 312082
rect 580901 312024 580906 312080
rect 580962 312024 584960 312080
rect 580901 312022 584960 312024
rect 580901 312019 580967 312022
rect 583520 311932 584960 312022
rect 226977 310586 227043 310589
rect 232773 310586 232839 310589
rect 226977 310584 232839 310586
rect 226977 310528 226982 310584
rect 227038 310528 232778 310584
rect 232834 310528 232839 310584
rect 226977 310526 232839 310528
rect 226977 310523 227043 310526
rect 232773 310523 232839 310526
rect 231853 310450 231919 310453
rect 232221 310450 232287 310453
rect 231853 310448 232287 310450
rect 231853 310392 231858 310448
rect 231914 310392 232226 310448
rect 232282 310392 232287 310448
rect 231853 310390 232287 310392
rect 231853 310387 231919 310390
rect 232221 310387 232287 310390
rect 97257 310314 97323 310317
rect 231209 310314 231275 310317
rect 234981 310314 235047 310317
rect 97257 310312 100188 310314
rect 97257 310256 97262 310312
rect 97318 310256 100188 310312
rect 97257 310254 100188 310256
rect 231209 310312 235047 310314
rect 231209 310256 231214 310312
rect 231270 310256 234986 310312
rect 235042 310256 235047 310312
rect 231209 310254 235047 310256
rect 97257 310251 97323 310254
rect 231209 310251 231275 310254
rect 234981 310251 235047 310254
rect 232630 309844 232636 309908
rect 232700 309906 232706 309908
rect 246205 309906 246271 309909
rect 232700 309904 246271 309906
rect 232700 309848 246210 309904
rect 246266 309848 246271 309904
rect 232700 309846 246271 309848
rect 232700 309844 232706 309846
rect 246205 309843 246271 309846
rect 170765 309770 170831 309773
rect 230013 309770 230079 309773
rect 246849 309770 246915 309773
rect 170765 309768 180810 309770
rect 170765 309712 170770 309768
rect 170826 309712 180810 309768
rect 170765 309710 180810 309712
rect 170765 309707 170831 309710
rect 172421 309634 172487 309637
rect 169924 309632 172487 309634
rect 169924 309576 172426 309632
rect 172482 309576 172487 309632
rect 169924 309574 172487 309576
rect 180750 309634 180810 309710
rect 230013 309768 246915 309770
rect 230013 309712 230018 309768
rect 230074 309712 246854 309768
rect 246910 309712 246915 309768
rect 230013 309710 246915 309712
rect 230013 309707 230079 309710
rect 246849 309707 246915 309710
rect 240501 309634 240567 309637
rect 180750 309632 240567 309634
rect 180750 309576 240506 309632
rect 240562 309576 240567 309632
rect 180750 309574 240567 309576
rect 172421 309571 172487 309574
rect 240501 309571 240567 309574
rect 173249 309498 173315 309501
rect 245285 309498 245351 309501
rect 173249 309496 245351 309498
rect 173249 309440 173254 309496
rect 173310 309440 245290 309496
rect 245346 309440 245351 309496
rect 173249 309438 245351 309440
rect 173249 309435 173315 309438
rect 245285 309435 245351 309438
rect 170949 309362 171015 309365
rect 245469 309362 245535 309365
rect 170949 309360 245535 309362
rect 170949 309304 170954 309360
rect 171010 309304 245474 309360
rect 245530 309304 245535 309360
rect 170949 309302 245535 309304
rect 170949 309299 171015 309302
rect 245469 309299 245535 309302
rect 174629 309226 174695 309229
rect 250253 309226 250319 309229
rect 174629 309224 250319 309226
rect 174629 309168 174634 309224
rect 174690 309168 250258 309224
rect 250314 309168 250319 309224
rect 174629 309166 250319 309168
rect 174629 309163 174695 309166
rect 250253 309163 250319 309166
rect 229921 309090 229987 309093
rect 234337 309090 234403 309093
rect 229921 309088 234403 309090
rect 229921 309032 229926 309088
rect 229982 309032 234342 309088
rect 234398 309032 234403 309088
rect 229921 309030 234403 309032
rect 229921 309027 229987 309030
rect 234337 309027 234403 309030
rect 234470 309028 234476 309092
rect 234540 309090 234546 309092
rect 235349 309090 235415 309093
rect 234540 309088 235415 309090
rect 234540 309032 235354 309088
rect 235410 309032 235415 309088
rect 234540 309030 235415 309032
rect 234540 309028 234546 309030
rect 235349 309027 235415 309030
rect 338665 309090 338731 309093
rect 362217 309090 362283 309093
rect 338665 309088 362283 309090
rect 338665 309032 338670 309088
rect 338726 309032 362222 309088
rect 362278 309032 362283 309088
rect 338665 309030 362283 309032
rect 338665 309027 338731 309030
rect 362217 309027 362283 309030
rect 173433 308954 173499 308957
rect 247033 308954 247099 308957
rect 173433 308952 247099 308954
rect 173433 308896 173438 308952
rect 173494 308896 247038 308952
rect 247094 308896 247099 308952
rect 173433 308894 247099 308896
rect 173433 308891 173499 308894
rect 247033 308891 247099 308894
rect 339217 308954 339283 308957
rect 362309 308954 362375 308957
rect 339217 308952 362375 308954
rect 339217 308896 339222 308952
rect 339278 308896 362314 308952
rect 362370 308896 362375 308952
rect 339217 308894 362375 308896
rect 339217 308891 339283 308894
rect 362309 308891 362375 308894
rect 173617 308818 173683 308821
rect 243353 308818 243419 308821
rect 173617 308816 243419 308818
rect 173617 308760 173622 308816
rect 173678 308760 243358 308816
rect 243414 308760 243419 308816
rect 173617 308758 243419 308760
rect 173617 308755 173683 308758
rect 243353 308755 243419 308758
rect 303981 308818 304047 308821
rect 360193 308818 360259 308821
rect 303981 308816 360259 308818
rect 303981 308760 303986 308816
rect 304042 308760 360198 308816
rect 360254 308760 360259 308816
rect 303981 308758 360259 308760
rect 303981 308755 304047 308758
rect 360193 308755 360259 308758
rect 231485 308682 231551 308685
rect 234470 308682 234476 308684
rect 231485 308680 234476 308682
rect 231485 308624 231490 308680
rect 231546 308624 234476 308680
rect 231485 308622 234476 308624
rect 231485 308619 231551 308622
rect 234470 308620 234476 308622
rect 234540 308620 234546 308684
rect 239397 308682 239463 308685
rect 251173 308682 251239 308685
rect 239397 308680 251239 308682
rect 239397 308624 239402 308680
rect 239458 308624 251178 308680
rect 251234 308624 251239 308680
rect 239397 308622 251239 308624
rect 239397 308619 239463 308622
rect 251173 308619 251239 308622
rect 298461 308682 298527 308685
rect 355409 308682 355475 308685
rect 298461 308680 355475 308682
rect 298461 308624 298466 308680
rect 298522 308624 355414 308680
rect 355470 308624 355475 308680
rect 298461 308622 355475 308624
rect 298461 308619 298527 308622
rect 355409 308619 355475 308622
rect 174537 308546 174603 308549
rect 250805 308546 250871 308549
rect 174537 308544 250871 308546
rect 174537 308488 174542 308544
rect 174598 308488 250810 308544
rect 250866 308488 250871 308544
rect 174537 308486 250871 308488
rect 174537 308483 174603 308486
rect 250805 308483 250871 308486
rect 299657 308546 299723 308549
rect 357525 308546 357591 308549
rect 299657 308544 357591 308546
rect 299657 308488 299662 308544
rect 299718 308488 357530 308544
rect 357586 308488 357591 308544
rect 299657 308486 357591 308488
rect 299657 308483 299723 308486
rect 357525 308483 357591 308486
rect 231301 308410 231367 308413
rect 239397 308410 239463 308413
rect 231301 308408 239463 308410
rect 231301 308352 231306 308408
rect 231362 308352 239402 308408
rect 239458 308352 239463 308408
rect 231301 308350 239463 308352
rect 231301 308347 231367 308350
rect 239397 308347 239463 308350
rect 298829 308410 298895 308413
rect 362493 308410 362559 308413
rect 298829 308408 362559 308410
rect 298829 308352 298834 308408
rect 298890 308352 362498 308408
rect 362554 308352 362559 308408
rect 298829 308350 362559 308352
rect 298829 308347 298895 308350
rect 362493 308347 362559 308350
rect 232446 308212 232452 308276
rect 232516 308274 232522 308276
rect 242433 308274 242499 308277
rect 232516 308272 242499 308274
rect 232516 308216 242438 308272
rect 242494 308216 242499 308272
rect 232516 308214 242499 308216
rect 232516 308212 232522 308214
rect 242433 308211 242499 308214
rect 338481 308274 338547 308277
rect 359549 308274 359615 308277
rect 338481 308272 359615 308274
rect 338481 308216 338486 308272
rect 338542 308216 359554 308272
rect 359610 308216 359615 308272
rect 338481 308214 359615 308216
rect 338481 308211 338547 308214
rect 359549 308211 359615 308214
rect 98637 307594 98703 307597
rect 98637 307592 100188 307594
rect 98637 307536 98642 307592
rect 98698 307536 100188 307592
rect 98637 307534 100188 307536
rect 98637 307531 98703 307534
rect 172421 306914 172487 306917
rect 169924 306912 172487 306914
rect 169924 306856 172426 306912
rect 172482 306856 172487 306912
rect 169924 306854 172487 306856
rect 172421 306851 172487 306854
rect 333145 306506 333211 306509
rect 333102 306504 333211 306506
rect 333102 306448 333150 306504
rect 333206 306448 333211 306504
rect 333102 306443 333211 306448
rect 306649 306370 306715 306373
rect 306606 306368 306715 306370
rect -960 306234 480 306324
rect 306606 306312 306654 306368
rect 306710 306312 306715 306368
rect 306606 306307 306715 306312
rect 3325 306234 3391 306237
rect -960 306232 3391 306234
rect -960 306176 3330 306232
rect 3386 306176 3391 306232
rect -960 306174 3391 306176
rect -960 306084 480 306174
rect 3325 306171 3391 306174
rect 219014 306172 219020 306236
rect 219084 306234 219090 306236
rect 284845 306234 284911 306237
rect 219084 306232 284911 306234
rect 219084 306176 284850 306232
rect 284906 306176 284911 306232
rect 219084 306174 284911 306176
rect 219084 306172 219090 306174
rect 284845 306171 284911 306174
rect 218830 306036 218836 306100
rect 218900 306098 218906 306100
rect 284293 306098 284359 306101
rect 218900 306096 284359 306098
rect 218900 306040 284298 306096
rect 284354 306040 284359 306096
rect 218900 306038 284359 306040
rect 218900 306036 218906 306038
rect 284293 306035 284359 306038
rect 306465 306098 306531 306101
rect 306606 306098 306666 306307
rect 333102 306237 333162 306443
rect 336917 306370 336983 306373
rect 340137 306370 340203 306373
rect 362401 306370 362467 306373
rect 336917 306368 338866 306370
rect 336917 306312 336922 306368
rect 336978 306312 338866 306368
rect 336917 306310 338866 306312
rect 336917 306307 336983 306310
rect 333053 306232 333162 306237
rect 333053 306176 333058 306232
rect 333114 306176 333162 306232
rect 333053 306174 333162 306176
rect 333053 306171 333119 306174
rect 306465 306096 306666 306098
rect 306465 306040 306470 306096
rect 306526 306040 306666 306096
rect 306465 306038 306666 306040
rect 306465 306035 306531 306038
rect 217542 305900 217548 305964
rect 217612 305962 217618 305964
rect 286961 305962 287027 305965
rect 217612 305960 287027 305962
rect 217612 305904 286966 305960
rect 287022 305904 287027 305960
rect 217612 305902 287027 305904
rect 217612 305900 217618 305902
rect 286961 305899 287027 305902
rect 217358 305764 217364 305828
rect 217428 305826 217434 305828
rect 285857 305826 285923 305829
rect 217428 305824 285923 305826
rect 217428 305768 285862 305824
rect 285918 305768 285923 305824
rect 217428 305766 285923 305768
rect 338806 305826 338866 306310
rect 340137 306368 362467 306370
rect 340137 306312 340142 306368
rect 340198 306312 362406 306368
rect 362462 306312 362467 306368
rect 340137 306310 362467 306312
rect 340137 306307 340203 306310
rect 362401 306307 362467 306310
rect 343725 306234 343791 306237
rect 368657 306234 368723 306237
rect 343725 306232 368723 306234
rect 343725 306176 343730 306232
rect 343786 306176 368662 306232
rect 368718 306176 368723 306232
rect 343725 306174 368723 306176
rect 343725 306171 343791 306174
rect 368657 306171 368723 306174
rect 340781 306098 340847 306101
rect 365989 306098 366055 306101
rect 340781 306096 366055 306098
rect 340781 306040 340786 306096
rect 340842 306040 365994 306096
rect 366050 306040 366055 306096
rect 340781 306038 366055 306040
rect 340781 306035 340847 306038
rect 365989 306035 366055 306038
rect 341517 305962 341583 305965
rect 368749 305962 368815 305965
rect 341517 305960 368815 305962
rect 341517 305904 341522 305960
rect 341578 305904 368754 305960
rect 368810 305904 368815 305960
rect 341517 305902 368815 305904
rect 341517 305899 341583 305902
rect 368749 305899 368815 305902
rect 378777 305826 378843 305829
rect 338806 305824 378843 305826
rect 338806 305768 378782 305824
rect 378838 305768 378843 305824
rect 338806 305766 378843 305768
rect 217428 305764 217434 305766
rect 285857 305763 285923 305766
rect 378777 305763 378843 305766
rect 170397 305690 170463 305693
rect 253473 305690 253539 305693
rect 170397 305688 253539 305690
rect 170397 305632 170402 305688
rect 170458 305632 253478 305688
rect 253534 305632 253539 305688
rect 170397 305630 253539 305632
rect 170397 305627 170463 305630
rect 253473 305627 253539 305630
rect 295057 305690 295123 305693
rect 357985 305690 358051 305693
rect 295057 305688 358051 305690
rect 295057 305632 295062 305688
rect 295118 305632 357990 305688
rect 358046 305632 358051 305688
rect 295057 305630 358051 305632
rect 295057 305627 295123 305630
rect 357985 305627 358051 305630
rect 97901 304874 97967 304877
rect 97901 304872 100188 304874
rect 97901 304816 97906 304872
rect 97962 304816 100188 304872
rect 97901 304814 100188 304816
rect 97901 304811 97967 304814
rect 172329 304194 172395 304197
rect 169924 304192 172395 304194
rect 169924 304136 172334 304192
rect 172390 304136 172395 304192
rect 169924 304134 172395 304136
rect 172329 304131 172395 304134
rect 344921 303514 344987 303517
rect 363689 303514 363755 303517
rect 344921 303512 363755 303514
rect 344921 303456 344926 303512
rect 344982 303456 363694 303512
rect 363750 303456 363755 303512
rect 344921 303454 363755 303456
rect 344921 303451 344987 303454
rect 363689 303451 363755 303454
rect 216438 303316 216444 303380
rect 216508 303378 216514 303380
rect 285029 303378 285095 303381
rect 216508 303376 285095 303378
rect 216508 303320 285034 303376
rect 285090 303320 285095 303376
rect 216508 303318 285095 303320
rect 216508 303316 216514 303318
rect 285029 303315 285095 303318
rect 345197 303378 345263 303381
rect 367921 303378 367987 303381
rect 345197 303376 367987 303378
rect 345197 303320 345202 303376
rect 345258 303320 367926 303376
rect 367982 303320 367987 303376
rect 345197 303318 367987 303320
rect 345197 303315 345263 303318
rect 367921 303315 367987 303318
rect 214782 303180 214788 303244
rect 214852 303242 214858 303244
rect 284109 303242 284175 303245
rect 214852 303240 284175 303242
rect 214852 303184 284114 303240
rect 284170 303184 284175 303240
rect 214852 303182 284175 303184
rect 214852 303180 214858 303182
rect 284109 303179 284175 303182
rect 339493 303242 339559 303245
rect 366449 303242 366515 303245
rect 339493 303240 366515 303242
rect 339493 303184 339498 303240
rect 339554 303184 366454 303240
rect 366510 303184 366515 303240
rect 339493 303182 366515 303184
rect 339493 303179 339559 303182
rect 366449 303179 366515 303182
rect 216070 303044 216076 303108
rect 216140 303106 216146 303108
rect 284661 303106 284727 303109
rect 216140 303104 284727 303106
rect 216140 303048 284666 303104
rect 284722 303048 284727 303104
rect 216140 303046 284727 303048
rect 216140 303044 216146 303046
rect 284661 303043 284727 303046
rect 338849 303106 338915 303109
rect 365161 303106 365227 303109
rect 338849 303104 365227 303106
rect 338849 303048 338854 303104
rect 338910 303048 365166 303104
rect 365222 303048 365227 303104
rect 338849 303046 365227 303048
rect 338849 303043 338915 303046
rect 365161 303043 365227 303046
rect 215150 302908 215156 302972
rect 215220 302970 215226 302972
rect 284477 302970 284543 302973
rect 215220 302968 284543 302970
rect 215220 302912 284482 302968
rect 284538 302912 284543 302968
rect 215220 302910 284543 302912
rect 215220 302908 215226 302910
rect 284477 302907 284543 302910
rect 305637 302970 305703 302973
rect 362902 302970 362908 302972
rect 305637 302968 362908 302970
rect 305637 302912 305642 302968
rect 305698 302912 362908 302968
rect 305637 302910 362908 302912
rect 305637 302907 305703 302910
rect 362902 302908 362908 302910
rect 362972 302908 362978 302972
rect 216990 302772 216996 302836
rect 217060 302834 217066 302836
rect 288709 302834 288775 302837
rect 217060 302832 288775 302834
rect 217060 302776 288714 302832
rect 288770 302776 288775 302832
rect 217060 302774 288775 302776
rect 217060 302772 217066 302774
rect 288709 302771 288775 302774
rect 294321 302834 294387 302837
rect 363781 302834 363847 302837
rect 294321 302832 363847 302834
rect 294321 302776 294326 302832
rect 294382 302776 363786 302832
rect 363842 302776 363847 302832
rect 294321 302774 363847 302776
rect 294321 302771 294387 302774
rect 363781 302771 363847 302774
rect 99833 302154 99899 302157
rect 99833 302152 100188 302154
rect 99833 302096 99838 302152
rect 99894 302096 100188 302152
rect 99833 302094 100188 302096
rect 99833 302091 99899 302094
rect 169753 301746 169819 301749
rect 169753 301744 171150 301746
rect 169753 301688 169758 301744
rect 169814 301688 171150 301744
rect 169753 301686 171150 301688
rect 169753 301683 169819 301686
rect 171090 301610 171150 301686
rect 214966 301684 214972 301748
rect 215036 301746 215042 301748
rect 283373 301746 283439 301749
rect 215036 301744 283439 301746
rect 215036 301688 283378 301744
rect 283434 301688 283439 301744
rect 215036 301686 283439 301688
rect 215036 301684 215042 301686
rect 283373 301683 283439 301686
rect 249977 301610 250043 301613
rect 171090 301608 250043 301610
rect 171090 301552 249982 301608
rect 250038 301552 250043 301608
rect 171090 301550 250043 301552
rect 249977 301547 250043 301550
rect 172421 301474 172487 301477
rect 169924 301472 172487 301474
rect 169924 301416 172426 301472
rect 172482 301416 172487 301472
rect 169924 301414 172487 301416
rect 172421 301411 172487 301414
rect 217174 301412 217180 301476
rect 217244 301474 217250 301476
rect 288617 301474 288683 301477
rect 217244 301472 288683 301474
rect 217244 301416 288622 301472
rect 288678 301416 288683 301472
rect 217244 301414 288683 301416
rect 217244 301412 217250 301414
rect 288617 301411 288683 301414
rect 169150 301140 169156 301204
rect 169220 301202 169226 301204
rect 239029 301202 239095 301205
rect 169220 301200 239095 301202
rect 169220 301144 239034 301200
rect 239090 301144 239095 301200
rect 169220 301142 239095 301144
rect 169220 301140 169226 301142
rect 239029 301139 239095 301142
rect 99281 300794 99347 300797
rect 244641 300794 244707 300797
rect 99281 300792 244707 300794
rect 99281 300736 99286 300792
rect 99342 300736 244646 300792
rect 244702 300736 244707 300792
rect 99281 300734 244707 300736
rect 99281 300731 99347 300734
rect 244641 300731 244707 300734
rect 166625 300658 166691 300661
rect 169845 300658 169911 300661
rect 166625 300656 169911 300658
rect 166625 300600 166630 300656
rect 166686 300600 169850 300656
rect 169906 300600 169911 300656
rect 166625 300598 169911 300600
rect 166625 300595 166691 300598
rect 169845 300595 169911 300598
rect 305545 300658 305611 300661
rect 358854 300658 358860 300660
rect 305545 300656 358860 300658
rect 305545 300600 305550 300656
rect 305606 300600 358860 300656
rect 305545 300598 358860 300600
rect 305545 300595 305611 300598
rect 358854 300596 358860 300598
rect 358924 300596 358930 300660
rect 211889 300522 211955 300525
rect 286133 300522 286199 300525
rect 211889 300520 286199 300522
rect 211889 300464 211894 300520
rect 211950 300464 286138 300520
rect 286194 300464 286199 300520
rect 211889 300462 286199 300464
rect 211889 300459 211955 300462
rect 286133 300459 286199 300462
rect 294229 300522 294295 300525
rect 358261 300522 358327 300525
rect 294229 300520 358327 300522
rect 294229 300464 294234 300520
rect 294290 300464 358266 300520
rect 358322 300464 358327 300520
rect 294229 300462 358327 300464
rect 294229 300459 294295 300462
rect 358261 300459 358327 300462
rect 168373 300386 168439 300389
rect 276473 300386 276539 300389
rect 168373 300384 276539 300386
rect 168373 300328 168378 300384
rect 168434 300328 276478 300384
rect 276534 300328 276539 300384
rect 168373 300326 276539 300328
rect 168373 300323 168439 300326
rect 276473 300323 276539 300326
rect 294689 300386 294755 300389
rect 366541 300386 366607 300389
rect 294689 300384 366607 300386
rect 294689 300328 294694 300384
rect 294750 300328 366546 300384
rect 366602 300328 366607 300384
rect 294689 300326 366607 300328
rect 294689 300323 294755 300326
rect 366541 300323 366607 300326
rect 160093 300250 160159 300253
rect 270033 300250 270099 300253
rect 160093 300248 270099 300250
rect 160093 300192 160098 300248
rect 160154 300192 270038 300248
rect 270094 300192 270099 300248
rect 160093 300190 270099 300192
rect 160093 300187 160159 300190
rect 270033 300187 270099 300190
rect 294781 300250 294847 300253
rect 370405 300250 370471 300253
rect 294781 300248 370471 300250
rect 294781 300192 294786 300248
rect 294842 300192 370410 300248
rect 370466 300192 370471 300248
rect 294781 300190 370471 300192
rect 294781 300187 294847 300190
rect 370405 300187 370471 300190
rect 32397 300114 32463 300117
rect 255865 300114 255931 300117
rect 32397 300112 255931 300114
rect 32397 300056 32402 300112
rect 32458 300056 255870 300112
rect 255926 300056 255931 300112
rect 32397 300054 255931 300056
rect 32397 300051 32463 300054
rect 255865 300051 255931 300054
rect 322105 300114 322171 300117
rect 467097 300114 467163 300117
rect 322105 300112 467163 300114
rect 322105 300056 322110 300112
rect 322166 300056 467102 300112
rect 467158 300056 467163 300112
rect 322105 300054 467163 300056
rect 322105 300051 322171 300054
rect 467097 300051 467163 300054
rect 97165 299434 97231 299437
rect 236453 299434 236519 299437
rect 97165 299432 236519 299434
rect 97165 299376 97170 299432
rect 97226 299376 236458 299432
rect 236514 299376 236519 299432
rect 97165 299374 236519 299376
rect 97165 299371 97231 299374
rect 236453 299371 236519 299374
rect 97533 299298 97599 299301
rect 233325 299298 233391 299301
rect 97533 299296 233391 299298
rect 97533 299240 97538 299296
rect 97594 299240 233330 299296
rect 233386 299240 233391 299296
rect 97533 299238 233391 299240
rect 97533 299235 97599 299238
rect 233325 299235 233391 299238
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 150893 297938 150959 297941
rect 169150 297938 169156 297940
rect 150893 297936 169156 297938
rect 150893 297880 150898 297936
rect 150954 297880 169156 297936
rect 150893 297878 169156 297880
rect 150893 297875 150959 297878
rect 169150 297876 169156 297878
rect 169220 297876 169226 297940
rect 214557 297938 214623 297941
rect 287605 297938 287671 297941
rect 214557 297936 287671 297938
rect 214557 297880 214562 297936
rect 214618 297880 287610 297936
rect 287666 297880 287671 297936
rect 214557 297878 287671 297880
rect 214557 297875 214623 297878
rect 287605 297875 287671 297878
rect 212349 297802 212415 297805
rect 287513 297802 287579 297805
rect 212349 297800 287579 297802
rect 212349 297744 212354 297800
rect 212410 297744 287518 297800
rect 287574 297744 287579 297800
rect 212349 297742 287579 297744
rect 212349 297739 212415 297742
rect 287513 297739 287579 297742
rect 211797 297666 211863 297669
rect 287421 297666 287487 297669
rect 211797 297664 287487 297666
rect 211797 297608 211802 297664
rect 211858 297608 287426 297664
rect 287482 297608 287487 297664
rect 211797 297606 287487 297608
rect 211797 297603 211863 297606
rect 287421 297603 287487 297606
rect 212165 297530 212231 297533
rect 289261 297530 289327 297533
rect 212165 297528 289327 297530
rect 212165 297472 212170 297528
rect 212226 297472 289266 297528
rect 289322 297472 289327 297528
rect 212165 297470 289327 297472
rect 212165 297467 212231 297470
rect 289261 297467 289327 297470
rect 211061 297394 211127 297397
rect 288893 297394 288959 297397
rect 211061 297392 288959 297394
rect 211061 297336 211066 297392
rect 211122 297336 288898 297392
rect 288954 297336 288959 297392
rect 211061 297334 288959 297336
rect 211061 297331 211127 297334
rect 288893 297331 288959 297334
rect 305453 296034 305519 296037
rect 360142 296034 360148 296036
rect 305453 296032 360148 296034
rect 305453 295976 305458 296032
rect 305514 295976 360148 296032
rect 305453 295974 360148 295976
rect 305453 295971 305519 295974
rect 360142 295972 360148 295974
rect 360212 295972 360218 296036
rect 305361 294538 305427 294541
rect 360878 294538 360884 294540
rect 305361 294536 360884 294538
rect 305361 294480 305366 294536
rect 305422 294480 360884 294536
rect 305361 294478 360884 294480
rect 305361 294475 305427 294478
rect 360878 294476 360884 294478
rect 360948 294476 360954 294540
rect -960 293178 480 293268
rect 3509 293178 3575 293181
rect -960 293176 3575 293178
rect -960 293120 3514 293176
rect 3570 293120 3575 293176
rect -960 293118 3575 293120
rect -960 293028 480 293118
rect 3509 293115 3575 293118
rect 219198 293116 219204 293180
rect 219268 293178 219274 293180
rect 283189 293178 283255 293181
rect 219268 293176 283255 293178
rect 219268 293120 283194 293176
rect 283250 293120 283255 293176
rect 219268 293118 283255 293120
rect 219268 293116 219274 293118
rect 283189 293115 283255 293118
rect 583520 285276 584960 285516
rect 216254 284820 216260 284884
rect 216324 284882 216330 284884
rect 283097 284882 283163 284885
rect 216324 284880 283163 284882
rect 216324 284824 283102 284880
rect 283158 284824 283163 284880
rect 216324 284822 283163 284824
rect 216324 284820 216330 284822
rect 283097 284819 283163 284822
rect 305269 283522 305335 283525
rect 365662 283522 365668 283524
rect 305269 283520 365668 283522
rect 305269 283464 305274 283520
rect 305330 283464 365668 283520
rect 305269 283462 365668 283464
rect 305269 283459 305335 283462
rect 365662 283460 365668 283462
rect 365732 283460 365738 283524
rect 305177 280802 305243 280805
rect 361614 280802 361620 280804
rect 305177 280800 361620 280802
rect 305177 280744 305182 280800
rect 305238 280744 361620 280800
rect 305177 280742 361620 280744
rect 305177 280739 305243 280742
rect 361614 280740 361620 280742
rect 361684 280740 361690 280804
rect -960 279972 480 280212
rect 306649 272506 306715 272509
rect 368422 272506 368428 272508
rect 306649 272504 368428 272506
rect 306649 272448 306654 272504
rect 306710 272448 368428 272504
rect 306649 272446 368428 272448
rect 306649 272443 306715 272446
rect 368422 272444 368428 272446
rect 368492 272444 368498 272508
rect 579981 272234 580047 272237
rect 583520 272234 584960 272324
rect 579981 272232 584960 272234
rect 579981 272176 579986 272232
rect 580042 272176 584960 272232
rect 579981 272174 584960 272176
rect 579981 272171 580047 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3509 267202 3575 267205
rect -960 267200 3575 267202
rect -960 267144 3514 267200
rect 3570 267144 3575 267200
rect -960 267142 3575 267144
rect -960 267052 480 267142
rect 3509 267139 3575 267142
rect 305085 267066 305151 267069
rect 364374 267066 364380 267068
rect 305085 267064 364380 267066
rect 305085 267008 305090 267064
rect 305146 267008 364380 267064
rect 305085 267006 364380 267008
rect 305085 267003 305151 267006
rect 364374 267004 364380 267006
rect 364444 267004 364450 267068
rect 212390 265508 212396 265572
rect 212460 265570 212466 265572
rect 281993 265570 282059 265573
rect 212460 265568 282059 265570
rect 212460 265512 281998 265568
rect 282054 265512 282059 265568
rect 212460 265510 282059 265512
rect 212460 265508 212466 265510
rect 281993 265507 282059 265510
rect 304993 265570 305059 265573
rect 367134 265570 367140 265572
rect 304993 265568 367140 265570
rect 304993 265512 304998 265568
rect 305054 265512 367140 265568
rect 304993 265510 367140 265512
rect 304993 265507 305059 265510
rect 367134 265508 367140 265510
rect 367204 265508 367210 265572
rect 213126 262788 213132 262852
rect 213196 262850 213202 262852
rect 282913 262850 282979 262853
rect 213196 262848 282979 262850
rect 213196 262792 282918 262848
rect 282974 262792 282979 262848
rect 213196 262790 282979 262792
rect 213196 262788 213202 262790
rect 282913 262787 282979 262790
rect 306465 262850 306531 262853
rect 369894 262850 369900 262852
rect 306465 262848 369900 262850
rect 306465 262792 306470 262848
rect 306526 262792 369900 262848
rect 306465 262790 369900 262792
rect 306465 262787 306531 262790
rect 369894 262788 369900 262790
rect 369964 262788 369970 262852
rect 579797 258906 579863 258909
rect 583520 258906 584960 258996
rect 579797 258904 584960 258906
rect 579797 258848 579802 258904
rect 579858 258848 584960 258904
rect 579797 258846 584960 258848
rect 579797 258843 579863 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3509 254146 3575 254149
rect -960 254144 3575 254146
rect -960 254088 3514 254144
rect 3570 254088 3575 254144
rect -960 254086 3575 254088
rect -960 253996 480 254086
rect 3509 254083 3575 254086
rect 303889 250882 303955 250885
rect 362534 250882 362540 250884
rect 303889 250880 362540 250882
rect 303889 250824 303894 250880
rect 303950 250824 362540 250880
rect 303889 250822 362540 250824
rect 303889 250819 303955 250822
rect 362534 250820 362540 250822
rect 362604 250820 362610 250884
rect 304073 250746 304139 250749
rect 363086 250746 363092 250748
rect 304073 250744 363092 250746
rect 304073 250688 304078 250744
rect 304134 250688 363092 250744
rect 304073 250686 363092 250688
rect 304073 250683 304139 250686
rect 363086 250684 363092 250686
rect 363156 250684 363162 250748
rect 302693 250610 302759 250613
rect 363270 250610 363276 250612
rect 302693 250608 363276 250610
rect 302693 250552 302698 250608
rect 302754 250552 363276 250608
rect 302693 250550 363276 250552
rect 302693 250547 302759 250550
rect 363270 250548 363276 250550
rect 363340 250548 363346 250612
rect 302877 250474 302943 250477
rect 363454 250474 363460 250476
rect 302877 250472 363460 250474
rect 302877 250416 302882 250472
rect 302938 250416 363460 250472
rect 302877 250414 363460 250416
rect 302877 250411 302943 250414
rect 363454 250412 363460 250414
rect 363524 250412 363530 250476
rect 303705 248298 303771 248301
rect 360326 248298 360332 248300
rect 303705 248296 360332 248298
rect 303705 248240 303710 248296
rect 303766 248240 360332 248296
rect 303705 248238 360332 248240
rect 303705 248235 303771 248238
rect 360326 248236 360332 248238
rect 360396 248236 360402 248300
rect 298185 248162 298251 248165
rect 364742 248162 364748 248164
rect 298185 248160 364748 248162
rect 298185 248104 298190 248160
rect 298246 248104 364748 248160
rect 298185 248102 364748 248104
rect 298185 248099 298251 248102
rect 364742 248100 364748 248102
rect 364812 248100 364818 248164
rect 296989 248026 297055 248029
rect 364558 248026 364564 248028
rect 296989 248024 364564 248026
rect 296989 247968 296994 248024
rect 297050 247968 364564 248024
rect 296989 247966 364564 247968
rect 296989 247963 297055 247966
rect 364558 247964 364564 247966
rect 364628 247964 364634 248028
rect 323025 247890 323091 247893
rect 483013 247890 483079 247893
rect 323025 247888 483079 247890
rect 323025 247832 323030 247888
rect 323086 247832 483018 247888
rect 483074 247832 483079 247888
rect 323025 247830 483079 247832
rect 323025 247827 323091 247830
rect 483013 247827 483079 247830
rect 328453 247754 328519 247757
rect 520273 247754 520339 247757
rect 328453 247752 520339 247754
rect 328453 247696 328458 247752
rect 328514 247696 520278 247752
rect 520334 247696 520339 247752
rect 328453 247694 520339 247696
rect 328453 247691 328519 247694
rect 520273 247691 520339 247694
rect 334157 247618 334223 247621
rect 557533 247618 557599 247621
rect 334157 247616 557599 247618
rect 334157 247560 334162 247616
rect 334218 247560 557538 247616
rect 557594 247560 557599 247616
rect 334157 247558 557599 247560
rect 334157 247555 334223 247558
rect 557533 247555 557599 247558
rect 303613 246258 303679 246261
rect 368606 246258 368612 246260
rect 303613 246256 368612 246258
rect 303613 246200 303618 246256
rect 303674 246200 368612 246256
rect 303613 246198 368612 246200
rect 303613 246195 303679 246198
rect 368606 246196 368612 246198
rect 368676 246196 368682 246260
rect 302417 245578 302483 245581
rect 359222 245578 359228 245580
rect 302417 245576 359228 245578
rect 302417 245520 302422 245576
rect 302478 245520 359228 245576
rect 302417 245518 359228 245520
rect 302417 245515 302483 245518
rect 359222 245516 359228 245518
rect 359292 245516 359298 245580
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 302233 245442 302299 245445
rect 359038 245442 359044 245444
rect 302233 245440 359044 245442
rect 302233 245384 302238 245440
rect 302294 245384 359044 245440
rect 302233 245382 359044 245384
rect 302233 245379 302299 245382
rect 359038 245380 359044 245382
rect 359108 245380 359114 245444
rect 583520 245428 584960 245518
rect 320173 245306 320239 245309
rect 467833 245306 467899 245309
rect 320173 245304 467899 245306
rect 320173 245248 320178 245304
rect 320234 245248 467838 245304
rect 467894 245248 467899 245304
rect 320173 245246 467899 245248
rect 320173 245243 320239 245246
rect 467833 245243 467899 245246
rect 322933 245170 322999 245173
rect 480253 245170 480319 245173
rect 322933 245168 480319 245170
rect 322933 245112 322938 245168
rect 322994 245112 480258 245168
rect 480314 245112 480319 245168
rect 322933 245110 480319 245112
rect 322933 245107 322999 245110
rect 480253 245107 480319 245110
rect 323117 245034 323183 245037
rect 481725 245034 481791 245037
rect 323117 245032 481791 245034
rect 323117 244976 323122 245032
rect 323178 244976 481730 245032
rect 481786 244976 481791 245032
rect 323117 244974 481791 244976
rect 323117 244971 323183 244974
rect 481725 244971 481791 244974
rect 332593 244898 332659 244901
rect 545113 244898 545179 244901
rect 332593 244896 545179 244898
rect 332593 244840 332598 244896
rect 332654 244840 545118 244896
rect 545174 244840 545179 244896
rect 332593 244838 545179 244840
rect 332593 244835 332659 244838
rect 545113 244835 545179 244838
rect 357893 244354 357959 244357
rect 358670 244354 358676 244356
rect 357893 244352 358676 244354
rect 357893 244296 357898 244352
rect 357954 244296 358676 244352
rect 357893 244294 358676 244296
rect 357893 244291 357959 244294
rect 358670 244292 358676 244294
rect 358740 244292 358746 244356
rect 218421 243538 218487 243541
rect 218646 243538 218652 243540
rect 218421 243536 218652 243538
rect 218421 243480 218426 243536
rect 218482 243480 218652 243536
rect 218421 243478 218652 243480
rect 218421 243475 218487 243478
rect 218646 243476 218652 243478
rect 218716 243476 218722 243540
rect 295425 243538 295491 243541
rect 364926 243538 364932 243540
rect 295425 243536 364932 243538
rect 295425 243480 295430 243536
rect 295486 243480 364932 243536
rect 295425 243478 364932 243480
rect 295425 243475 295491 243478
rect 364926 243476 364932 243478
rect 364996 243476 365002 243540
rect -960 241090 480 241180
rect 3509 241090 3575 241093
rect -960 241088 3575 241090
rect -960 241032 3514 241088
rect 3570 241032 3575 241088
rect -960 241030 3575 241032
rect -960 240940 480 241030
rect 3509 241027 3575 241030
rect 580809 232386 580875 232389
rect 583520 232386 584960 232476
rect 580809 232384 584960 232386
rect 580809 232328 580814 232384
rect 580870 232328 584960 232384
rect 580809 232326 584960 232328
rect 580809 232323 580875 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 579705 219058 579771 219061
rect 583520 219058 584960 219148
rect 579705 219056 584960 219058
rect 579705 219000 579710 219056
rect 579766 219000 584960 219056
rect 579705 218998 584960 219000
rect 579705 218995 579771 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 579613 205730 579679 205733
rect 583520 205730 584960 205820
rect 579613 205728 584960 205730
rect 579613 205672 579618 205728
rect 579674 205672 584960 205728
rect 579613 205670 584960 205672
rect 579613 205667 579679 205670
rect 358077 205594 358143 205597
rect 364926 205594 364932 205596
rect 358077 205592 364932 205594
rect 358077 205536 358082 205592
rect 358138 205536 364932 205592
rect 358077 205534 364932 205536
rect 358077 205531 358143 205534
rect 364926 205532 364932 205534
rect 364996 205532 365002 205596
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3049 201922 3115 201925
rect -960 201920 3115 201922
rect -960 201864 3054 201920
rect 3110 201864 3115 201920
rect -960 201862 3115 201864
rect -960 201772 480 201862
rect 3049 201859 3115 201862
rect 217133 196890 217199 196893
rect 219390 196890 220064 196924
rect 217133 196888 220064 196890
rect 217133 196832 217138 196888
rect 217194 196864 220064 196888
rect 217194 196832 219450 196864
rect 217133 196830 219450 196832
rect 217133 196827 217199 196830
rect 217409 195938 217475 195941
rect 219390 195938 220064 195972
rect 217409 195936 220064 195938
rect 217409 195880 217414 195936
rect 217470 195912 220064 195936
rect 217470 195880 219450 195912
rect 217409 195878 219450 195880
rect 217409 195875 217475 195878
rect 217685 193762 217751 193765
rect 219390 193762 220064 193796
rect 217685 193760 220064 193762
rect 217685 193704 217690 193760
rect 217746 193736 220064 193760
rect 217746 193704 219450 193736
rect 217685 193702 219450 193704
rect 217685 193699 217751 193702
rect 217041 192810 217107 192813
rect 219390 192810 220064 192844
rect 217041 192808 220064 192810
rect 217041 192752 217046 192808
rect 217102 192784 220064 192808
rect 217102 192752 219450 192784
rect 217041 192750 219450 192752
rect 217041 192747 217107 192750
rect 580717 192538 580783 192541
rect 583520 192538 584960 192628
rect 580717 192536 584960 192538
rect 580717 192480 580722 192536
rect 580778 192480 584960 192536
rect 580717 192478 584960 192480
rect 580717 192475 580783 192478
rect 583520 192388 584960 192478
rect 218513 191042 218579 191045
rect 219390 191042 220064 191076
rect 218513 191040 220064 191042
rect 218513 190984 218518 191040
rect 218574 191016 220064 191040
rect 218574 190984 219450 191016
rect 218513 190982 219450 190984
rect 218513 190979 218579 190982
rect 218697 189954 218763 189957
rect 219390 189954 220064 189988
rect 218697 189952 220064 189954
rect 218697 189896 218702 189952
rect 218758 189928 220064 189952
rect 218758 189896 219450 189928
rect 218697 189894 219450 189896
rect 218697 189891 218763 189894
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 216673 188186 216739 188189
rect 219390 188186 220064 188220
rect 216673 188184 220064 188186
rect 216673 188128 216678 188184
rect 216734 188160 220064 188184
rect 216734 188128 219450 188160
rect 216673 188126 219450 188128
rect 216673 188123 216739 188126
rect 579705 179210 579771 179213
rect 583520 179210 584960 179300
rect 579705 179208 584960 179210
rect 579705 179152 579710 179208
rect 579766 179152 584960 179208
rect 579705 179150 584960 179152
rect 579705 179147 579771 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 217593 169962 217659 169965
rect 219390 169962 220064 169996
rect 217593 169960 220064 169962
rect 217593 169904 217598 169960
rect 217654 169936 220064 169960
rect 217654 169904 219450 169936
rect 217593 169902 219450 169904
rect 217593 169899 217659 169902
rect 217225 168330 217291 168333
rect 219390 168330 220064 168364
rect 217225 168328 220064 168330
rect 217225 168272 217230 168328
rect 217286 168304 220064 168328
rect 217286 168272 219450 168304
rect 217225 168270 219450 168272
rect 217225 168267 217291 168270
rect 217777 168058 217843 168061
rect 219390 168058 220064 168092
rect 217777 168056 220064 168058
rect 217777 168000 217782 168056
rect 217838 168032 220064 168056
rect 217838 168000 219450 168032
rect 217777 167998 219450 168000
rect 217777 167995 217843 167998
rect 583520 165882 584960 165972
rect 567150 165822 584960 165882
rect 358486 165684 358492 165748
rect 358556 165746 358562 165748
rect 567150 165746 567210 165822
rect 358556 165686 567210 165746
rect 583520 165732 584960 165822
rect 358556 165684 358562 165686
rect -960 162890 480 162980
rect 214414 162890 214420 162892
rect -960 162830 214420 162890
rect -960 162740 480 162830
rect 214414 162828 214420 162830
rect 214484 162828 214490 162892
rect 238201 159900 238267 159901
rect 239581 159900 239647 159901
rect 241697 159900 241763 159901
rect 273621 159900 273687 159901
rect 276105 159900 276171 159901
rect 278497 159900 278563 159901
rect 293493 159900 293559 159901
rect 238201 159896 238230 159900
rect 238294 159898 238300 159900
rect 238201 159840 238206 159896
rect 238201 159836 238230 159840
rect 238294 159838 238358 159898
rect 239581 159896 239590 159900
rect 239654 159898 239660 159900
rect 239581 159840 239586 159896
rect 238294 159836 238300 159838
rect 239581 159836 239590 159840
rect 239654 159838 239738 159898
rect 241697 159896 241766 159900
rect 241697 159840 241702 159896
rect 241758 159840 241766 159896
rect 239654 159836 239660 159838
rect 241697 159836 241766 159840
rect 241830 159898 241836 159900
rect 273584 159898 273590 159900
rect 241830 159838 241854 159898
rect 273530 159838 273590 159898
rect 273654 159896 273687 159900
rect 276032 159898 276038 159900
rect 273682 159840 273687 159896
rect 241830 159836 241836 159838
rect 273584 159836 273590 159838
rect 273654 159836 273687 159840
rect 276014 159838 276038 159898
rect 276032 159836 276038 159838
rect 276102 159896 276171 159900
rect 278480 159898 278486 159900
rect 276102 159840 276110 159896
rect 276166 159840 276171 159896
rect 276102 159836 276171 159840
rect 278406 159838 278486 159898
rect 278550 159896 278563 159900
rect 293440 159898 293446 159900
rect 278558 159840 278563 159896
rect 278480 159836 278486 159838
rect 278550 159836 278563 159840
rect 293402 159838 293446 159898
rect 293510 159896 293559 159900
rect 293554 159840 293559 159896
rect 293440 159836 293446 159838
rect 293510 159836 293559 159840
rect 238201 159835 238267 159836
rect 239581 159835 239647 159836
rect 241697 159835 241763 159836
rect 273621 159835 273687 159836
rect 276105 159835 276171 159836
rect 278497 159835 278563 159836
rect 293493 159835 293559 159836
rect 295885 159900 295951 159901
rect 303521 159900 303587 159901
rect 295885 159896 295894 159900
rect 295958 159898 295964 159900
rect 303504 159898 303510 159900
rect 295885 159840 295890 159896
rect 295885 159836 295894 159840
rect 295958 159838 296042 159898
rect 303430 159838 303510 159898
rect 303574 159896 303587 159900
rect 303582 159840 303587 159896
rect 295958 159836 295964 159838
rect 303504 159836 303510 159838
rect 303574 159836 303587 159840
rect 295885 159835 295951 159836
rect 303521 159835 303587 159836
rect 310973 159900 311039 159901
rect 313457 159900 313523 159901
rect 310973 159896 310990 159900
rect 311054 159898 311060 159900
rect 313432 159898 313438 159900
rect 310973 159840 310978 159896
rect 310973 159836 310990 159840
rect 311054 159838 311130 159898
rect 313366 159838 313438 159898
rect 313502 159896 313523 159900
rect 313518 159840 313523 159896
rect 311054 159836 311060 159838
rect 313432 159836 313438 159838
rect 313502 159836 313523 159840
rect 310973 159835 311039 159836
rect 313457 159835 313523 159836
rect 298461 159764 298527 159765
rect 298461 159760 298478 159764
rect 298542 159762 298548 159764
rect 298461 159704 298466 159760
rect 298461 159700 298478 159704
rect 298542 159702 298618 159762
rect 298542 159700 298548 159702
rect 298461 159699 298527 159700
rect 255957 159628 256023 159629
rect 265341 159628 265407 159629
rect 271045 159628 271111 159629
rect 255904 159626 255910 159628
rect 255866 159566 255910 159626
rect 255974 159624 256023 159628
rect 265288 159626 265294 159628
rect 256018 159568 256023 159624
rect 255904 159564 255910 159566
rect 255974 159564 256023 159568
rect 265250 159566 265294 159626
rect 265358 159624 265407 159628
rect 271000 159626 271006 159628
rect 265402 159568 265407 159624
rect 265288 159564 265294 159566
rect 265358 159564 265407 159568
rect 270954 159566 271006 159626
rect 271070 159624 271111 159628
rect 271106 159568 271111 159624
rect 271000 159564 271006 159566
rect 271070 159564 271111 159568
rect 255957 159563 256023 159564
rect 265341 159563 265407 159564
rect 271045 159563 271111 159564
rect 261702 159020 261708 159084
rect 261772 159082 261778 159084
rect 364977 159082 365043 159085
rect 261772 159080 365043 159082
rect 261772 159024 364982 159080
rect 365038 159024 365043 159080
rect 261772 159022 365043 159024
rect 261772 159020 261778 159022
rect 364977 159019 365043 159022
rect 260782 158884 260788 158948
rect 260852 158946 260858 158948
rect 364885 158946 364951 158949
rect 260852 158944 364951 158946
rect 260852 158888 364890 158944
rect 364946 158888 364951 158944
rect 260852 158886 364951 158888
rect 260852 158884 260858 158886
rect 364885 158883 364951 158886
rect 244222 158748 244228 158812
rect 244292 158810 244298 158812
rect 364793 158810 364859 158813
rect 244292 158808 364859 158810
rect 244292 158752 364798 158808
rect 364854 158752 364859 158808
rect 244292 158750 364859 158752
rect 244292 158748 244298 158750
rect 364793 158747 364859 158750
rect 368606 158748 368612 158812
rect 368676 158810 368682 158812
rect 369393 158810 369459 158813
rect 368676 158808 369459 158810
rect 368676 158752 369398 158808
rect 369454 158752 369459 158808
rect 368676 158750 369459 158752
rect 368676 158748 368682 158750
rect 369393 158747 369459 158750
rect 218830 158612 218836 158676
rect 218900 158674 218906 158676
rect 220813 158674 220879 158677
rect 218900 158672 220879 158674
rect 218900 158616 220818 158672
rect 220874 158616 220879 158672
rect 218900 158614 220879 158616
rect 218900 158612 218906 158614
rect 220813 158611 220879 158614
rect 240501 158676 240567 158677
rect 248321 158676 248387 158677
rect 250161 158676 250227 158677
rect 251449 158676 251515 158677
rect 254577 158676 254643 158677
rect 256049 158676 256115 158677
rect 257153 158676 257219 158677
rect 258257 158676 258323 158677
rect 258625 158676 258691 158677
rect 259545 158676 259611 158677
rect 261201 158676 261267 158677
rect 262857 158676 262923 158677
rect 263961 158676 264027 158677
rect 265985 158676 266051 158677
rect 240501 158672 240548 158676
rect 240612 158674 240618 158676
rect 248270 158674 248276 158676
rect 240501 158616 240506 158672
rect 240501 158612 240548 158616
rect 240612 158614 240658 158674
rect 248230 158614 248276 158674
rect 248340 158672 248387 158676
rect 250110 158674 250116 158676
rect 248382 158616 248387 158672
rect 240612 158612 240618 158614
rect 248270 158612 248276 158614
rect 248340 158612 248387 158616
rect 250070 158614 250116 158674
rect 250180 158672 250227 158676
rect 251398 158674 251404 158676
rect 250222 158616 250227 158672
rect 250110 158612 250116 158614
rect 250180 158612 250227 158616
rect 251358 158614 251404 158674
rect 251468 158672 251515 158676
rect 254526 158674 254532 158676
rect 251510 158616 251515 158672
rect 251398 158612 251404 158614
rect 251468 158612 251515 158616
rect 254486 158614 254532 158674
rect 254596 158672 254643 158676
rect 255998 158674 256004 158676
rect 254638 158616 254643 158672
rect 254526 158612 254532 158614
rect 254596 158612 254643 158616
rect 255958 158614 256004 158674
rect 256068 158672 256115 158676
rect 257102 158674 257108 158676
rect 256110 158616 256115 158672
rect 255998 158612 256004 158614
rect 256068 158612 256115 158616
rect 257062 158614 257108 158674
rect 257172 158672 257219 158676
rect 258206 158674 258212 158676
rect 257214 158616 257219 158672
rect 257102 158612 257108 158614
rect 257172 158612 257219 158616
rect 258166 158614 258212 158674
rect 258276 158672 258323 158676
rect 258574 158674 258580 158676
rect 258318 158616 258323 158672
rect 258206 158612 258212 158614
rect 258276 158612 258323 158616
rect 258534 158614 258580 158674
rect 258644 158672 258691 158676
rect 259494 158674 259500 158676
rect 258686 158616 258691 158672
rect 258574 158612 258580 158614
rect 258644 158612 258691 158616
rect 259454 158614 259500 158674
rect 259564 158672 259611 158676
rect 261150 158674 261156 158676
rect 259606 158616 259611 158672
rect 259494 158612 259500 158614
rect 259564 158612 259611 158616
rect 261110 158614 261156 158674
rect 261220 158672 261267 158676
rect 262806 158674 262812 158676
rect 261262 158616 261267 158672
rect 261150 158612 261156 158614
rect 261220 158612 261267 158616
rect 262766 158614 262812 158674
rect 262876 158672 262923 158676
rect 263910 158674 263916 158676
rect 262918 158616 262923 158672
rect 262806 158612 262812 158614
rect 262876 158612 262923 158616
rect 263870 158614 263916 158674
rect 263980 158672 264027 158676
rect 265934 158674 265940 158676
rect 264022 158616 264027 158672
rect 263910 158612 263916 158614
rect 263980 158612 264027 158616
rect 265894 158614 265940 158674
rect 266004 158672 266051 158676
rect 266046 158616 266051 158672
rect 265934 158612 265940 158614
rect 266004 158612 266051 158616
rect 266486 158612 266492 158676
rect 266556 158674 266562 158676
rect 266813 158674 266879 158677
rect 267641 158676 267707 158677
rect 268745 158676 268811 158677
rect 269849 158676 269915 158677
rect 271137 158676 271203 158677
rect 272241 158676 272307 158677
rect 267590 158674 267596 158676
rect 266556 158672 266879 158674
rect 266556 158616 266818 158672
rect 266874 158616 266879 158672
rect 266556 158614 266879 158616
rect 267550 158614 267596 158674
rect 267660 158672 267707 158676
rect 268694 158674 268700 158676
rect 267702 158616 267707 158672
rect 266556 158612 266562 158614
rect 240501 158611 240567 158612
rect 248321 158611 248387 158612
rect 250161 158611 250227 158612
rect 251449 158611 251515 158612
rect 254577 158611 254643 158612
rect 256049 158611 256115 158612
rect 257153 158611 257219 158612
rect 258257 158611 258323 158612
rect 258625 158611 258691 158612
rect 259545 158611 259611 158612
rect 261201 158611 261267 158612
rect 262857 158611 262923 158612
rect 263961 158611 264027 158612
rect 265985 158611 266051 158612
rect 266813 158611 266879 158614
rect 267590 158612 267596 158614
rect 267660 158612 267707 158616
rect 268654 158614 268700 158674
rect 268764 158672 268811 158676
rect 269798 158674 269804 158676
rect 268806 158616 268811 158672
rect 268694 158612 268700 158614
rect 268764 158612 268811 158616
rect 269758 158614 269804 158674
rect 269868 158672 269915 158676
rect 271086 158674 271092 158676
rect 269910 158616 269915 158672
rect 269798 158612 269804 158614
rect 269868 158612 269915 158616
rect 271046 158614 271092 158674
rect 271156 158672 271203 158676
rect 272190 158674 272196 158676
rect 271198 158616 271203 158672
rect 271086 158612 271092 158614
rect 271156 158612 271203 158616
rect 272150 158614 272196 158674
rect 272260 158672 272307 158676
rect 272302 158616 272307 158672
rect 272190 158612 272196 158614
rect 272260 158612 272307 158616
rect 273294 158612 273300 158676
rect 273364 158674 273370 158676
rect 274173 158674 274239 158677
rect 274449 158676 274515 158677
rect 275921 158676 275987 158677
rect 281073 158676 281139 158677
rect 291009 158676 291075 158677
rect 300945 158676 301011 158677
rect 308673 158676 308739 158677
rect 274398 158674 274404 158676
rect 273364 158672 274239 158674
rect 273364 158616 274178 158672
rect 274234 158616 274239 158672
rect 273364 158614 274239 158616
rect 274358 158614 274404 158674
rect 274468 158672 274515 158676
rect 275870 158674 275876 158676
rect 274510 158616 274515 158672
rect 273364 158612 273370 158614
rect 267641 158611 267707 158612
rect 268745 158611 268811 158612
rect 269849 158611 269915 158612
rect 271137 158611 271203 158612
rect 272241 158611 272307 158612
rect 274173 158611 274239 158614
rect 274398 158612 274404 158614
rect 274468 158612 274515 158616
rect 275830 158614 275876 158674
rect 275940 158672 275987 158676
rect 281022 158674 281028 158676
rect 275982 158616 275987 158672
rect 275870 158612 275876 158614
rect 275940 158612 275987 158616
rect 280982 158614 281028 158674
rect 281092 158672 281139 158676
rect 290958 158674 290964 158676
rect 281134 158616 281139 158672
rect 281022 158612 281028 158614
rect 281092 158612 281139 158616
rect 290918 158614 290964 158674
rect 291028 158672 291075 158676
rect 300894 158674 300900 158676
rect 291070 158616 291075 158672
rect 290958 158612 290964 158614
rect 291028 158612 291075 158616
rect 300854 158614 300900 158674
rect 300964 158672 301011 158676
rect 308622 158674 308628 158676
rect 301006 158616 301011 158672
rect 300894 158612 300900 158614
rect 300964 158612 301011 158616
rect 308582 158614 308628 158674
rect 308692 158672 308739 158676
rect 308734 158616 308739 158672
rect 308622 158612 308628 158614
rect 308692 158612 308739 158616
rect 320950 158612 320956 158676
rect 321020 158674 321026 158676
rect 321093 158674 321159 158677
rect 323393 158676 323459 158677
rect 325969 158676 326035 158677
rect 323342 158674 323348 158676
rect 321020 158672 321159 158674
rect 321020 158616 321098 158672
rect 321154 158616 321159 158672
rect 321020 158614 321159 158616
rect 323302 158614 323348 158674
rect 323412 158672 323459 158676
rect 325918 158674 325924 158676
rect 323454 158616 323459 158672
rect 321020 158612 321026 158614
rect 274449 158611 274515 158612
rect 275921 158611 275987 158612
rect 281073 158611 281139 158612
rect 291009 158611 291075 158612
rect 300945 158611 301011 158612
rect 308673 158611 308739 158612
rect 321093 158611 321159 158614
rect 323342 158612 323348 158614
rect 323412 158612 323459 158616
rect 325878 158614 325924 158674
rect 325988 158672 326035 158676
rect 326030 158616 326035 158672
rect 325918 158612 325924 158614
rect 325988 158612 326035 158616
rect 323393 158611 323459 158612
rect 325969 158611 326035 158612
rect 219014 158476 219020 158540
rect 219084 158538 219090 158540
rect 224953 158538 225019 158541
rect 219084 158536 225019 158538
rect 219084 158480 224958 158536
rect 225014 158480 225019 158536
rect 219084 158478 225019 158480
rect 219084 158476 219090 158478
rect 224953 158475 225019 158478
rect 236126 158476 236132 158540
rect 236196 158538 236202 158540
rect 359549 158538 359615 158541
rect 236196 158536 359615 158538
rect 236196 158480 359554 158536
rect 359610 158480 359615 158536
rect 236196 158478 359615 158480
rect 236196 158476 236202 158478
rect 359549 158475 359615 158478
rect 216070 158340 216076 158404
rect 216140 158402 216146 158404
rect 223573 158402 223639 158405
rect 216140 158400 223639 158402
rect 216140 158344 223578 158400
rect 223634 158344 223639 158400
rect 216140 158342 223639 158344
rect 216140 158340 216146 158342
rect 223573 158339 223639 158342
rect 248638 158340 248644 158404
rect 248708 158402 248714 158404
rect 368933 158402 368999 158405
rect 248708 158400 368999 158402
rect 248708 158344 368938 158400
rect 368994 158344 368999 158400
rect 248708 158342 368999 158344
rect 248708 158340 248714 158342
rect 368933 158339 368999 158342
rect 217358 158204 217364 158268
rect 217428 158266 217434 158268
rect 231853 158266 231919 158269
rect 217428 158264 231919 158266
rect 217428 158208 231858 158264
rect 231914 158208 231919 158264
rect 217428 158206 231919 158208
rect 217428 158204 217434 158206
rect 231853 158203 231919 158206
rect 243118 158204 243124 158268
rect 243188 158266 243194 158268
rect 362217 158266 362283 158269
rect 243188 158264 362283 158266
rect 243188 158208 362222 158264
rect 362278 158208 362283 158264
rect 243188 158206 362283 158208
rect 243188 158204 243194 158206
rect 362217 158203 362283 158206
rect 217542 158068 217548 158132
rect 217612 158130 217618 158132
rect 238753 158130 238819 158133
rect 217612 158128 238819 158130
rect 217612 158072 238758 158128
rect 238814 158072 238819 158128
rect 217612 158070 238819 158072
rect 217612 158068 217618 158070
rect 238753 158067 238819 158070
rect 250846 158068 250852 158132
rect 250916 158130 250922 158132
rect 251081 158130 251147 158133
rect 250916 158128 251147 158130
rect 250916 158072 251086 158128
rect 251142 158072 251147 158128
rect 250916 158070 251147 158072
rect 250916 158068 250922 158070
rect 251081 158067 251147 158070
rect 276974 158068 276980 158132
rect 277044 158130 277050 158132
rect 277117 158130 277183 158133
rect 278129 158132 278195 158133
rect 278078 158130 278084 158132
rect 277044 158128 277183 158130
rect 277044 158072 277122 158128
rect 277178 158072 277183 158128
rect 277044 158070 277183 158072
rect 278038 158070 278084 158130
rect 278148 158128 278195 158132
rect 278190 158072 278195 158128
rect 277044 158068 277050 158070
rect 277117 158067 277183 158070
rect 278078 158068 278084 158070
rect 278148 158068 278195 158072
rect 279182 158068 279188 158132
rect 279252 158130 279258 158132
rect 279969 158130 280035 158133
rect 279252 158128 280035 158130
rect 279252 158072 279974 158128
rect 280030 158072 280035 158128
rect 279252 158070 280035 158072
rect 279252 158068 279258 158070
rect 278129 158067 278195 158068
rect 279969 158067 280035 158070
rect 353937 158130 354003 158133
rect 358077 158130 358143 158133
rect 353937 158128 358143 158130
rect 353937 158072 353942 158128
rect 353998 158072 358082 158128
rect 358138 158072 358143 158128
rect 353937 158070 358143 158072
rect 353937 158067 354003 158070
rect 358077 158067 358143 158070
rect 216990 157932 216996 157996
rect 217060 157994 217066 157996
rect 251173 157994 251239 157997
rect 252369 157996 252435 157997
rect 252318 157994 252324 157996
rect 217060 157992 251239 157994
rect 217060 157936 251178 157992
rect 251234 157936 251239 157992
rect 217060 157934 251239 157936
rect 252278 157934 252324 157994
rect 252388 157992 252435 157996
rect 252430 157936 252435 157992
rect 217060 157932 217066 157934
rect 251173 157931 251239 157934
rect 252318 157932 252324 157934
rect 252388 157932 252435 157936
rect 253422 157932 253428 157996
rect 253492 157994 253498 157996
rect 253565 157994 253631 157997
rect 253492 157992 253631 157994
rect 253492 157936 253570 157992
rect 253626 157936 253631 157992
rect 253492 157934 253631 157936
rect 253492 157932 253498 157934
rect 252369 157931 252435 157932
rect 253565 157931 253631 157934
rect 268326 157932 268332 157996
rect 268396 157994 268402 157996
rect 268929 157994 268995 157997
rect 268396 157992 268995 157994
rect 268396 157936 268934 157992
rect 268990 157936 268995 157992
rect 268396 157934 268995 157936
rect 268396 157932 268402 157934
rect 268929 157931 268995 157934
rect 354121 157994 354187 157997
rect 358353 157994 358419 157997
rect 354121 157992 358419 157994
rect 354121 157936 354126 157992
rect 354182 157936 358358 157992
rect 358414 157936 358419 157992
rect 354121 157934 358419 157936
rect 354121 157931 354187 157934
rect 358353 157931 358419 157934
rect 214782 157796 214788 157860
rect 214852 157858 214858 157860
rect 219433 157858 219499 157861
rect 214852 157856 219499 157858
rect 214852 157800 219438 157856
rect 219494 157800 219499 157856
rect 214852 157798 219499 157800
rect 214852 157796 214858 157798
rect 219433 157795 219499 157798
rect 283598 157796 283604 157860
rect 283668 157858 283674 157860
rect 283741 157858 283807 157861
rect 283668 157856 283807 157858
rect 283668 157800 283746 157856
rect 283802 157800 283807 157856
rect 283668 157798 283807 157800
rect 283668 157796 283674 157798
rect 283741 157795 283807 157798
rect 285990 157796 285996 157860
rect 286060 157858 286066 157860
rect 286501 157858 286567 157861
rect 286060 157856 286567 157858
rect 286060 157800 286506 157856
rect 286562 157800 286567 157856
rect 286060 157798 286567 157800
rect 286060 157796 286066 157798
rect 286501 157795 286567 157798
rect 237230 157524 237236 157588
rect 237300 157586 237306 157588
rect 362309 157586 362375 157589
rect 237300 157584 362375 157586
rect 237300 157528 362314 157584
rect 362370 157528 362375 157584
rect 237300 157526 362375 157528
rect 237300 157524 237306 157526
rect 362309 157523 362375 157526
rect 253657 157452 253723 157453
rect 245510 157388 245516 157452
rect 245580 157388 245586 157452
rect 246614 157388 246620 157452
rect 246684 157388 246690 157452
rect 247718 157388 247724 157452
rect 247788 157450 247794 157452
rect 253606 157450 253612 157452
rect 247788 157390 248430 157450
rect 253566 157390 253612 157450
rect 253676 157448 253723 157452
rect 253718 157392 253723 157448
rect 247788 157388 247794 157390
rect 245518 157042 245578 157388
rect 246622 157178 246682 157388
rect 248370 157314 248430 157390
rect 253606 157388 253612 157390
rect 253676 157388 253723 157392
rect 263542 157388 263548 157452
rect 263612 157450 263618 157452
rect 263961 157450 264027 157453
rect 288249 157452 288315 157453
rect 306097 157452 306163 157453
rect 315849 157452 315915 157453
rect 318609 157452 318675 157453
rect 288198 157450 288204 157452
rect 263612 157448 264027 157450
rect 263612 157392 263966 157448
rect 264022 157392 264027 157448
rect 263612 157390 264027 157392
rect 288158 157390 288204 157450
rect 288268 157448 288315 157452
rect 306046 157450 306052 157452
rect 288310 157392 288315 157448
rect 263612 157388 263618 157390
rect 253657 157387 253723 157388
rect 263961 157387 264027 157390
rect 288198 157388 288204 157390
rect 288268 157388 288315 157392
rect 306006 157390 306052 157450
rect 306116 157448 306163 157452
rect 315798 157450 315804 157452
rect 306158 157392 306163 157448
rect 306046 157388 306052 157390
rect 306116 157388 306163 157392
rect 315758 157390 315804 157450
rect 315868 157448 315915 157452
rect 318558 157450 318564 157452
rect 315910 157392 315915 157448
rect 315798 157388 315804 157390
rect 315868 157388 315915 157392
rect 318518 157390 318564 157450
rect 318628 157448 318675 157452
rect 318670 157392 318675 157448
rect 318558 157388 318564 157390
rect 318628 157388 318675 157392
rect 360326 157388 360332 157452
rect 360396 157450 360402 157452
rect 360929 157450 360995 157453
rect 360396 157448 360995 157450
rect 360396 157392 360934 157448
rect 360990 157392 360995 157448
rect 360396 157390 360995 157392
rect 360396 157388 360402 157390
rect 288249 157387 288315 157388
rect 306097 157387 306163 157388
rect 315849 157387 315915 157388
rect 318609 157387 318675 157388
rect 360929 157387 360995 157390
rect 362217 157450 362283 157453
rect 362534 157450 362540 157452
rect 362217 157448 362540 157450
rect 362217 157392 362222 157448
rect 362278 157392 362540 157448
rect 362217 157390 362540 157392
rect 362217 157387 362283 157390
rect 362534 157388 362540 157390
rect 362604 157388 362610 157452
rect 368749 157314 368815 157317
rect 248370 157312 368815 157314
rect 248370 157256 368754 157312
rect 368810 157256 368815 157312
rect 248370 157254 368815 157256
rect 368749 157251 368815 157254
rect 365989 157178 366055 157181
rect 246622 157176 366055 157178
rect 246622 157120 365994 157176
rect 366050 157120 366055 157176
rect 246622 157118 366055 157120
rect 365989 157115 366055 157118
rect 362493 157042 362559 157045
rect 245518 157040 362559 157042
rect 245518 156984 362498 157040
rect 362554 156984 362559 157040
rect 245518 156982 362559 156984
rect 362493 156979 362559 156982
rect 217174 155212 217180 155276
rect 217244 155274 217250 155276
rect 251265 155274 251331 155277
rect 217244 155272 251331 155274
rect 217244 155216 251270 155272
rect 251326 155216 251331 155272
rect 217244 155214 251331 155216
rect 217244 155212 217250 155214
rect 251265 155211 251331 155214
rect 580533 152690 580599 152693
rect 583520 152690 584960 152780
rect 580533 152688 584960 152690
rect 580533 152632 580538 152688
rect 580594 152632 584960 152688
rect 580533 152630 584960 152632
rect 580533 152627 580599 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3509 149834 3575 149837
rect -960 149832 3575 149834
rect -960 149776 3514 149832
rect 3570 149776 3575 149832
rect -960 149774 3575 149776
rect -960 149684 480 149774
rect 3509 149771 3575 149774
rect 580625 139362 580691 139365
rect 583520 139362 584960 139452
rect 580625 139360 584960 139362
rect 580625 139304 580630 139360
rect 580686 139304 584960 139360
rect 580625 139302 584960 139304
rect 580625 139299 580691 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 580441 126034 580507 126037
rect 583520 126034 584960 126124
rect 580441 126032 584960 126034
rect 580441 125976 580446 126032
rect 580502 125976 584960 126032
rect 580441 125974 584960 125976
rect 580441 125971 580507 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 583520 112842 584960 112932
rect 583342 112782 584960 112842
rect 583342 112706 583402 112782
rect 583520 112706 584960 112782
rect 583342 112692 584960 112706
rect 583342 112646 583586 112692
rect 358302 111828 358308 111892
rect 358372 111890 358378 111892
rect 583526 111890 583586 112646
rect 358372 111830 583586 111890
rect 358372 111828 358378 111830
rect -960 110666 480 110756
rect -960 110606 6930 110666
rect -960 110516 480 110606
rect 6870 110530 6930 110606
rect 211654 110530 211660 110532
rect 6870 110470 211660 110530
rect 211654 110468 211660 110470
rect 211724 110468 211730 110532
rect 368974 99452 368980 99516
rect 369044 99514 369050 99516
rect 583520 99514 584960 99604
rect 369044 99454 584960 99514
rect 369044 99452 369050 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3509 97610 3575 97613
rect -960 97608 3575 97610
rect -960 97552 3514 97608
rect 3570 97552 3575 97608
rect -960 97550 3575 97552
rect -960 97460 480 97550
rect 3509 97547 3575 97550
rect 583520 86186 584960 86276
rect 583342 86126 584960 86186
rect 583342 86050 583402 86126
rect 583520 86050 584960 86126
rect 583342 86036 584960 86050
rect 583342 85990 583586 86036
rect 360694 85580 360700 85644
rect 360764 85642 360770 85644
rect 583526 85642 583586 85990
rect 360764 85582 583586 85642
rect 360764 85580 360770 85582
rect -960 84690 480 84780
rect 3509 84690 3575 84693
rect -960 84688 3575 84690
rect -960 84632 3514 84688
rect 3570 84632 3575 84688
rect -960 84630 3575 84632
rect -960 84540 480 84630
rect 3509 84627 3575 84630
rect 583520 72994 584960 73084
rect 583342 72934 584960 72994
rect 583342 72858 583402 72934
rect 583520 72858 584960 72934
rect 583342 72844 584960 72858
rect 583342 72798 583586 72844
rect 358118 71844 358124 71908
rect 358188 71906 358194 71908
rect 583526 71906 583586 72798
rect 358188 71846 583586 71906
rect 358188 71844 358194 71846
rect -960 71634 480 71724
rect 3509 71634 3575 71637
rect -960 71632 3575 71634
rect -960 71576 3514 71632
rect 3570 71576 3575 71632
rect -960 71574 3575 71576
rect -960 71484 480 71574
rect 3509 71571 3575 71574
rect 583520 59666 584960 59756
rect 567150 59606 584960 59666
rect 367686 59332 367692 59396
rect 367756 59394 367762 59396
rect 567150 59394 567210 59606
rect 583520 59516 584960 59606
rect 367756 59334 567210 59394
rect 367756 59332 367762 59334
rect -960 58578 480 58668
rect 3509 58578 3575 58581
rect -960 58576 3575 58578
rect -960 58520 3514 58576
rect 3570 58520 3575 58576
rect -960 58518 3575 58520
rect -960 58428 480 58518
rect 3509 58515 3575 58518
rect 583520 46338 584960 46428
rect 583342 46278 584960 46338
rect 583342 46202 583402 46278
rect 583520 46202 584960 46278
rect 583342 46188 584960 46202
rect 583342 46142 583586 46188
rect -960 45522 480 45612
rect 359406 45596 359412 45660
rect 359476 45658 359482 45660
rect 583526 45658 583586 46142
rect 359476 45598 583586 45658
rect 359476 45596 359482 45598
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 580349 33146 580415 33149
rect 583520 33146 584960 33236
rect 580349 33144 584960 33146
rect 580349 33088 580354 33144
rect 580410 33088 584960 33144
rect 580349 33086 584960 33088
rect 580349 33083 580415 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect -960 32406 674 32466
rect -960 32330 480 32406
rect 614 32330 674 32406
rect -960 32316 674 32330
rect 246 32270 674 32316
rect 246 31786 306 32270
rect 215886 31786 215892 31788
rect 246 31726 215892 31786
rect 215886 31724 215892 31726
rect 215956 31724 215962 31788
rect 583520 19818 584960 19908
rect 583342 19758 584960 19818
rect 583342 19682 583402 19758
rect 583520 19682 584960 19758
rect 583342 19668 584960 19682
rect 583342 19622 583586 19668
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 358670 19348 358676 19412
rect 358740 19410 358746 19412
rect 583526 19410 583586 19622
rect 358740 19350 583586 19410
rect 358740 19348 358746 19350
rect 319713 9074 319779 9077
rect 364742 9074 364748 9076
rect 319713 9072 364748 9074
rect 319713 9016 319718 9072
rect 319774 9016 364748 9072
rect 319713 9014 364748 9016
rect 319713 9011 319779 9014
rect 364742 9012 364748 9014
rect 364812 9012 364818 9076
rect 305545 8938 305611 8941
rect 364558 8938 364564 8940
rect 305545 8936 364564 8938
rect 305545 8880 305550 8936
rect 305606 8880 364564 8936
rect 305545 8878 364564 8880
rect 305545 8875 305611 8878
rect 364558 8876 364564 8878
rect 364628 8876 364634 8940
rect 351637 6898 351703 6901
rect 363086 6898 363092 6900
rect 351637 6896 363092 6898
rect 351637 6840 351642 6896
rect 351698 6840 363092 6896
rect 351637 6838 363092 6840
rect 351637 6835 351703 6838
rect 363086 6836 363092 6838
rect 363156 6836 363162 6900
rect 348049 6762 348115 6765
rect 363454 6762 363460 6764
rect 348049 6760 363460 6762
rect 348049 6704 348054 6760
rect 348110 6704 363460 6760
rect 348049 6702 363460 6704
rect 348049 6699 348115 6702
rect 363454 6700 363460 6702
rect 363524 6700 363530 6764
rect 344553 6626 344619 6629
rect 363270 6626 363276 6628
rect 344553 6624 363276 6626
rect -960 6490 480 6580
rect 344553 6568 344558 6624
rect 344614 6568 363276 6624
rect 344553 6566 363276 6568
rect 344553 6563 344619 6566
rect 363270 6564 363276 6566
rect 363340 6564 363346 6628
rect 580257 6626 580323 6629
rect 583520 6626 584960 6716
rect 580257 6624 584960 6626
rect 580257 6568 580262 6624
rect 580318 6568 584960 6624
rect 580257 6566 584960 6568
rect 580257 6563 580323 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 340965 6490 341031 6493
rect 363229 6490 363295 6493
rect 340965 6488 363295 6490
rect 340965 6432 340970 6488
rect 341026 6432 363234 6488
rect 363290 6432 363295 6488
rect 583520 6476 584960 6566
rect 340965 6430 363295 6432
rect 340965 6427 341031 6430
rect 363229 6427 363295 6430
rect 337469 6354 337535 6357
rect 363045 6354 363111 6357
rect 337469 6352 363111 6354
rect 337469 6296 337474 6352
rect 337530 6296 363050 6352
rect 363106 6296 363111 6352
rect 337469 6294 363111 6296
rect 337469 6291 337535 6294
rect 363045 6291 363111 6294
rect 333881 6218 333947 6221
rect 362953 6218 363019 6221
rect 333881 6216 363019 6218
rect 333881 6160 333886 6216
rect 333942 6160 362958 6216
rect 363014 6160 363019 6216
rect 333881 6158 363019 6160
rect 333881 6155 333947 6158
rect 362953 6155 363019 6158
rect 346945 4042 347011 4045
rect 360377 4042 360443 4045
rect 346945 4040 360443 4042
rect 346945 3984 346950 4040
rect 347006 3984 360382 4040
rect 360438 3984 360443 4040
rect 346945 3982 360443 3984
rect 346945 3979 347011 3982
rect 360377 3979 360443 3982
rect 215150 3844 215156 3908
rect 215220 3906 215226 3908
rect 222745 3906 222811 3909
rect 215220 3904 222811 3906
rect 215220 3848 222750 3904
rect 222806 3848 222811 3904
rect 215220 3846 222811 3848
rect 215220 3844 215226 3846
rect 222745 3843 222811 3846
rect 345749 3906 345815 3909
rect 359222 3906 359228 3908
rect 345749 3904 359228 3906
rect 345749 3848 345754 3904
rect 345810 3848 359228 3904
rect 345749 3846 359228 3848
rect 345749 3843 345815 3846
rect 359222 3844 359228 3846
rect 359292 3844 359298 3908
rect 360878 3844 360884 3908
rect 360948 3906 360954 3908
rect 367001 3906 367067 3909
rect 360948 3904 367067 3906
rect 360948 3848 367006 3904
rect 367062 3848 367067 3904
rect 360948 3846 367067 3848
rect 360948 3844 360954 3846
rect 367001 3843 367067 3846
rect 216438 3708 216444 3772
rect 216508 3770 216514 3772
rect 219249 3770 219315 3773
rect 216508 3768 219315 3770
rect 216508 3712 219254 3768
rect 219310 3712 219315 3768
rect 216508 3710 219315 3712
rect 216508 3708 216514 3710
rect 219249 3707 219315 3710
rect 342161 3770 342227 3773
rect 359038 3770 359044 3772
rect 342161 3768 359044 3770
rect 342161 3712 342166 3768
rect 342222 3712 359044 3768
rect 342161 3710 359044 3712
rect 342161 3707 342227 3710
rect 359038 3708 359044 3710
rect 359108 3708 359114 3772
rect 218053 3634 218119 3637
rect 219198 3634 219204 3636
rect 218053 3632 219204 3634
rect 218053 3576 218058 3632
rect 218114 3576 219204 3632
rect 218053 3574 219204 3576
rect 218053 3571 218119 3574
rect 219198 3572 219204 3574
rect 219268 3572 219274 3636
rect 219341 3634 219407 3637
rect 226333 3634 226399 3637
rect 219341 3632 226399 3634
rect 219341 3576 219346 3632
rect 219402 3576 226338 3632
rect 226394 3576 226399 3632
rect 219341 3574 226399 3576
rect 219341 3571 219407 3574
rect 226333 3571 226399 3574
rect 343357 3634 343423 3637
rect 356697 3634 356763 3637
rect 359089 3634 359155 3637
rect 343357 3632 356763 3634
rect 343357 3576 343362 3632
rect 343418 3576 356702 3632
rect 356758 3576 356763 3632
rect 343357 3574 356763 3576
rect 343357 3571 343423 3574
rect 356697 3571 356763 3574
rect 356838 3632 359155 3634
rect 356838 3576 359094 3632
rect 359150 3576 359155 3632
rect 356838 3574 359155 3576
rect 212165 3498 212231 3501
rect 212390 3498 212396 3500
rect 212165 3496 212396 3498
rect 212165 3440 212170 3496
rect 212226 3440 212396 3496
rect 212165 3438 212396 3440
rect 212165 3435 212231 3438
rect 212390 3436 212396 3438
rect 212460 3436 212466 3500
rect 213126 3436 213132 3500
rect 213196 3498 213202 3500
rect 213361 3498 213427 3501
rect 213196 3496 213427 3498
rect 213196 3440 213366 3496
rect 213422 3440 213427 3496
rect 213196 3438 213427 3440
rect 213196 3436 213202 3438
rect 213361 3435 213427 3438
rect 214465 3498 214531 3501
rect 214966 3498 214972 3500
rect 214465 3496 214972 3498
rect 214465 3440 214470 3496
rect 214526 3440 214972 3496
rect 214465 3438 214972 3440
rect 214465 3435 214531 3438
rect 214966 3436 214972 3438
rect 215036 3436 215042 3500
rect 215661 3498 215727 3501
rect 216254 3498 216260 3500
rect 215661 3496 216260 3498
rect 215661 3440 215666 3496
rect 215722 3440 216260 3496
rect 215661 3438 216260 3440
rect 215661 3435 215727 3438
rect 216254 3436 216260 3438
rect 216324 3436 216330 3500
rect 218646 3436 218652 3500
rect 218716 3498 218722 3500
rect 219249 3498 219315 3501
rect 218716 3496 219315 3498
rect 218716 3440 219254 3496
rect 219310 3440 219315 3496
rect 218716 3438 219315 3440
rect 218716 3436 218722 3438
rect 219249 3435 219315 3438
rect 338665 3498 338731 3501
rect 356838 3498 356898 3574
rect 359089 3571 359155 3574
rect 338665 3496 356898 3498
rect 338665 3440 338670 3496
rect 338726 3440 356898 3496
rect 338665 3438 356898 3440
rect 338665 3435 338731 3438
rect 358854 3436 358860 3500
rect 358924 3498 358930 3500
rect 359917 3498 359983 3501
rect 358924 3496 359983 3498
rect 358924 3440 359922 3496
rect 359978 3440 359983 3496
rect 358924 3438 359983 3440
rect 358924 3436 358930 3438
rect 359917 3435 359983 3438
rect 360142 3436 360148 3500
rect 360212 3498 360218 3500
rect 361113 3498 361179 3501
rect 360212 3496 361179 3498
rect 360212 3440 361118 3496
rect 361174 3440 361179 3496
rect 360212 3438 361179 3440
rect 360212 3436 360218 3438
rect 361113 3435 361179 3438
rect 361614 3436 361620 3500
rect 361684 3498 361690 3500
rect 362309 3498 362375 3501
rect 361684 3496 362375 3498
rect 361684 3440 362314 3496
rect 362370 3440 362375 3496
rect 361684 3438 362375 3440
rect 361684 3436 361690 3438
rect 362309 3435 362375 3438
rect 362902 3436 362908 3500
rect 362972 3498 362978 3500
rect 363505 3498 363571 3501
rect 362972 3496 363571 3498
rect 362972 3440 363510 3496
rect 363566 3440 363571 3496
rect 362972 3438 363571 3440
rect 362972 3436 362978 3438
rect 363505 3435 363571 3438
rect 364374 3436 364380 3500
rect 364444 3498 364450 3500
rect 364609 3498 364675 3501
rect 364444 3496 364675 3498
rect 364444 3440 364614 3496
rect 364670 3440 364675 3496
rect 364444 3438 364675 3440
rect 364444 3436 364450 3438
rect 364609 3435 364675 3438
rect 365662 3436 365668 3500
rect 365732 3498 365738 3500
rect 365805 3498 365871 3501
rect 365732 3496 365871 3498
rect 365732 3440 365810 3496
rect 365866 3440 365871 3496
rect 365732 3438 365871 3440
rect 365732 3436 365738 3438
rect 365805 3435 365871 3438
rect 367134 3436 367140 3500
rect 367204 3498 367210 3500
rect 368197 3498 368263 3501
rect 367204 3496 368263 3498
rect 367204 3440 368202 3496
rect 368258 3440 368263 3496
rect 367204 3438 368263 3440
rect 367204 3436 367210 3438
rect 368197 3435 368263 3438
rect 368422 3436 368428 3500
rect 368492 3498 368498 3500
rect 369393 3498 369459 3501
rect 368492 3496 369459 3498
rect 368492 3440 369398 3496
rect 369454 3440 369459 3496
rect 368492 3438 369459 3440
rect 368492 3436 368498 3438
rect 369393 3435 369459 3438
rect 369894 3436 369900 3500
rect 369964 3498 369970 3500
rect 370589 3498 370655 3501
rect 369964 3496 370655 3498
rect 369964 3440 370594 3496
rect 370650 3440 370655 3496
rect 369964 3438 370655 3440
rect 369964 3436 369970 3438
rect 370589 3435 370655 3438
rect 216489 3362 216555 3365
rect 240501 3362 240567 3365
rect 216489 3360 240567 3362
rect 216489 3304 216494 3360
rect 216550 3304 240506 3360
rect 240562 3304 240567 3360
rect 216489 3302 240567 3304
rect 216489 3299 216555 3302
rect 240501 3299 240567 3302
rect 339861 3362 339927 3365
rect 360561 3362 360627 3365
rect 339861 3360 360627 3362
rect 339861 3304 339866 3360
rect 339922 3304 360566 3360
rect 360622 3304 360627 3360
rect 339861 3302 360627 3304
rect 339861 3299 339927 3302
rect 360561 3299 360627 3302
rect 215109 3226 215175 3229
rect 227529 3226 227595 3229
rect 215109 3224 227595 3226
rect 215109 3168 215114 3224
rect 215170 3168 227534 3224
rect 227590 3168 227595 3224
rect 215109 3166 227595 3168
rect 215109 3163 215175 3166
rect 227529 3163 227595 3166
rect 352833 3226 352899 3229
rect 360193 3226 360259 3229
rect 352833 3224 360259 3226
rect 352833 3168 352838 3224
rect 352894 3168 360198 3224
rect 360254 3168 360259 3224
rect 352833 3166 360259 3168
rect 352833 3163 352899 3166
rect 360193 3163 360259 3166
rect 356697 3090 356763 3093
rect 361757 3090 361823 3093
rect 356697 3088 361823 3090
rect 356697 3032 356702 3088
rect 356758 3032 361762 3088
rect 361818 3032 361823 3088
rect 356697 3030 361823 3032
rect 356697 3027 356763 3030
rect 361757 3027 361823 3030
<< via3 >>
rect 238340 477260 238404 477324
rect 268332 477260 268396 477324
rect 241836 477124 241900 477188
rect 306052 477048 306116 477052
rect 306052 476992 306102 477048
rect 306102 476992 306116 477048
rect 306052 476988 306116 476992
rect 320956 476988 321020 477052
rect 239628 476852 239692 476916
rect 240548 476852 240612 476916
rect 281028 476852 281092 476916
rect 308628 476716 308692 476780
rect 248276 476580 248340 476644
rect 258028 476580 258092 476644
rect 263548 476580 263612 476644
rect 313412 476580 313476 476644
rect 253612 476444 253676 476508
rect 259132 476444 259196 476508
rect 273668 476444 273732 476508
rect 318564 476444 318628 476508
rect 236132 476308 236196 476372
rect 244228 476308 244292 476372
rect 246620 476308 246684 476372
rect 250116 476308 250180 476372
rect 251404 476308 251468 476372
rect 255820 476308 255884 476372
rect 259500 476308 259564 476372
rect 261156 476308 261220 476372
rect 265388 476308 265452 476372
rect 266492 476308 266556 476372
rect 270908 476308 270972 476372
rect 273300 476308 273364 476372
rect 276060 476308 276124 476372
rect 278084 476308 278148 476372
rect 303476 476368 303540 476372
rect 303476 476312 303526 476368
rect 303526 476312 303540 476368
rect 303476 476308 303540 476312
rect 323348 476308 323412 476372
rect 237236 476232 237300 476236
rect 237236 476176 237286 476232
rect 237286 476176 237300 476232
rect 237236 476172 237300 476176
rect 243124 476172 243188 476236
rect 245516 476172 245580 476236
rect 247724 476172 247788 476236
rect 248644 476172 248708 476236
rect 250852 476172 250916 476236
rect 252324 476172 252388 476236
rect 253428 476172 253492 476236
rect 254532 476172 254596 476236
rect 256188 476172 256252 476236
rect 257108 476172 257172 476236
rect 260604 476172 260668 476236
rect 261708 476172 261772 476236
rect 262812 476172 262876 476236
rect 263916 476172 263980 476236
rect 265940 476172 266004 476236
rect 267596 476232 267660 476236
rect 267596 476176 267646 476232
rect 267646 476176 267660 476232
rect 267596 476172 267660 476176
rect 268700 476172 268764 476236
rect 269804 476172 269868 476236
rect 271276 476172 271340 476236
rect 272196 476172 272260 476236
rect 274404 476232 274468 476236
rect 274404 476176 274418 476232
rect 274418 476176 274468 476232
rect 274404 476172 274468 476176
rect 275876 476232 275940 476236
rect 275876 476176 275926 476232
rect 275926 476176 275940 476232
rect 275876 476172 275940 476176
rect 276980 476172 277044 476236
rect 278452 476172 278516 476236
rect 279188 476172 279252 476236
rect 283604 476172 283668 476236
rect 285996 476172 286060 476236
rect 288204 476172 288268 476236
rect 290964 476172 291028 476236
rect 293540 476172 293604 476236
rect 295932 476172 295996 476236
rect 298508 476172 298572 476236
rect 300900 476172 300964 476236
rect 311020 476172 311084 476236
rect 315804 476172 315868 476236
rect 326660 476172 326724 476236
rect 368980 436188 369044 436252
rect 367692 436052 367756 436116
rect 214420 435236 214484 435300
rect 215892 435100 215956 435164
rect 211660 434964 211724 435028
rect 360700 434828 360764 434892
rect 359412 434692 359476 434756
rect 358492 432244 358556 432308
rect 358308 432108 358372 432172
rect 358124 431972 358188 432036
rect 245700 431700 245764 431764
rect 245700 430612 245764 430676
rect 232084 374036 232148 374100
rect 232084 372676 232148 372740
rect 232636 309844 232700 309908
rect 234476 309028 234540 309092
rect 234476 308620 234540 308684
rect 232452 308212 232516 308276
rect 219020 306172 219084 306236
rect 218836 306036 218900 306100
rect 217548 305900 217612 305964
rect 217364 305764 217428 305828
rect 216444 303316 216508 303380
rect 214788 303180 214852 303244
rect 216076 303044 216140 303108
rect 215156 302908 215220 302972
rect 362908 302908 362972 302972
rect 216996 302772 217060 302836
rect 214972 301684 215036 301748
rect 217180 301412 217244 301476
rect 169156 301140 169220 301204
rect 358860 300596 358924 300660
rect 169156 297876 169220 297940
rect 360148 295972 360212 296036
rect 360884 294476 360948 294540
rect 219204 293116 219268 293180
rect 216260 284820 216324 284884
rect 365668 283460 365732 283524
rect 361620 280740 361684 280804
rect 368428 272444 368492 272508
rect 364380 267004 364444 267068
rect 212396 265508 212460 265572
rect 367140 265508 367204 265572
rect 213132 262788 213196 262852
rect 369900 262788 369964 262852
rect 362540 250820 362604 250884
rect 363092 250684 363156 250748
rect 363276 250548 363340 250612
rect 363460 250412 363524 250476
rect 360332 248236 360396 248300
rect 364748 248100 364812 248164
rect 364564 247964 364628 248028
rect 368612 246196 368676 246260
rect 359228 245516 359292 245580
rect 359044 245380 359108 245444
rect 358676 244292 358740 244356
rect 218652 243476 218716 243540
rect 364932 243476 364996 243540
rect 364932 205532 364996 205596
rect 358492 165684 358556 165748
rect 214420 162828 214484 162892
rect 238230 159896 238294 159900
rect 238230 159840 238262 159896
rect 238262 159840 238294 159896
rect 238230 159836 238294 159840
rect 239590 159896 239654 159900
rect 239590 159840 239642 159896
rect 239642 159840 239654 159896
rect 239590 159836 239654 159840
rect 241766 159836 241830 159900
rect 273590 159896 273654 159900
rect 273590 159840 273626 159896
rect 273626 159840 273654 159896
rect 273590 159836 273654 159840
rect 276038 159836 276102 159900
rect 278486 159896 278550 159900
rect 278486 159840 278502 159896
rect 278502 159840 278550 159896
rect 278486 159836 278550 159840
rect 293446 159896 293510 159900
rect 293446 159840 293498 159896
rect 293498 159840 293510 159896
rect 293446 159836 293510 159840
rect 295894 159896 295958 159900
rect 295894 159840 295946 159896
rect 295946 159840 295958 159896
rect 295894 159836 295958 159840
rect 303510 159896 303574 159900
rect 303510 159840 303526 159896
rect 303526 159840 303574 159896
rect 303510 159836 303574 159840
rect 310990 159896 311054 159900
rect 310990 159840 311034 159896
rect 311034 159840 311054 159896
rect 310990 159836 311054 159840
rect 313438 159896 313502 159900
rect 313438 159840 313462 159896
rect 313462 159840 313502 159896
rect 313438 159836 313502 159840
rect 298478 159760 298542 159764
rect 298478 159704 298522 159760
rect 298522 159704 298542 159760
rect 298478 159700 298542 159704
rect 255910 159624 255974 159628
rect 255910 159568 255962 159624
rect 255962 159568 255974 159624
rect 255910 159564 255974 159568
rect 265294 159624 265358 159628
rect 265294 159568 265346 159624
rect 265346 159568 265358 159624
rect 265294 159564 265358 159568
rect 271006 159624 271070 159628
rect 271006 159568 271050 159624
rect 271050 159568 271070 159624
rect 271006 159564 271070 159568
rect 261708 159020 261772 159084
rect 260788 158884 260852 158948
rect 244228 158748 244292 158812
rect 368612 158748 368676 158812
rect 218836 158612 218900 158676
rect 240548 158672 240612 158676
rect 240548 158616 240562 158672
rect 240562 158616 240612 158672
rect 240548 158612 240612 158616
rect 248276 158672 248340 158676
rect 248276 158616 248326 158672
rect 248326 158616 248340 158672
rect 248276 158612 248340 158616
rect 250116 158672 250180 158676
rect 250116 158616 250166 158672
rect 250166 158616 250180 158672
rect 250116 158612 250180 158616
rect 251404 158672 251468 158676
rect 251404 158616 251454 158672
rect 251454 158616 251468 158672
rect 251404 158612 251468 158616
rect 254532 158672 254596 158676
rect 254532 158616 254582 158672
rect 254582 158616 254596 158672
rect 254532 158612 254596 158616
rect 256004 158672 256068 158676
rect 256004 158616 256054 158672
rect 256054 158616 256068 158672
rect 256004 158612 256068 158616
rect 257108 158672 257172 158676
rect 257108 158616 257158 158672
rect 257158 158616 257172 158672
rect 257108 158612 257172 158616
rect 258212 158672 258276 158676
rect 258212 158616 258262 158672
rect 258262 158616 258276 158672
rect 258212 158612 258276 158616
rect 258580 158672 258644 158676
rect 258580 158616 258630 158672
rect 258630 158616 258644 158672
rect 258580 158612 258644 158616
rect 259500 158672 259564 158676
rect 259500 158616 259550 158672
rect 259550 158616 259564 158672
rect 259500 158612 259564 158616
rect 261156 158672 261220 158676
rect 261156 158616 261206 158672
rect 261206 158616 261220 158672
rect 261156 158612 261220 158616
rect 262812 158672 262876 158676
rect 262812 158616 262862 158672
rect 262862 158616 262876 158672
rect 262812 158612 262876 158616
rect 263916 158672 263980 158676
rect 263916 158616 263966 158672
rect 263966 158616 263980 158672
rect 263916 158612 263980 158616
rect 265940 158672 266004 158676
rect 265940 158616 265990 158672
rect 265990 158616 266004 158672
rect 265940 158612 266004 158616
rect 266492 158612 266556 158676
rect 267596 158672 267660 158676
rect 267596 158616 267646 158672
rect 267646 158616 267660 158672
rect 267596 158612 267660 158616
rect 268700 158672 268764 158676
rect 268700 158616 268750 158672
rect 268750 158616 268764 158672
rect 268700 158612 268764 158616
rect 269804 158672 269868 158676
rect 269804 158616 269854 158672
rect 269854 158616 269868 158672
rect 269804 158612 269868 158616
rect 271092 158672 271156 158676
rect 271092 158616 271142 158672
rect 271142 158616 271156 158672
rect 271092 158612 271156 158616
rect 272196 158672 272260 158676
rect 272196 158616 272246 158672
rect 272246 158616 272260 158672
rect 272196 158612 272260 158616
rect 273300 158612 273364 158676
rect 274404 158672 274468 158676
rect 274404 158616 274454 158672
rect 274454 158616 274468 158672
rect 274404 158612 274468 158616
rect 275876 158672 275940 158676
rect 275876 158616 275926 158672
rect 275926 158616 275940 158672
rect 275876 158612 275940 158616
rect 281028 158672 281092 158676
rect 281028 158616 281078 158672
rect 281078 158616 281092 158672
rect 281028 158612 281092 158616
rect 290964 158672 291028 158676
rect 290964 158616 291014 158672
rect 291014 158616 291028 158672
rect 290964 158612 291028 158616
rect 300900 158672 300964 158676
rect 300900 158616 300950 158672
rect 300950 158616 300964 158672
rect 300900 158612 300964 158616
rect 308628 158672 308692 158676
rect 308628 158616 308678 158672
rect 308678 158616 308692 158672
rect 308628 158612 308692 158616
rect 320956 158612 321020 158676
rect 323348 158672 323412 158676
rect 323348 158616 323398 158672
rect 323398 158616 323412 158672
rect 323348 158612 323412 158616
rect 325924 158672 325988 158676
rect 325924 158616 325974 158672
rect 325974 158616 325988 158672
rect 325924 158612 325988 158616
rect 219020 158476 219084 158540
rect 236132 158476 236196 158540
rect 216076 158340 216140 158404
rect 248644 158340 248708 158404
rect 217364 158204 217428 158268
rect 243124 158204 243188 158268
rect 217548 158068 217612 158132
rect 250852 158068 250916 158132
rect 276980 158068 277044 158132
rect 278084 158128 278148 158132
rect 278084 158072 278134 158128
rect 278134 158072 278148 158128
rect 278084 158068 278148 158072
rect 279188 158068 279252 158132
rect 216996 157932 217060 157996
rect 252324 157992 252388 157996
rect 252324 157936 252374 157992
rect 252374 157936 252388 157992
rect 252324 157932 252388 157936
rect 253428 157932 253492 157996
rect 268332 157932 268396 157996
rect 214788 157796 214852 157860
rect 283604 157796 283668 157860
rect 285996 157796 286060 157860
rect 237236 157524 237300 157588
rect 245516 157388 245580 157452
rect 246620 157388 246684 157452
rect 247724 157388 247788 157452
rect 253612 157448 253676 157452
rect 253612 157392 253662 157448
rect 253662 157392 253676 157448
rect 253612 157388 253676 157392
rect 263548 157388 263612 157452
rect 288204 157448 288268 157452
rect 288204 157392 288254 157448
rect 288254 157392 288268 157448
rect 288204 157388 288268 157392
rect 306052 157448 306116 157452
rect 306052 157392 306102 157448
rect 306102 157392 306116 157448
rect 306052 157388 306116 157392
rect 315804 157448 315868 157452
rect 315804 157392 315854 157448
rect 315854 157392 315868 157448
rect 315804 157388 315868 157392
rect 318564 157448 318628 157452
rect 318564 157392 318614 157448
rect 318614 157392 318628 157448
rect 318564 157388 318628 157392
rect 360332 157388 360396 157452
rect 362540 157388 362604 157452
rect 217180 155212 217244 155276
rect 358308 111828 358372 111892
rect 211660 110468 211724 110532
rect 368980 99452 369044 99516
rect 360700 85580 360764 85644
rect 358124 71844 358188 71908
rect 367692 59332 367756 59396
rect 359412 45596 359476 45660
rect 215892 31724 215956 31788
rect 358676 19348 358740 19412
rect 364748 9012 364812 9076
rect 364564 8876 364628 8940
rect 363092 6836 363156 6900
rect 363460 6700 363524 6764
rect 363276 6564 363340 6628
rect 215156 3844 215220 3908
rect 359228 3844 359292 3908
rect 360884 3844 360948 3908
rect 216444 3708 216508 3772
rect 359044 3708 359108 3772
rect 219204 3572 219268 3636
rect 212396 3436 212460 3500
rect 213132 3436 213196 3500
rect 214972 3436 215036 3500
rect 216260 3436 216324 3500
rect 218652 3436 218716 3500
rect 358860 3436 358924 3500
rect 360148 3436 360212 3500
rect 361620 3436 361684 3500
rect 362908 3436 362972 3500
rect 364380 3436 364444 3500
rect 365668 3436 365732 3500
rect 367140 3436 367204 3500
rect 368428 3436 368492 3500
rect 369900 3436 369964 3500
<< metal4 >>
rect -9036 711868 -8416 711900
rect -9036 711632 -9004 711868
rect -8768 711632 -8684 711868
rect -8448 711632 -8416 711868
rect -9036 711548 -8416 711632
rect -9036 711312 -9004 711548
rect -8768 711312 -8684 711548
rect -8448 711312 -8416 711548
rect -9036 682954 -8416 711312
rect -9036 682718 -9004 682954
rect -8768 682718 -8684 682954
rect -8448 682718 -8416 682954
rect -9036 682634 -8416 682718
rect -9036 682398 -9004 682634
rect -8768 682398 -8684 682634
rect -8448 682398 -8416 682634
rect -9036 646954 -8416 682398
rect -9036 646718 -9004 646954
rect -8768 646718 -8684 646954
rect -8448 646718 -8416 646954
rect -9036 646634 -8416 646718
rect -9036 646398 -9004 646634
rect -8768 646398 -8684 646634
rect -8448 646398 -8416 646634
rect -9036 610954 -8416 646398
rect -9036 610718 -9004 610954
rect -8768 610718 -8684 610954
rect -8448 610718 -8416 610954
rect -9036 610634 -8416 610718
rect -9036 610398 -9004 610634
rect -8768 610398 -8684 610634
rect -8448 610398 -8416 610634
rect -9036 574954 -8416 610398
rect -9036 574718 -9004 574954
rect -8768 574718 -8684 574954
rect -8448 574718 -8416 574954
rect -9036 574634 -8416 574718
rect -9036 574398 -9004 574634
rect -8768 574398 -8684 574634
rect -8448 574398 -8416 574634
rect -9036 538954 -8416 574398
rect -9036 538718 -9004 538954
rect -8768 538718 -8684 538954
rect -8448 538718 -8416 538954
rect -9036 538634 -8416 538718
rect -9036 538398 -9004 538634
rect -8768 538398 -8684 538634
rect -8448 538398 -8416 538634
rect -9036 502954 -8416 538398
rect -9036 502718 -9004 502954
rect -8768 502718 -8684 502954
rect -8448 502718 -8416 502954
rect -9036 502634 -8416 502718
rect -9036 502398 -9004 502634
rect -8768 502398 -8684 502634
rect -8448 502398 -8416 502634
rect -9036 466954 -8416 502398
rect -9036 466718 -9004 466954
rect -8768 466718 -8684 466954
rect -8448 466718 -8416 466954
rect -9036 466634 -8416 466718
rect -9036 466398 -9004 466634
rect -8768 466398 -8684 466634
rect -8448 466398 -8416 466634
rect -9036 430954 -8416 466398
rect -9036 430718 -9004 430954
rect -8768 430718 -8684 430954
rect -8448 430718 -8416 430954
rect -9036 430634 -8416 430718
rect -9036 430398 -9004 430634
rect -8768 430398 -8684 430634
rect -8448 430398 -8416 430634
rect -9036 394954 -8416 430398
rect -9036 394718 -9004 394954
rect -8768 394718 -8684 394954
rect -8448 394718 -8416 394954
rect -9036 394634 -8416 394718
rect -9036 394398 -9004 394634
rect -8768 394398 -8684 394634
rect -8448 394398 -8416 394634
rect -9036 358954 -8416 394398
rect -9036 358718 -9004 358954
rect -8768 358718 -8684 358954
rect -8448 358718 -8416 358954
rect -9036 358634 -8416 358718
rect -9036 358398 -9004 358634
rect -8768 358398 -8684 358634
rect -8448 358398 -8416 358634
rect -9036 322954 -8416 358398
rect -9036 322718 -9004 322954
rect -8768 322718 -8684 322954
rect -8448 322718 -8416 322954
rect -9036 322634 -8416 322718
rect -9036 322398 -9004 322634
rect -8768 322398 -8684 322634
rect -8448 322398 -8416 322634
rect -9036 286954 -8416 322398
rect -9036 286718 -9004 286954
rect -8768 286718 -8684 286954
rect -8448 286718 -8416 286954
rect -9036 286634 -8416 286718
rect -9036 286398 -9004 286634
rect -8768 286398 -8684 286634
rect -8448 286398 -8416 286634
rect -9036 250954 -8416 286398
rect -9036 250718 -9004 250954
rect -8768 250718 -8684 250954
rect -8448 250718 -8416 250954
rect -9036 250634 -8416 250718
rect -9036 250398 -9004 250634
rect -8768 250398 -8684 250634
rect -8448 250398 -8416 250634
rect -9036 214954 -8416 250398
rect -9036 214718 -9004 214954
rect -8768 214718 -8684 214954
rect -8448 214718 -8416 214954
rect -9036 214634 -8416 214718
rect -9036 214398 -9004 214634
rect -8768 214398 -8684 214634
rect -8448 214398 -8416 214634
rect -9036 178954 -8416 214398
rect -9036 178718 -9004 178954
rect -8768 178718 -8684 178954
rect -8448 178718 -8416 178954
rect -9036 178634 -8416 178718
rect -9036 178398 -9004 178634
rect -8768 178398 -8684 178634
rect -8448 178398 -8416 178634
rect -9036 142954 -8416 178398
rect -9036 142718 -9004 142954
rect -8768 142718 -8684 142954
rect -8448 142718 -8416 142954
rect -9036 142634 -8416 142718
rect -9036 142398 -9004 142634
rect -8768 142398 -8684 142634
rect -8448 142398 -8416 142634
rect -9036 106954 -8416 142398
rect -9036 106718 -9004 106954
rect -8768 106718 -8684 106954
rect -8448 106718 -8416 106954
rect -9036 106634 -8416 106718
rect -9036 106398 -9004 106634
rect -8768 106398 -8684 106634
rect -8448 106398 -8416 106634
rect -9036 70954 -8416 106398
rect -9036 70718 -9004 70954
rect -8768 70718 -8684 70954
rect -8448 70718 -8416 70954
rect -9036 70634 -8416 70718
rect -9036 70398 -9004 70634
rect -8768 70398 -8684 70634
rect -8448 70398 -8416 70634
rect -9036 34954 -8416 70398
rect -9036 34718 -9004 34954
rect -8768 34718 -8684 34954
rect -8448 34718 -8416 34954
rect -9036 34634 -8416 34718
rect -9036 34398 -9004 34634
rect -8768 34398 -8684 34634
rect -8448 34398 -8416 34634
rect -9036 -7376 -8416 34398
rect -8076 710908 -7456 710940
rect -8076 710672 -8044 710908
rect -7808 710672 -7724 710908
rect -7488 710672 -7456 710908
rect -8076 710588 -7456 710672
rect -8076 710352 -8044 710588
rect -7808 710352 -7724 710588
rect -7488 710352 -7456 710588
rect -8076 678454 -7456 710352
rect -8076 678218 -8044 678454
rect -7808 678218 -7724 678454
rect -7488 678218 -7456 678454
rect -8076 678134 -7456 678218
rect -8076 677898 -8044 678134
rect -7808 677898 -7724 678134
rect -7488 677898 -7456 678134
rect -8076 642454 -7456 677898
rect -8076 642218 -8044 642454
rect -7808 642218 -7724 642454
rect -7488 642218 -7456 642454
rect -8076 642134 -7456 642218
rect -8076 641898 -8044 642134
rect -7808 641898 -7724 642134
rect -7488 641898 -7456 642134
rect -8076 606454 -7456 641898
rect -8076 606218 -8044 606454
rect -7808 606218 -7724 606454
rect -7488 606218 -7456 606454
rect -8076 606134 -7456 606218
rect -8076 605898 -8044 606134
rect -7808 605898 -7724 606134
rect -7488 605898 -7456 606134
rect -8076 570454 -7456 605898
rect -8076 570218 -8044 570454
rect -7808 570218 -7724 570454
rect -7488 570218 -7456 570454
rect -8076 570134 -7456 570218
rect -8076 569898 -8044 570134
rect -7808 569898 -7724 570134
rect -7488 569898 -7456 570134
rect -8076 534454 -7456 569898
rect -8076 534218 -8044 534454
rect -7808 534218 -7724 534454
rect -7488 534218 -7456 534454
rect -8076 534134 -7456 534218
rect -8076 533898 -8044 534134
rect -7808 533898 -7724 534134
rect -7488 533898 -7456 534134
rect -8076 498454 -7456 533898
rect -8076 498218 -8044 498454
rect -7808 498218 -7724 498454
rect -7488 498218 -7456 498454
rect -8076 498134 -7456 498218
rect -8076 497898 -8044 498134
rect -7808 497898 -7724 498134
rect -7488 497898 -7456 498134
rect -8076 462454 -7456 497898
rect -8076 462218 -8044 462454
rect -7808 462218 -7724 462454
rect -7488 462218 -7456 462454
rect -8076 462134 -7456 462218
rect -8076 461898 -8044 462134
rect -7808 461898 -7724 462134
rect -7488 461898 -7456 462134
rect -8076 426454 -7456 461898
rect -8076 426218 -8044 426454
rect -7808 426218 -7724 426454
rect -7488 426218 -7456 426454
rect -8076 426134 -7456 426218
rect -8076 425898 -8044 426134
rect -7808 425898 -7724 426134
rect -7488 425898 -7456 426134
rect -8076 390454 -7456 425898
rect -8076 390218 -8044 390454
rect -7808 390218 -7724 390454
rect -7488 390218 -7456 390454
rect -8076 390134 -7456 390218
rect -8076 389898 -8044 390134
rect -7808 389898 -7724 390134
rect -7488 389898 -7456 390134
rect -8076 354454 -7456 389898
rect -8076 354218 -8044 354454
rect -7808 354218 -7724 354454
rect -7488 354218 -7456 354454
rect -8076 354134 -7456 354218
rect -8076 353898 -8044 354134
rect -7808 353898 -7724 354134
rect -7488 353898 -7456 354134
rect -8076 318454 -7456 353898
rect -8076 318218 -8044 318454
rect -7808 318218 -7724 318454
rect -7488 318218 -7456 318454
rect -8076 318134 -7456 318218
rect -8076 317898 -8044 318134
rect -7808 317898 -7724 318134
rect -7488 317898 -7456 318134
rect -8076 282454 -7456 317898
rect -8076 282218 -8044 282454
rect -7808 282218 -7724 282454
rect -7488 282218 -7456 282454
rect -8076 282134 -7456 282218
rect -8076 281898 -8044 282134
rect -7808 281898 -7724 282134
rect -7488 281898 -7456 282134
rect -8076 246454 -7456 281898
rect -8076 246218 -8044 246454
rect -7808 246218 -7724 246454
rect -7488 246218 -7456 246454
rect -8076 246134 -7456 246218
rect -8076 245898 -8044 246134
rect -7808 245898 -7724 246134
rect -7488 245898 -7456 246134
rect -8076 210454 -7456 245898
rect -8076 210218 -8044 210454
rect -7808 210218 -7724 210454
rect -7488 210218 -7456 210454
rect -8076 210134 -7456 210218
rect -8076 209898 -8044 210134
rect -7808 209898 -7724 210134
rect -7488 209898 -7456 210134
rect -8076 174454 -7456 209898
rect -8076 174218 -8044 174454
rect -7808 174218 -7724 174454
rect -7488 174218 -7456 174454
rect -8076 174134 -7456 174218
rect -8076 173898 -8044 174134
rect -7808 173898 -7724 174134
rect -7488 173898 -7456 174134
rect -8076 138454 -7456 173898
rect -8076 138218 -8044 138454
rect -7808 138218 -7724 138454
rect -7488 138218 -7456 138454
rect -8076 138134 -7456 138218
rect -8076 137898 -8044 138134
rect -7808 137898 -7724 138134
rect -7488 137898 -7456 138134
rect -8076 102454 -7456 137898
rect -8076 102218 -8044 102454
rect -7808 102218 -7724 102454
rect -7488 102218 -7456 102454
rect -8076 102134 -7456 102218
rect -8076 101898 -8044 102134
rect -7808 101898 -7724 102134
rect -7488 101898 -7456 102134
rect -8076 66454 -7456 101898
rect -8076 66218 -8044 66454
rect -7808 66218 -7724 66454
rect -7488 66218 -7456 66454
rect -8076 66134 -7456 66218
rect -8076 65898 -8044 66134
rect -7808 65898 -7724 66134
rect -7488 65898 -7456 66134
rect -8076 30454 -7456 65898
rect -8076 30218 -8044 30454
rect -7808 30218 -7724 30454
rect -7488 30218 -7456 30454
rect -8076 30134 -7456 30218
rect -8076 29898 -8044 30134
rect -7808 29898 -7724 30134
rect -7488 29898 -7456 30134
rect -8076 -6416 -7456 29898
rect -7116 709948 -6496 709980
rect -7116 709712 -7084 709948
rect -6848 709712 -6764 709948
rect -6528 709712 -6496 709948
rect -7116 709628 -6496 709712
rect -7116 709392 -7084 709628
rect -6848 709392 -6764 709628
rect -6528 709392 -6496 709628
rect -7116 673954 -6496 709392
rect -7116 673718 -7084 673954
rect -6848 673718 -6764 673954
rect -6528 673718 -6496 673954
rect -7116 673634 -6496 673718
rect -7116 673398 -7084 673634
rect -6848 673398 -6764 673634
rect -6528 673398 -6496 673634
rect -7116 637954 -6496 673398
rect -7116 637718 -7084 637954
rect -6848 637718 -6764 637954
rect -6528 637718 -6496 637954
rect -7116 637634 -6496 637718
rect -7116 637398 -7084 637634
rect -6848 637398 -6764 637634
rect -6528 637398 -6496 637634
rect -7116 601954 -6496 637398
rect -7116 601718 -7084 601954
rect -6848 601718 -6764 601954
rect -6528 601718 -6496 601954
rect -7116 601634 -6496 601718
rect -7116 601398 -7084 601634
rect -6848 601398 -6764 601634
rect -6528 601398 -6496 601634
rect -7116 565954 -6496 601398
rect -7116 565718 -7084 565954
rect -6848 565718 -6764 565954
rect -6528 565718 -6496 565954
rect -7116 565634 -6496 565718
rect -7116 565398 -7084 565634
rect -6848 565398 -6764 565634
rect -6528 565398 -6496 565634
rect -7116 529954 -6496 565398
rect -7116 529718 -7084 529954
rect -6848 529718 -6764 529954
rect -6528 529718 -6496 529954
rect -7116 529634 -6496 529718
rect -7116 529398 -7084 529634
rect -6848 529398 -6764 529634
rect -6528 529398 -6496 529634
rect -7116 493954 -6496 529398
rect -7116 493718 -7084 493954
rect -6848 493718 -6764 493954
rect -6528 493718 -6496 493954
rect -7116 493634 -6496 493718
rect -7116 493398 -7084 493634
rect -6848 493398 -6764 493634
rect -6528 493398 -6496 493634
rect -7116 457954 -6496 493398
rect -7116 457718 -7084 457954
rect -6848 457718 -6764 457954
rect -6528 457718 -6496 457954
rect -7116 457634 -6496 457718
rect -7116 457398 -7084 457634
rect -6848 457398 -6764 457634
rect -6528 457398 -6496 457634
rect -7116 421954 -6496 457398
rect -7116 421718 -7084 421954
rect -6848 421718 -6764 421954
rect -6528 421718 -6496 421954
rect -7116 421634 -6496 421718
rect -7116 421398 -7084 421634
rect -6848 421398 -6764 421634
rect -6528 421398 -6496 421634
rect -7116 385954 -6496 421398
rect -7116 385718 -7084 385954
rect -6848 385718 -6764 385954
rect -6528 385718 -6496 385954
rect -7116 385634 -6496 385718
rect -7116 385398 -7084 385634
rect -6848 385398 -6764 385634
rect -6528 385398 -6496 385634
rect -7116 349954 -6496 385398
rect -7116 349718 -7084 349954
rect -6848 349718 -6764 349954
rect -6528 349718 -6496 349954
rect -7116 349634 -6496 349718
rect -7116 349398 -7084 349634
rect -6848 349398 -6764 349634
rect -6528 349398 -6496 349634
rect -7116 313954 -6496 349398
rect -7116 313718 -7084 313954
rect -6848 313718 -6764 313954
rect -6528 313718 -6496 313954
rect -7116 313634 -6496 313718
rect -7116 313398 -7084 313634
rect -6848 313398 -6764 313634
rect -6528 313398 -6496 313634
rect -7116 277954 -6496 313398
rect -7116 277718 -7084 277954
rect -6848 277718 -6764 277954
rect -6528 277718 -6496 277954
rect -7116 277634 -6496 277718
rect -7116 277398 -7084 277634
rect -6848 277398 -6764 277634
rect -6528 277398 -6496 277634
rect -7116 241954 -6496 277398
rect -7116 241718 -7084 241954
rect -6848 241718 -6764 241954
rect -6528 241718 -6496 241954
rect -7116 241634 -6496 241718
rect -7116 241398 -7084 241634
rect -6848 241398 -6764 241634
rect -6528 241398 -6496 241634
rect -7116 205954 -6496 241398
rect -7116 205718 -7084 205954
rect -6848 205718 -6764 205954
rect -6528 205718 -6496 205954
rect -7116 205634 -6496 205718
rect -7116 205398 -7084 205634
rect -6848 205398 -6764 205634
rect -6528 205398 -6496 205634
rect -7116 169954 -6496 205398
rect -7116 169718 -7084 169954
rect -6848 169718 -6764 169954
rect -6528 169718 -6496 169954
rect -7116 169634 -6496 169718
rect -7116 169398 -7084 169634
rect -6848 169398 -6764 169634
rect -6528 169398 -6496 169634
rect -7116 133954 -6496 169398
rect -7116 133718 -7084 133954
rect -6848 133718 -6764 133954
rect -6528 133718 -6496 133954
rect -7116 133634 -6496 133718
rect -7116 133398 -7084 133634
rect -6848 133398 -6764 133634
rect -6528 133398 -6496 133634
rect -7116 97954 -6496 133398
rect -7116 97718 -7084 97954
rect -6848 97718 -6764 97954
rect -6528 97718 -6496 97954
rect -7116 97634 -6496 97718
rect -7116 97398 -7084 97634
rect -6848 97398 -6764 97634
rect -6528 97398 -6496 97634
rect -7116 61954 -6496 97398
rect -7116 61718 -7084 61954
rect -6848 61718 -6764 61954
rect -6528 61718 -6496 61954
rect -7116 61634 -6496 61718
rect -7116 61398 -7084 61634
rect -6848 61398 -6764 61634
rect -6528 61398 -6496 61634
rect -7116 25954 -6496 61398
rect -7116 25718 -7084 25954
rect -6848 25718 -6764 25954
rect -6528 25718 -6496 25954
rect -7116 25634 -6496 25718
rect -7116 25398 -7084 25634
rect -6848 25398 -6764 25634
rect -6528 25398 -6496 25634
rect -7116 -5456 -6496 25398
rect -6156 708988 -5536 709020
rect -6156 708752 -6124 708988
rect -5888 708752 -5804 708988
rect -5568 708752 -5536 708988
rect -6156 708668 -5536 708752
rect -6156 708432 -6124 708668
rect -5888 708432 -5804 708668
rect -5568 708432 -5536 708668
rect -6156 669454 -5536 708432
rect -6156 669218 -6124 669454
rect -5888 669218 -5804 669454
rect -5568 669218 -5536 669454
rect -6156 669134 -5536 669218
rect -6156 668898 -6124 669134
rect -5888 668898 -5804 669134
rect -5568 668898 -5536 669134
rect -6156 633454 -5536 668898
rect -6156 633218 -6124 633454
rect -5888 633218 -5804 633454
rect -5568 633218 -5536 633454
rect -6156 633134 -5536 633218
rect -6156 632898 -6124 633134
rect -5888 632898 -5804 633134
rect -5568 632898 -5536 633134
rect -6156 597454 -5536 632898
rect -6156 597218 -6124 597454
rect -5888 597218 -5804 597454
rect -5568 597218 -5536 597454
rect -6156 597134 -5536 597218
rect -6156 596898 -6124 597134
rect -5888 596898 -5804 597134
rect -5568 596898 -5536 597134
rect -6156 561454 -5536 596898
rect -6156 561218 -6124 561454
rect -5888 561218 -5804 561454
rect -5568 561218 -5536 561454
rect -6156 561134 -5536 561218
rect -6156 560898 -6124 561134
rect -5888 560898 -5804 561134
rect -5568 560898 -5536 561134
rect -6156 525454 -5536 560898
rect -6156 525218 -6124 525454
rect -5888 525218 -5804 525454
rect -5568 525218 -5536 525454
rect -6156 525134 -5536 525218
rect -6156 524898 -6124 525134
rect -5888 524898 -5804 525134
rect -5568 524898 -5536 525134
rect -6156 489454 -5536 524898
rect -6156 489218 -6124 489454
rect -5888 489218 -5804 489454
rect -5568 489218 -5536 489454
rect -6156 489134 -5536 489218
rect -6156 488898 -6124 489134
rect -5888 488898 -5804 489134
rect -5568 488898 -5536 489134
rect -6156 453454 -5536 488898
rect -6156 453218 -6124 453454
rect -5888 453218 -5804 453454
rect -5568 453218 -5536 453454
rect -6156 453134 -5536 453218
rect -6156 452898 -6124 453134
rect -5888 452898 -5804 453134
rect -5568 452898 -5536 453134
rect -6156 417454 -5536 452898
rect -6156 417218 -6124 417454
rect -5888 417218 -5804 417454
rect -5568 417218 -5536 417454
rect -6156 417134 -5536 417218
rect -6156 416898 -6124 417134
rect -5888 416898 -5804 417134
rect -5568 416898 -5536 417134
rect -6156 381454 -5536 416898
rect -6156 381218 -6124 381454
rect -5888 381218 -5804 381454
rect -5568 381218 -5536 381454
rect -6156 381134 -5536 381218
rect -6156 380898 -6124 381134
rect -5888 380898 -5804 381134
rect -5568 380898 -5536 381134
rect -6156 345454 -5536 380898
rect -6156 345218 -6124 345454
rect -5888 345218 -5804 345454
rect -5568 345218 -5536 345454
rect -6156 345134 -5536 345218
rect -6156 344898 -6124 345134
rect -5888 344898 -5804 345134
rect -5568 344898 -5536 345134
rect -6156 309454 -5536 344898
rect -6156 309218 -6124 309454
rect -5888 309218 -5804 309454
rect -5568 309218 -5536 309454
rect -6156 309134 -5536 309218
rect -6156 308898 -6124 309134
rect -5888 308898 -5804 309134
rect -5568 308898 -5536 309134
rect -6156 273454 -5536 308898
rect -6156 273218 -6124 273454
rect -5888 273218 -5804 273454
rect -5568 273218 -5536 273454
rect -6156 273134 -5536 273218
rect -6156 272898 -6124 273134
rect -5888 272898 -5804 273134
rect -5568 272898 -5536 273134
rect -6156 237454 -5536 272898
rect -6156 237218 -6124 237454
rect -5888 237218 -5804 237454
rect -5568 237218 -5536 237454
rect -6156 237134 -5536 237218
rect -6156 236898 -6124 237134
rect -5888 236898 -5804 237134
rect -5568 236898 -5536 237134
rect -6156 201454 -5536 236898
rect -6156 201218 -6124 201454
rect -5888 201218 -5804 201454
rect -5568 201218 -5536 201454
rect -6156 201134 -5536 201218
rect -6156 200898 -6124 201134
rect -5888 200898 -5804 201134
rect -5568 200898 -5536 201134
rect -6156 165454 -5536 200898
rect -6156 165218 -6124 165454
rect -5888 165218 -5804 165454
rect -5568 165218 -5536 165454
rect -6156 165134 -5536 165218
rect -6156 164898 -6124 165134
rect -5888 164898 -5804 165134
rect -5568 164898 -5536 165134
rect -6156 129454 -5536 164898
rect -6156 129218 -6124 129454
rect -5888 129218 -5804 129454
rect -5568 129218 -5536 129454
rect -6156 129134 -5536 129218
rect -6156 128898 -6124 129134
rect -5888 128898 -5804 129134
rect -5568 128898 -5536 129134
rect -6156 93454 -5536 128898
rect -6156 93218 -6124 93454
rect -5888 93218 -5804 93454
rect -5568 93218 -5536 93454
rect -6156 93134 -5536 93218
rect -6156 92898 -6124 93134
rect -5888 92898 -5804 93134
rect -5568 92898 -5536 93134
rect -6156 57454 -5536 92898
rect -6156 57218 -6124 57454
rect -5888 57218 -5804 57454
rect -5568 57218 -5536 57454
rect -6156 57134 -5536 57218
rect -6156 56898 -6124 57134
rect -5888 56898 -5804 57134
rect -5568 56898 -5536 57134
rect -6156 21454 -5536 56898
rect -6156 21218 -6124 21454
rect -5888 21218 -5804 21454
rect -5568 21218 -5536 21454
rect -6156 21134 -5536 21218
rect -6156 20898 -6124 21134
rect -5888 20898 -5804 21134
rect -5568 20898 -5536 21134
rect -6156 -4496 -5536 20898
rect -5196 708028 -4576 708060
rect -5196 707792 -5164 708028
rect -4928 707792 -4844 708028
rect -4608 707792 -4576 708028
rect -5196 707708 -4576 707792
rect -5196 707472 -5164 707708
rect -4928 707472 -4844 707708
rect -4608 707472 -4576 707708
rect -5196 700954 -4576 707472
rect -5196 700718 -5164 700954
rect -4928 700718 -4844 700954
rect -4608 700718 -4576 700954
rect -5196 700634 -4576 700718
rect -5196 700398 -5164 700634
rect -4928 700398 -4844 700634
rect -4608 700398 -4576 700634
rect -5196 664954 -4576 700398
rect -5196 664718 -5164 664954
rect -4928 664718 -4844 664954
rect -4608 664718 -4576 664954
rect -5196 664634 -4576 664718
rect -5196 664398 -5164 664634
rect -4928 664398 -4844 664634
rect -4608 664398 -4576 664634
rect -5196 628954 -4576 664398
rect -5196 628718 -5164 628954
rect -4928 628718 -4844 628954
rect -4608 628718 -4576 628954
rect -5196 628634 -4576 628718
rect -5196 628398 -5164 628634
rect -4928 628398 -4844 628634
rect -4608 628398 -4576 628634
rect -5196 592954 -4576 628398
rect -5196 592718 -5164 592954
rect -4928 592718 -4844 592954
rect -4608 592718 -4576 592954
rect -5196 592634 -4576 592718
rect -5196 592398 -5164 592634
rect -4928 592398 -4844 592634
rect -4608 592398 -4576 592634
rect -5196 556954 -4576 592398
rect -5196 556718 -5164 556954
rect -4928 556718 -4844 556954
rect -4608 556718 -4576 556954
rect -5196 556634 -4576 556718
rect -5196 556398 -5164 556634
rect -4928 556398 -4844 556634
rect -4608 556398 -4576 556634
rect -5196 520954 -4576 556398
rect -5196 520718 -5164 520954
rect -4928 520718 -4844 520954
rect -4608 520718 -4576 520954
rect -5196 520634 -4576 520718
rect -5196 520398 -5164 520634
rect -4928 520398 -4844 520634
rect -4608 520398 -4576 520634
rect -5196 484954 -4576 520398
rect -5196 484718 -5164 484954
rect -4928 484718 -4844 484954
rect -4608 484718 -4576 484954
rect -5196 484634 -4576 484718
rect -5196 484398 -5164 484634
rect -4928 484398 -4844 484634
rect -4608 484398 -4576 484634
rect -5196 448954 -4576 484398
rect -5196 448718 -5164 448954
rect -4928 448718 -4844 448954
rect -4608 448718 -4576 448954
rect -5196 448634 -4576 448718
rect -5196 448398 -5164 448634
rect -4928 448398 -4844 448634
rect -4608 448398 -4576 448634
rect -5196 412954 -4576 448398
rect -5196 412718 -5164 412954
rect -4928 412718 -4844 412954
rect -4608 412718 -4576 412954
rect -5196 412634 -4576 412718
rect -5196 412398 -5164 412634
rect -4928 412398 -4844 412634
rect -4608 412398 -4576 412634
rect -5196 376954 -4576 412398
rect -5196 376718 -5164 376954
rect -4928 376718 -4844 376954
rect -4608 376718 -4576 376954
rect -5196 376634 -4576 376718
rect -5196 376398 -5164 376634
rect -4928 376398 -4844 376634
rect -4608 376398 -4576 376634
rect -5196 340954 -4576 376398
rect -5196 340718 -5164 340954
rect -4928 340718 -4844 340954
rect -4608 340718 -4576 340954
rect -5196 340634 -4576 340718
rect -5196 340398 -5164 340634
rect -4928 340398 -4844 340634
rect -4608 340398 -4576 340634
rect -5196 304954 -4576 340398
rect -5196 304718 -5164 304954
rect -4928 304718 -4844 304954
rect -4608 304718 -4576 304954
rect -5196 304634 -4576 304718
rect -5196 304398 -5164 304634
rect -4928 304398 -4844 304634
rect -4608 304398 -4576 304634
rect -5196 268954 -4576 304398
rect -5196 268718 -5164 268954
rect -4928 268718 -4844 268954
rect -4608 268718 -4576 268954
rect -5196 268634 -4576 268718
rect -5196 268398 -5164 268634
rect -4928 268398 -4844 268634
rect -4608 268398 -4576 268634
rect -5196 232954 -4576 268398
rect -5196 232718 -5164 232954
rect -4928 232718 -4844 232954
rect -4608 232718 -4576 232954
rect -5196 232634 -4576 232718
rect -5196 232398 -5164 232634
rect -4928 232398 -4844 232634
rect -4608 232398 -4576 232634
rect -5196 196954 -4576 232398
rect -5196 196718 -5164 196954
rect -4928 196718 -4844 196954
rect -4608 196718 -4576 196954
rect -5196 196634 -4576 196718
rect -5196 196398 -5164 196634
rect -4928 196398 -4844 196634
rect -4608 196398 -4576 196634
rect -5196 160954 -4576 196398
rect -5196 160718 -5164 160954
rect -4928 160718 -4844 160954
rect -4608 160718 -4576 160954
rect -5196 160634 -4576 160718
rect -5196 160398 -5164 160634
rect -4928 160398 -4844 160634
rect -4608 160398 -4576 160634
rect -5196 124954 -4576 160398
rect -5196 124718 -5164 124954
rect -4928 124718 -4844 124954
rect -4608 124718 -4576 124954
rect -5196 124634 -4576 124718
rect -5196 124398 -5164 124634
rect -4928 124398 -4844 124634
rect -4608 124398 -4576 124634
rect -5196 88954 -4576 124398
rect -5196 88718 -5164 88954
rect -4928 88718 -4844 88954
rect -4608 88718 -4576 88954
rect -5196 88634 -4576 88718
rect -5196 88398 -5164 88634
rect -4928 88398 -4844 88634
rect -4608 88398 -4576 88634
rect -5196 52954 -4576 88398
rect -5196 52718 -5164 52954
rect -4928 52718 -4844 52954
rect -4608 52718 -4576 52954
rect -5196 52634 -4576 52718
rect -5196 52398 -5164 52634
rect -4928 52398 -4844 52634
rect -4608 52398 -4576 52634
rect -5196 16954 -4576 52398
rect -5196 16718 -5164 16954
rect -4928 16718 -4844 16954
rect -4608 16718 -4576 16954
rect -5196 16634 -4576 16718
rect -5196 16398 -5164 16634
rect -4928 16398 -4844 16634
rect -4608 16398 -4576 16634
rect -5196 -3536 -4576 16398
rect -4236 707068 -3616 707100
rect -4236 706832 -4204 707068
rect -3968 706832 -3884 707068
rect -3648 706832 -3616 707068
rect -4236 706748 -3616 706832
rect -4236 706512 -4204 706748
rect -3968 706512 -3884 706748
rect -3648 706512 -3616 706748
rect -4236 696454 -3616 706512
rect -4236 696218 -4204 696454
rect -3968 696218 -3884 696454
rect -3648 696218 -3616 696454
rect -4236 696134 -3616 696218
rect -4236 695898 -4204 696134
rect -3968 695898 -3884 696134
rect -3648 695898 -3616 696134
rect -4236 660454 -3616 695898
rect -4236 660218 -4204 660454
rect -3968 660218 -3884 660454
rect -3648 660218 -3616 660454
rect -4236 660134 -3616 660218
rect -4236 659898 -4204 660134
rect -3968 659898 -3884 660134
rect -3648 659898 -3616 660134
rect -4236 624454 -3616 659898
rect -4236 624218 -4204 624454
rect -3968 624218 -3884 624454
rect -3648 624218 -3616 624454
rect -4236 624134 -3616 624218
rect -4236 623898 -4204 624134
rect -3968 623898 -3884 624134
rect -3648 623898 -3616 624134
rect -4236 588454 -3616 623898
rect -4236 588218 -4204 588454
rect -3968 588218 -3884 588454
rect -3648 588218 -3616 588454
rect -4236 588134 -3616 588218
rect -4236 587898 -4204 588134
rect -3968 587898 -3884 588134
rect -3648 587898 -3616 588134
rect -4236 552454 -3616 587898
rect -4236 552218 -4204 552454
rect -3968 552218 -3884 552454
rect -3648 552218 -3616 552454
rect -4236 552134 -3616 552218
rect -4236 551898 -4204 552134
rect -3968 551898 -3884 552134
rect -3648 551898 -3616 552134
rect -4236 516454 -3616 551898
rect -4236 516218 -4204 516454
rect -3968 516218 -3884 516454
rect -3648 516218 -3616 516454
rect -4236 516134 -3616 516218
rect -4236 515898 -4204 516134
rect -3968 515898 -3884 516134
rect -3648 515898 -3616 516134
rect -4236 480454 -3616 515898
rect -4236 480218 -4204 480454
rect -3968 480218 -3884 480454
rect -3648 480218 -3616 480454
rect -4236 480134 -3616 480218
rect -4236 479898 -4204 480134
rect -3968 479898 -3884 480134
rect -3648 479898 -3616 480134
rect -4236 444454 -3616 479898
rect -4236 444218 -4204 444454
rect -3968 444218 -3884 444454
rect -3648 444218 -3616 444454
rect -4236 444134 -3616 444218
rect -4236 443898 -4204 444134
rect -3968 443898 -3884 444134
rect -3648 443898 -3616 444134
rect -4236 408454 -3616 443898
rect -4236 408218 -4204 408454
rect -3968 408218 -3884 408454
rect -3648 408218 -3616 408454
rect -4236 408134 -3616 408218
rect -4236 407898 -4204 408134
rect -3968 407898 -3884 408134
rect -3648 407898 -3616 408134
rect -4236 372454 -3616 407898
rect -4236 372218 -4204 372454
rect -3968 372218 -3884 372454
rect -3648 372218 -3616 372454
rect -4236 372134 -3616 372218
rect -4236 371898 -4204 372134
rect -3968 371898 -3884 372134
rect -3648 371898 -3616 372134
rect -4236 336454 -3616 371898
rect -4236 336218 -4204 336454
rect -3968 336218 -3884 336454
rect -3648 336218 -3616 336454
rect -4236 336134 -3616 336218
rect -4236 335898 -4204 336134
rect -3968 335898 -3884 336134
rect -3648 335898 -3616 336134
rect -4236 300454 -3616 335898
rect -4236 300218 -4204 300454
rect -3968 300218 -3884 300454
rect -3648 300218 -3616 300454
rect -4236 300134 -3616 300218
rect -4236 299898 -4204 300134
rect -3968 299898 -3884 300134
rect -3648 299898 -3616 300134
rect -4236 264454 -3616 299898
rect -4236 264218 -4204 264454
rect -3968 264218 -3884 264454
rect -3648 264218 -3616 264454
rect -4236 264134 -3616 264218
rect -4236 263898 -4204 264134
rect -3968 263898 -3884 264134
rect -3648 263898 -3616 264134
rect -4236 228454 -3616 263898
rect -4236 228218 -4204 228454
rect -3968 228218 -3884 228454
rect -3648 228218 -3616 228454
rect -4236 228134 -3616 228218
rect -4236 227898 -4204 228134
rect -3968 227898 -3884 228134
rect -3648 227898 -3616 228134
rect -4236 192454 -3616 227898
rect -4236 192218 -4204 192454
rect -3968 192218 -3884 192454
rect -3648 192218 -3616 192454
rect -4236 192134 -3616 192218
rect -4236 191898 -4204 192134
rect -3968 191898 -3884 192134
rect -3648 191898 -3616 192134
rect -4236 156454 -3616 191898
rect -4236 156218 -4204 156454
rect -3968 156218 -3884 156454
rect -3648 156218 -3616 156454
rect -4236 156134 -3616 156218
rect -4236 155898 -4204 156134
rect -3968 155898 -3884 156134
rect -3648 155898 -3616 156134
rect -4236 120454 -3616 155898
rect -4236 120218 -4204 120454
rect -3968 120218 -3884 120454
rect -3648 120218 -3616 120454
rect -4236 120134 -3616 120218
rect -4236 119898 -4204 120134
rect -3968 119898 -3884 120134
rect -3648 119898 -3616 120134
rect -4236 84454 -3616 119898
rect -4236 84218 -4204 84454
rect -3968 84218 -3884 84454
rect -3648 84218 -3616 84454
rect -4236 84134 -3616 84218
rect -4236 83898 -4204 84134
rect -3968 83898 -3884 84134
rect -3648 83898 -3616 84134
rect -4236 48454 -3616 83898
rect -4236 48218 -4204 48454
rect -3968 48218 -3884 48454
rect -3648 48218 -3616 48454
rect -4236 48134 -3616 48218
rect -4236 47898 -4204 48134
rect -3968 47898 -3884 48134
rect -3648 47898 -3616 48134
rect -4236 12454 -3616 47898
rect -4236 12218 -4204 12454
rect -3968 12218 -3884 12454
rect -3648 12218 -3616 12454
rect -4236 12134 -3616 12218
rect -4236 11898 -4204 12134
rect -3968 11898 -3884 12134
rect -3648 11898 -3616 12134
rect -4236 -2576 -3616 11898
rect -3276 706108 -2656 706140
rect -3276 705872 -3244 706108
rect -3008 705872 -2924 706108
rect -2688 705872 -2656 706108
rect -3276 705788 -2656 705872
rect -3276 705552 -3244 705788
rect -3008 705552 -2924 705788
rect -2688 705552 -2656 705788
rect -3276 691954 -2656 705552
rect -3276 691718 -3244 691954
rect -3008 691718 -2924 691954
rect -2688 691718 -2656 691954
rect -3276 691634 -2656 691718
rect -3276 691398 -3244 691634
rect -3008 691398 -2924 691634
rect -2688 691398 -2656 691634
rect -3276 655954 -2656 691398
rect -3276 655718 -3244 655954
rect -3008 655718 -2924 655954
rect -2688 655718 -2656 655954
rect -3276 655634 -2656 655718
rect -3276 655398 -3244 655634
rect -3008 655398 -2924 655634
rect -2688 655398 -2656 655634
rect -3276 619954 -2656 655398
rect -3276 619718 -3244 619954
rect -3008 619718 -2924 619954
rect -2688 619718 -2656 619954
rect -3276 619634 -2656 619718
rect -3276 619398 -3244 619634
rect -3008 619398 -2924 619634
rect -2688 619398 -2656 619634
rect -3276 583954 -2656 619398
rect -3276 583718 -3244 583954
rect -3008 583718 -2924 583954
rect -2688 583718 -2656 583954
rect -3276 583634 -2656 583718
rect -3276 583398 -3244 583634
rect -3008 583398 -2924 583634
rect -2688 583398 -2656 583634
rect -3276 547954 -2656 583398
rect -3276 547718 -3244 547954
rect -3008 547718 -2924 547954
rect -2688 547718 -2656 547954
rect -3276 547634 -2656 547718
rect -3276 547398 -3244 547634
rect -3008 547398 -2924 547634
rect -2688 547398 -2656 547634
rect -3276 511954 -2656 547398
rect -3276 511718 -3244 511954
rect -3008 511718 -2924 511954
rect -2688 511718 -2656 511954
rect -3276 511634 -2656 511718
rect -3276 511398 -3244 511634
rect -3008 511398 -2924 511634
rect -2688 511398 -2656 511634
rect -3276 475954 -2656 511398
rect -3276 475718 -3244 475954
rect -3008 475718 -2924 475954
rect -2688 475718 -2656 475954
rect -3276 475634 -2656 475718
rect -3276 475398 -3244 475634
rect -3008 475398 -2924 475634
rect -2688 475398 -2656 475634
rect -3276 439954 -2656 475398
rect -3276 439718 -3244 439954
rect -3008 439718 -2924 439954
rect -2688 439718 -2656 439954
rect -3276 439634 -2656 439718
rect -3276 439398 -3244 439634
rect -3008 439398 -2924 439634
rect -2688 439398 -2656 439634
rect -3276 403954 -2656 439398
rect -3276 403718 -3244 403954
rect -3008 403718 -2924 403954
rect -2688 403718 -2656 403954
rect -3276 403634 -2656 403718
rect -3276 403398 -3244 403634
rect -3008 403398 -2924 403634
rect -2688 403398 -2656 403634
rect -3276 367954 -2656 403398
rect -3276 367718 -3244 367954
rect -3008 367718 -2924 367954
rect -2688 367718 -2656 367954
rect -3276 367634 -2656 367718
rect -3276 367398 -3244 367634
rect -3008 367398 -2924 367634
rect -2688 367398 -2656 367634
rect -3276 331954 -2656 367398
rect -3276 331718 -3244 331954
rect -3008 331718 -2924 331954
rect -2688 331718 -2656 331954
rect -3276 331634 -2656 331718
rect -3276 331398 -3244 331634
rect -3008 331398 -2924 331634
rect -2688 331398 -2656 331634
rect -3276 295954 -2656 331398
rect -3276 295718 -3244 295954
rect -3008 295718 -2924 295954
rect -2688 295718 -2656 295954
rect -3276 295634 -2656 295718
rect -3276 295398 -3244 295634
rect -3008 295398 -2924 295634
rect -2688 295398 -2656 295634
rect -3276 259954 -2656 295398
rect -3276 259718 -3244 259954
rect -3008 259718 -2924 259954
rect -2688 259718 -2656 259954
rect -3276 259634 -2656 259718
rect -3276 259398 -3244 259634
rect -3008 259398 -2924 259634
rect -2688 259398 -2656 259634
rect -3276 223954 -2656 259398
rect -3276 223718 -3244 223954
rect -3008 223718 -2924 223954
rect -2688 223718 -2656 223954
rect -3276 223634 -2656 223718
rect -3276 223398 -3244 223634
rect -3008 223398 -2924 223634
rect -2688 223398 -2656 223634
rect -3276 187954 -2656 223398
rect -3276 187718 -3244 187954
rect -3008 187718 -2924 187954
rect -2688 187718 -2656 187954
rect -3276 187634 -2656 187718
rect -3276 187398 -3244 187634
rect -3008 187398 -2924 187634
rect -2688 187398 -2656 187634
rect -3276 151954 -2656 187398
rect -3276 151718 -3244 151954
rect -3008 151718 -2924 151954
rect -2688 151718 -2656 151954
rect -3276 151634 -2656 151718
rect -3276 151398 -3244 151634
rect -3008 151398 -2924 151634
rect -2688 151398 -2656 151634
rect -3276 115954 -2656 151398
rect -3276 115718 -3244 115954
rect -3008 115718 -2924 115954
rect -2688 115718 -2656 115954
rect -3276 115634 -2656 115718
rect -3276 115398 -3244 115634
rect -3008 115398 -2924 115634
rect -2688 115398 -2656 115634
rect -3276 79954 -2656 115398
rect -3276 79718 -3244 79954
rect -3008 79718 -2924 79954
rect -2688 79718 -2656 79954
rect -3276 79634 -2656 79718
rect -3276 79398 -3244 79634
rect -3008 79398 -2924 79634
rect -2688 79398 -2656 79634
rect -3276 43954 -2656 79398
rect -3276 43718 -3244 43954
rect -3008 43718 -2924 43954
rect -2688 43718 -2656 43954
rect -3276 43634 -2656 43718
rect -3276 43398 -3244 43634
rect -3008 43398 -2924 43634
rect -2688 43398 -2656 43634
rect -3276 7954 -2656 43398
rect -3276 7718 -3244 7954
rect -3008 7718 -2924 7954
rect -2688 7718 -2656 7954
rect -3276 7634 -2656 7718
rect -3276 7398 -3244 7634
rect -3008 7398 -2924 7634
rect -2688 7398 -2656 7634
rect -3276 -1616 -2656 7398
rect -2316 705148 -1696 705180
rect -2316 704912 -2284 705148
rect -2048 704912 -1964 705148
rect -1728 704912 -1696 705148
rect -2316 704828 -1696 704912
rect -2316 704592 -2284 704828
rect -2048 704592 -1964 704828
rect -1728 704592 -1696 704828
rect -2316 687454 -1696 704592
rect -2316 687218 -2284 687454
rect -2048 687218 -1964 687454
rect -1728 687218 -1696 687454
rect -2316 687134 -1696 687218
rect -2316 686898 -2284 687134
rect -2048 686898 -1964 687134
rect -1728 686898 -1696 687134
rect -2316 651454 -1696 686898
rect -2316 651218 -2284 651454
rect -2048 651218 -1964 651454
rect -1728 651218 -1696 651454
rect -2316 651134 -1696 651218
rect -2316 650898 -2284 651134
rect -2048 650898 -1964 651134
rect -1728 650898 -1696 651134
rect -2316 615454 -1696 650898
rect -2316 615218 -2284 615454
rect -2048 615218 -1964 615454
rect -1728 615218 -1696 615454
rect -2316 615134 -1696 615218
rect -2316 614898 -2284 615134
rect -2048 614898 -1964 615134
rect -1728 614898 -1696 615134
rect -2316 579454 -1696 614898
rect -2316 579218 -2284 579454
rect -2048 579218 -1964 579454
rect -1728 579218 -1696 579454
rect -2316 579134 -1696 579218
rect -2316 578898 -2284 579134
rect -2048 578898 -1964 579134
rect -1728 578898 -1696 579134
rect -2316 543454 -1696 578898
rect -2316 543218 -2284 543454
rect -2048 543218 -1964 543454
rect -1728 543218 -1696 543454
rect -2316 543134 -1696 543218
rect -2316 542898 -2284 543134
rect -2048 542898 -1964 543134
rect -1728 542898 -1696 543134
rect -2316 507454 -1696 542898
rect -2316 507218 -2284 507454
rect -2048 507218 -1964 507454
rect -1728 507218 -1696 507454
rect -2316 507134 -1696 507218
rect -2316 506898 -2284 507134
rect -2048 506898 -1964 507134
rect -1728 506898 -1696 507134
rect -2316 471454 -1696 506898
rect -2316 471218 -2284 471454
rect -2048 471218 -1964 471454
rect -1728 471218 -1696 471454
rect -2316 471134 -1696 471218
rect -2316 470898 -2284 471134
rect -2048 470898 -1964 471134
rect -1728 470898 -1696 471134
rect -2316 435454 -1696 470898
rect -2316 435218 -2284 435454
rect -2048 435218 -1964 435454
rect -1728 435218 -1696 435454
rect -2316 435134 -1696 435218
rect -2316 434898 -2284 435134
rect -2048 434898 -1964 435134
rect -1728 434898 -1696 435134
rect -2316 399454 -1696 434898
rect -2316 399218 -2284 399454
rect -2048 399218 -1964 399454
rect -1728 399218 -1696 399454
rect -2316 399134 -1696 399218
rect -2316 398898 -2284 399134
rect -2048 398898 -1964 399134
rect -1728 398898 -1696 399134
rect -2316 363454 -1696 398898
rect -2316 363218 -2284 363454
rect -2048 363218 -1964 363454
rect -1728 363218 -1696 363454
rect -2316 363134 -1696 363218
rect -2316 362898 -2284 363134
rect -2048 362898 -1964 363134
rect -1728 362898 -1696 363134
rect -2316 327454 -1696 362898
rect -2316 327218 -2284 327454
rect -2048 327218 -1964 327454
rect -1728 327218 -1696 327454
rect -2316 327134 -1696 327218
rect -2316 326898 -2284 327134
rect -2048 326898 -1964 327134
rect -1728 326898 -1696 327134
rect -2316 291454 -1696 326898
rect -2316 291218 -2284 291454
rect -2048 291218 -1964 291454
rect -1728 291218 -1696 291454
rect -2316 291134 -1696 291218
rect -2316 290898 -2284 291134
rect -2048 290898 -1964 291134
rect -1728 290898 -1696 291134
rect -2316 255454 -1696 290898
rect -2316 255218 -2284 255454
rect -2048 255218 -1964 255454
rect -1728 255218 -1696 255454
rect -2316 255134 -1696 255218
rect -2316 254898 -2284 255134
rect -2048 254898 -1964 255134
rect -1728 254898 -1696 255134
rect -2316 219454 -1696 254898
rect -2316 219218 -2284 219454
rect -2048 219218 -1964 219454
rect -1728 219218 -1696 219454
rect -2316 219134 -1696 219218
rect -2316 218898 -2284 219134
rect -2048 218898 -1964 219134
rect -1728 218898 -1696 219134
rect -2316 183454 -1696 218898
rect -2316 183218 -2284 183454
rect -2048 183218 -1964 183454
rect -1728 183218 -1696 183454
rect -2316 183134 -1696 183218
rect -2316 182898 -2284 183134
rect -2048 182898 -1964 183134
rect -1728 182898 -1696 183134
rect -2316 147454 -1696 182898
rect -2316 147218 -2284 147454
rect -2048 147218 -1964 147454
rect -1728 147218 -1696 147454
rect -2316 147134 -1696 147218
rect -2316 146898 -2284 147134
rect -2048 146898 -1964 147134
rect -1728 146898 -1696 147134
rect -2316 111454 -1696 146898
rect -2316 111218 -2284 111454
rect -2048 111218 -1964 111454
rect -1728 111218 -1696 111454
rect -2316 111134 -1696 111218
rect -2316 110898 -2284 111134
rect -2048 110898 -1964 111134
rect -1728 110898 -1696 111134
rect -2316 75454 -1696 110898
rect -2316 75218 -2284 75454
rect -2048 75218 -1964 75454
rect -1728 75218 -1696 75454
rect -2316 75134 -1696 75218
rect -2316 74898 -2284 75134
rect -2048 74898 -1964 75134
rect -1728 74898 -1696 75134
rect -2316 39454 -1696 74898
rect -2316 39218 -2284 39454
rect -2048 39218 -1964 39454
rect -1728 39218 -1696 39454
rect -2316 39134 -1696 39218
rect -2316 38898 -2284 39134
rect -2048 38898 -1964 39134
rect -1728 38898 -1696 39134
rect -2316 3454 -1696 38898
rect -2316 3218 -2284 3454
rect -2048 3218 -1964 3454
rect -1728 3218 -1696 3454
rect -2316 3134 -1696 3218
rect -2316 2898 -2284 3134
rect -2048 2898 -1964 3134
rect -1728 2898 -1696 3134
rect -2316 -656 -1696 2898
rect -2316 -892 -2284 -656
rect -2048 -892 -1964 -656
rect -1728 -892 -1696 -656
rect -2316 -976 -1696 -892
rect -2316 -1212 -2284 -976
rect -2048 -1212 -1964 -976
rect -1728 -1212 -1696 -976
rect -2316 -1244 -1696 -1212
rect 1794 705148 2414 711900
rect 1794 704912 1826 705148
rect 2062 704912 2146 705148
rect 2382 704912 2414 705148
rect 1794 704828 2414 704912
rect 1794 704592 1826 704828
rect 2062 704592 2146 704828
rect 2382 704592 2414 704828
rect 1794 687454 2414 704592
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -656 2414 2898
rect 1794 -892 1826 -656
rect 2062 -892 2146 -656
rect 2382 -892 2414 -656
rect 1794 -976 2414 -892
rect 1794 -1212 1826 -976
rect 2062 -1212 2146 -976
rect 2382 -1212 2414 -976
rect -3276 -1852 -3244 -1616
rect -3008 -1852 -2924 -1616
rect -2688 -1852 -2656 -1616
rect -3276 -1936 -2656 -1852
rect -3276 -2172 -3244 -1936
rect -3008 -2172 -2924 -1936
rect -2688 -2172 -2656 -1936
rect -3276 -2204 -2656 -2172
rect -4236 -2812 -4204 -2576
rect -3968 -2812 -3884 -2576
rect -3648 -2812 -3616 -2576
rect -4236 -2896 -3616 -2812
rect -4236 -3132 -4204 -2896
rect -3968 -3132 -3884 -2896
rect -3648 -3132 -3616 -2896
rect -4236 -3164 -3616 -3132
rect -5196 -3772 -5164 -3536
rect -4928 -3772 -4844 -3536
rect -4608 -3772 -4576 -3536
rect -5196 -3856 -4576 -3772
rect -5196 -4092 -5164 -3856
rect -4928 -4092 -4844 -3856
rect -4608 -4092 -4576 -3856
rect -5196 -4124 -4576 -4092
rect -6156 -4732 -6124 -4496
rect -5888 -4732 -5804 -4496
rect -5568 -4732 -5536 -4496
rect -6156 -4816 -5536 -4732
rect -6156 -5052 -6124 -4816
rect -5888 -5052 -5804 -4816
rect -5568 -5052 -5536 -4816
rect -6156 -5084 -5536 -5052
rect -7116 -5692 -7084 -5456
rect -6848 -5692 -6764 -5456
rect -6528 -5692 -6496 -5456
rect -7116 -5776 -6496 -5692
rect -7116 -6012 -7084 -5776
rect -6848 -6012 -6764 -5776
rect -6528 -6012 -6496 -5776
rect -7116 -6044 -6496 -6012
rect -8076 -6652 -8044 -6416
rect -7808 -6652 -7724 -6416
rect -7488 -6652 -7456 -6416
rect -8076 -6736 -7456 -6652
rect -8076 -6972 -8044 -6736
rect -7808 -6972 -7724 -6736
rect -7488 -6972 -7456 -6736
rect -8076 -7004 -7456 -6972
rect -9036 -7612 -9004 -7376
rect -8768 -7612 -8684 -7376
rect -8448 -7612 -8416 -7376
rect -9036 -7696 -8416 -7612
rect -9036 -7932 -9004 -7696
rect -8768 -7932 -8684 -7696
rect -8448 -7932 -8416 -7696
rect -9036 -7964 -8416 -7932
rect 1794 -7964 2414 -1212
rect 6294 706108 6914 711900
rect 6294 705872 6326 706108
rect 6562 705872 6646 706108
rect 6882 705872 6914 706108
rect 6294 705788 6914 705872
rect 6294 705552 6326 705788
rect 6562 705552 6646 705788
rect 6882 705552 6914 705788
rect 6294 691954 6914 705552
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1616 6914 7398
rect 6294 -1852 6326 -1616
rect 6562 -1852 6646 -1616
rect 6882 -1852 6914 -1616
rect 6294 -1936 6914 -1852
rect 6294 -2172 6326 -1936
rect 6562 -2172 6646 -1936
rect 6882 -2172 6914 -1936
rect 6294 -7964 6914 -2172
rect 10794 707068 11414 711900
rect 10794 706832 10826 707068
rect 11062 706832 11146 707068
rect 11382 706832 11414 707068
rect 10794 706748 11414 706832
rect 10794 706512 10826 706748
rect 11062 706512 11146 706748
rect 11382 706512 11414 706748
rect 10794 696454 11414 706512
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2576 11414 11898
rect 10794 -2812 10826 -2576
rect 11062 -2812 11146 -2576
rect 11382 -2812 11414 -2576
rect 10794 -2896 11414 -2812
rect 10794 -3132 10826 -2896
rect 11062 -3132 11146 -2896
rect 11382 -3132 11414 -2896
rect 10794 -7964 11414 -3132
rect 15294 708028 15914 711900
rect 15294 707792 15326 708028
rect 15562 707792 15646 708028
rect 15882 707792 15914 708028
rect 15294 707708 15914 707792
rect 15294 707472 15326 707708
rect 15562 707472 15646 707708
rect 15882 707472 15914 707708
rect 15294 700954 15914 707472
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3536 15914 16398
rect 15294 -3772 15326 -3536
rect 15562 -3772 15646 -3536
rect 15882 -3772 15914 -3536
rect 15294 -3856 15914 -3772
rect 15294 -4092 15326 -3856
rect 15562 -4092 15646 -3856
rect 15882 -4092 15914 -3856
rect 15294 -7964 15914 -4092
rect 19794 708988 20414 711900
rect 19794 708752 19826 708988
rect 20062 708752 20146 708988
rect 20382 708752 20414 708988
rect 19794 708668 20414 708752
rect 19794 708432 19826 708668
rect 20062 708432 20146 708668
rect 20382 708432 20414 708668
rect 19794 669454 20414 708432
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4496 20414 20898
rect 19794 -4732 19826 -4496
rect 20062 -4732 20146 -4496
rect 20382 -4732 20414 -4496
rect 19794 -4816 20414 -4732
rect 19794 -5052 19826 -4816
rect 20062 -5052 20146 -4816
rect 20382 -5052 20414 -4816
rect 19794 -7964 20414 -5052
rect 24294 709948 24914 711900
rect 24294 709712 24326 709948
rect 24562 709712 24646 709948
rect 24882 709712 24914 709948
rect 24294 709628 24914 709712
rect 24294 709392 24326 709628
rect 24562 709392 24646 709628
rect 24882 709392 24914 709628
rect 24294 673954 24914 709392
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5456 24914 25398
rect 24294 -5692 24326 -5456
rect 24562 -5692 24646 -5456
rect 24882 -5692 24914 -5456
rect 24294 -5776 24914 -5692
rect 24294 -6012 24326 -5776
rect 24562 -6012 24646 -5776
rect 24882 -6012 24914 -5776
rect 24294 -7964 24914 -6012
rect 28794 710908 29414 711900
rect 28794 710672 28826 710908
rect 29062 710672 29146 710908
rect 29382 710672 29414 710908
rect 28794 710588 29414 710672
rect 28794 710352 28826 710588
rect 29062 710352 29146 710588
rect 29382 710352 29414 710588
rect 28794 678454 29414 710352
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6416 29414 29898
rect 28794 -6652 28826 -6416
rect 29062 -6652 29146 -6416
rect 29382 -6652 29414 -6416
rect 28794 -6736 29414 -6652
rect 28794 -6972 28826 -6736
rect 29062 -6972 29146 -6736
rect 29382 -6972 29414 -6736
rect 28794 -7964 29414 -6972
rect 33294 711868 33914 711900
rect 33294 711632 33326 711868
rect 33562 711632 33646 711868
rect 33882 711632 33914 711868
rect 33294 711548 33914 711632
rect 33294 711312 33326 711548
rect 33562 711312 33646 711548
rect 33882 711312 33914 711548
rect 33294 682954 33914 711312
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7376 33914 34398
rect 33294 -7612 33326 -7376
rect 33562 -7612 33646 -7376
rect 33882 -7612 33914 -7376
rect 33294 -7696 33914 -7612
rect 33294 -7932 33326 -7696
rect 33562 -7932 33646 -7696
rect 33882 -7932 33914 -7696
rect 33294 -7964 33914 -7932
rect 37794 705148 38414 711900
rect 37794 704912 37826 705148
rect 38062 704912 38146 705148
rect 38382 704912 38414 705148
rect 37794 704828 38414 704912
rect 37794 704592 37826 704828
rect 38062 704592 38146 704828
rect 38382 704592 38414 704828
rect 37794 687454 38414 704592
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -656 38414 2898
rect 37794 -892 37826 -656
rect 38062 -892 38146 -656
rect 38382 -892 38414 -656
rect 37794 -976 38414 -892
rect 37794 -1212 37826 -976
rect 38062 -1212 38146 -976
rect 38382 -1212 38414 -976
rect 37794 -7964 38414 -1212
rect 42294 706108 42914 711900
rect 42294 705872 42326 706108
rect 42562 705872 42646 706108
rect 42882 705872 42914 706108
rect 42294 705788 42914 705872
rect 42294 705552 42326 705788
rect 42562 705552 42646 705788
rect 42882 705552 42914 705788
rect 42294 691954 42914 705552
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1616 42914 7398
rect 42294 -1852 42326 -1616
rect 42562 -1852 42646 -1616
rect 42882 -1852 42914 -1616
rect 42294 -1936 42914 -1852
rect 42294 -2172 42326 -1936
rect 42562 -2172 42646 -1936
rect 42882 -2172 42914 -1936
rect 42294 -7964 42914 -2172
rect 46794 707068 47414 711900
rect 46794 706832 46826 707068
rect 47062 706832 47146 707068
rect 47382 706832 47414 707068
rect 46794 706748 47414 706832
rect 46794 706512 46826 706748
rect 47062 706512 47146 706748
rect 47382 706512 47414 706748
rect 46794 696454 47414 706512
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2576 47414 11898
rect 46794 -2812 46826 -2576
rect 47062 -2812 47146 -2576
rect 47382 -2812 47414 -2576
rect 46794 -2896 47414 -2812
rect 46794 -3132 46826 -2896
rect 47062 -3132 47146 -2896
rect 47382 -3132 47414 -2896
rect 46794 -7964 47414 -3132
rect 51294 708028 51914 711900
rect 51294 707792 51326 708028
rect 51562 707792 51646 708028
rect 51882 707792 51914 708028
rect 51294 707708 51914 707792
rect 51294 707472 51326 707708
rect 51562 707472 51646 707708
rect 51882 707472 51914 707708
rect 51294 700954 51914 707472
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3536 51914 16398
rect 51294 -3772 51326 -3536
rect 51562 -3772 51646 -3536
rect 51882 -3772 51914 -3536
rect 51294 -3856 51914 -3772
rect 51294 -4092 51326 -3856
rect 51562 -4092 51646 -3856
rect 51882 -4092 51914 -3856
rect 51294 -7964 51914 -4092
rect 55794 708988 56414 711900
rect 55794 708752 55826 708988
rect 56062 708752 56146 708988
rect 56382 708752 56414 708988
rect 55794 708668 56414 708752
rect 55794 708432 55826 708668
rect 56062 708432 56146 708668
rect 56382 708432 56414 708668
rect 55794 669454 56414 708432
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4496 56414 20898
rect 55794 -4732 55826 -4496
rect 56062 -4732 56146 -4496
rect 56382 -4732 56414 -4496
rect 55794 -4816 56414 -4732
rect 55794 -5052 55826 -4816
rect 56062 -5052 56146 -4816
rect 56382 -5052 56414 -4816
rect 55794 -7964 56414 -5052
rect 60294 709948 60914 711900
rect 60294 709712 60326 709948
rect 60562 709712 60646 709948
rect 60882 709712 60914 709948
rect 60294 709628 60914 709712
rect 60294 709392 60326 709628
rect 60562 709392 60646 709628
rect 60882 709392 60914 709628
rect 60294 673954 60914 709392
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 60294 205954 60914 241398
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5456 60914 25398
rect 60294 -5692 60326 -5456
rect 60562 -5692 60646 -5456
rect 60882 -5692 60914 -5456
rect 60294 -5776 60914 -5692
rect 60294 -6012 60326 -5776
rect 60562 -6012 60646 -5776
rect 60882 -6012 60914 -5776
rect 60294 -7964 60914 -6012
rect 64794 710908 65414 711900
rect 64794 710672 64826 710908
rect 65062 710672 65146 710908
rect 65382 710672 65414 710908
rect 64794 710588 65414 710672
rect 64794 710352 64826 710588
rect 65062 710352 65146 710588
rect 65382 710352 65414 710588
rect 64794 678454 65414 710352
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6416 65414 29898
rect 64794 -6652 64826 -6416
rect 65062 -6652 65146 -6416
rect 65382 -6652 65414 -6416
rect 64794 -6736 65414 -6652
rect 64794 -6972 64826 -6736
rect 65062 -6972 65146 -6736
rect 65382 -6972 65414 -6736
rect 64794 -7964 65414 -6972
rect 69294 711868 69914 711900
rect 69294 711632 69326 711868
rect 69562 711632 69646 711868
rect 69882 711632 69914 711868
rect 69294 711548 69914 711632
rect 69294 711312 69326 711548
rect 69562 711312 69646 711548
rect 69882 711312 69914 711548
rect 69294 682954 69914 711312
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 214954 69914 250398
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7376 69914 34398
rect 69294 -7612 69326 -7376
rect 69562 -7612 69646 -7376
rect 69882 -7612 69914 -7376
rect 69294 -7696 69914 -7612
rect 69294 -7932 69326 -7696
rect 69562 -7932 69646 -7696
rect 69882 -7932 69914 -7696
rect 69294 -7964 69914 -7932
rect 73794 705148 74414 711900
rect 73794 704912 73826 705148
rect 74062 704912 74146 705148
rect 74382 704912 74414 705148
rect 73794 704828 74414 704912
rect 73794 704592 73826 704828
rect 74062 704592 74146 704828
rect 74382 704592 74414 704828
rect 73794 687454 74414 704592
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -656 74414 2898
rect 73794 -892 73826 -656
rect 74062 -892 74146 -656
rect 74382 -892 74414 -656
rect 73794 -976 74414 -892
rect 73794 -1212 73826 -976
rect 74062 -1212 74146 -976
rect 74382 -1212 74414 -976
rect 73794 -7964 74414 -1212
rect 78294 706108 78914 711900
rect 78294 705872 78326 706108
rect 78562 705872 78646 706108
rect 78882 705872 78914 706108
rect 78294 705788 78914 705872
rect 78294 705552 78326 705788
rect 78562 705552 78646 705788
rect 78882 705552 78914 705788
rect 78294 691954 78914 705552
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 223954 78914 259398
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1616 78914 7398
rect 78294 -1852 78326 -1616
rect 78562 -1852 78646 -1616
rect 78882 -1852 78914 -1616
rect 78294 -1936 78914 -1852
rect 78294 -2172 78326 -1936
rect 78562 -2172 78646 -1936
rect 78882 -2172 78914 -1936
rect 78294 -7964 78914 -2172
rect 82794 707068 83414 711900
rect 82794 706832 82826 707068
rect 83062 706832 83146 707068
rect 83382 706832 83414 707068
rect 82794 706748 83414 706832
rect 82794 706512 82826 706748
rect 83062 706512 83146 706748
rect 83382 706512 83414 706748
rect 82794 696454 83414 706512
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 228454 83414 263898
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2576 83414 11898
rect 82794 -2812 82826 -2576
rect 83062 -2812 83146 -2576
rect 83382 -2812 83414 -2576
rect 82794 -2896 83414 -2812
rect 82794 -3132 82826 -2896
rect 83062 -3132 83146 -2896
rect 83382 -3132 83414 -2896
rect 82794 -7964 83414 -3132
rect 87294 708028 87914 711900
rect 87294 707792 87326 708028
rect 87562 707792 87646 708028
rect 87882 707792 87914 708028
rect 87294 707708 87914 707792
rect 87294 707472 87326 707708
rect 87562 707472 87646 707708
rect 87882 707472 87914 707708
rect 87294 700954 87914 707472
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 232954 87914 268398
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3536 87914 16398
rect 87294 -3772 87326 -3536
rect 87562 -3772 87646 -3536
rect 87882 -3772 87914 -3536
rect 87294 -3856 87914 -3772
rect 87294 -4092 87326 -3856
rect 87562 -4092 87646 -3856
rect 87882 -4092 87914 -3856
rect 87294 -7964 87914 -4092
rect 91794 708988 92414 711900
rect 91794 708752 91826 708988
rect 92062 708752 92146 708988
rect 92382 708752 92414 708988
rect 91794 708668 92414 708752
rect 91794 708432 91826 708668
rect 92062 708432 92146 708668
rect 92382 708432 92414 708668
rect 91794 669454 92414 708432
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4496 92414 20898
rect 91794 -4732 91826 -4496
rect 92062 -4732 92146 -4496
rect 92382 -4732 92414 -4496
rect 91794 -4816 92414 -4732
rect 91794 -5052 91826 -4816
rect 92062 -5052 92146 -4816
rect 92382 -5052 92414 -4816
rect 91794 -7964 92414 -5052
rect 96294 709948 96914 711900
rect 96294 709712 96326 709948
rect 96562 709712 96646 709948
rect 96882 709712 96914 709948
rect 96294 709628 96914 709712
rect 96294 709392 96326 709628
rect 96562 709392 96646 709628
rect 96882 709392 96914 709628
rect 96294 673954 96914 709392
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 100794 710908 101414 711900
rect 100794 710672 100826 710908
rect 101062 710672 101146 710908
rect 101382 710672 101414 710908
rect 100794 710588 101414 710672
rect 100794 710352 100826 710588
rect 101062 710352 101146 710588
rect 101382 710352 101414 710588
rect 100794 678454 101414 710352
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 374164 101414 389898
rect 105294 711868 105914 711900
rect 105294 711632 105326 711868
rect 105562 711632 105646 711868
rect 105882 711632 105914 711868
rect 105294 711548 105914 711632
rect 105294 711312 105326 711548
rect 105562 711312 105646 711548
rect 105882 711312 105914 711548
rect 105294 682954 105914 711312
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 374164 105914 394398
rect 109794 705148 110414 711900
rect 109794 704912 109826 705148
rect 110062 704912 110146 705148
rect 110382 704912 110414 705148
rect 109794 704828 110414 704912
rect 109794 704592 109826 704828
rect 110062 704592 110146 704828
rect 110382 704592 110414 704828
rect 109794 687454 110414 704592
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 374164 110414 398898
rect 114294 706108 114914 711900
rect 114294 705872 114326 706108
rect 114562 705872 114646 706108
rect 114882 705872 114914 706108
rect 114294 705788 114914 705872
rect 114294 705552 114326 705788
rect 114562 705552 114646 705788
rect 114882 705552 114914 705788
rect 114294 691954 114914 705552
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 374164 114914 403398
rect 118794 707068 119414 711900
rect 118794 706832 118826 707068
rect 119062 706832 119146 707068
rect 119382 706832 119414 707068
rect 118794 706748 119414 706832
rect 118794 706512 118826 706748
rect 119062 706512 119146 706748
rect 119382 706512 119414 706748
rect 118794 696454 119414 706512
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 374164 119414 407898
rect 123294 708028 123914 711900
rect 123294 707792 123326 708028
rect 123562 707792 123646 708028
rect 123882 707792 123914 708028
rect 123294 707708 123914 707792
rect 123294 707472 123326 707708
rect 123562 707472 123646 707708
rect 123882 707472 123914 707708
rect 123294 700954 123914 707472
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 374164 123914 376398
rect 127794 708988 128414 711900
rect 127794 708752 127826 708988
rect 128062 708752 128146 708988
rect 128382 708752 128414 708988
rect 127794 708668 128414 708752
rect 127794 708432 127826 708668
rect 128062 708432 128146 708668
rect 128382 708432 128414 708668
rect 127794 669454 128414 708432
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 374164 128414 380898
rect 132294 709948 132914 711900
rect 132294 709712 132326 709948
rect 132562 709712 132646 709948
rect 132882 709712 132914 709948
rect 132294 709628 132914 709712
rect 132294 709392 132326 709628
rect 132562 709392 132646 709628
rect 132882 709392 132914 709628
rect 132294 673954 132914 709392
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 374164 132914 385398
rect 136794 710908 137414 711900
rect 136794 710672 136826 710908
rect 137062 710672 137146 710908
rect 137382 710672 137414 710908
rect 136794 710588 137414 710672
rect 136794 710352 136826 710588
rect 137062 710352 137146 710588
rect 137382 710352 137414 710588
rect 136794 678454 137414 710352
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 374164 137414 389898
rect 141294 711868 141914 711900
rect 141294 711632 141326 711868
rect 141562 711632 141646 711868
rect 141882 711632 141914 711868
rect 141294 711548 141914 711632
rect 141294 711312 141326 711548
rect 141562 711312 141646 711548
rect 141882 711312 141914 711548
rect 141294 682954 141914 711312
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 374164 141914 394398
rect 145794 705148 146414 711900
rect 145794 704912 145826 705148
rect 146062 704912 146146 705148
rect 146382 704912 146414 705148
rect 145794 704828 146414 704912
rect 145794 704592 145826 704828
rect 146062 704592 146146 704828
rect 146382 704592 146414 704828
rect 145794 687454 146414 704592
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 374164 146414 398898
rect 150294 706108 150914 711900
rect 150294 705872 150326 706108
rect 150562 705872 150646 706108
rect 150882 705872 150914 706108
rect 150294 705788 150914 705872
rect 150294 705552 150326 705788
rect 150562 705552 150646 705788
rect 150882 705552 150914 705788
rect 150294 691954 150914 705552
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 374164 150914 403398
rect 154794 707068 155414 711900
rect 154794 706832 154826 707068
rect 155062 706832 155146 707068
rect 155382 706832 155414 707068
rect 154794 706748 155414 706832
rect 154794 706512 154826 706748
rect 155062 706512 155146 706748
rect 155382 706512 155414 706748
rect 154794 696454 155414 706512
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 374164 155414 407898
rect 159294 708028 159914 711900
rect 159294 707792 159326 708028
rect 159562 707792 159646 708028
rect 159882 707792 159914 708028
rect 159294 707708 159914 707792
rect 159294 707472 159326 707708
rect 159562 707472 159646 707708
rect 159882 707472 159914 707708
rect 159294 700954 159914 707472
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 374164 159914 376398
rect 163794 708988 164414 711900
rect 163794 708752 163826 708988
rect 164062 708752 164146 708988
rect 164382 708752 164414 708988
rect 163794 708668 164414 708752
rect 163794 708432 163826 708668
rect 164062 708432 164146 708668
rect 164382 708432 164414 708668
rect 163794 669454 164414 708432
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 374164 164414 380898
rect 168294 709948 168914 711900
rect 168294 709712 168326 709948
rect 168562 709712 168646 709948
rect 168882 709712 168914 709948
rect 168294 709628 168914 709712
rect 168294 709392 168326 709628
rect 168562 709392 168646 709628
rect 168882 709392 168914 709628
rect 168294 673954 168914 709392
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 374164 168914 385398
rect 172794 710908 173414 711900
rect 172794 710672 172826 710908
rect 173062 710672 173146 710908
rect 173382 710672 173414 710908
rect 172794 710588 173414 710672
rect 172794 710352 172826 710588
rect 173062 710352 173146 710588
rect 173382 710352 173414 710588
rect 172794 678454 173414 710352
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 119568 367954 119888 367986
rect 119568 367718 119610 367954
rect 119846 367718 119888 367954
rect 119568 367634 119888 367718
rect 119568 367398 119610 367634
rect 119846 367398 119888 367634
rect 119568 367366 119888 367398
rect 150288 367954 150608 367986
rect 150288 367718 150330 367954
rect 150566 367718 150608 367954
rect 150288 367634 150608 367718
rect 150288 367398 150330 367634
rect 150566 367398 150608 367634
rect 150288 367366 150608 367398
rect 104208 363454 104528 363486
rect 104208 363218 104250 363454
rect 104486 363218 104528 363454
rect 104208 363134 104528 363218
rect 104208 362898 104250 363134
rect 104486 362898 104528 363134
rect 104208 362866 104528 362898
rect 134928 363454 135248 363486
rect 134928 363218 134970 363454
rect 135206 363218 135248 363454
rect 134928 363134 135248 363218
rect 134928 362898 134970 363134
rect 135206 362898 135248 363134
rect 134928 362866 135248 362898
rect 165648 363454 165968 363486
rect 165648 363218 165690 363454
rect 165926 363218 165968 363454
rect 165648 363134 165968 363218
rect 165648 362898 165690 363134
rect 165926 362898 165968 363134
rect 165648 362866 165968 362898
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 119568 331954 119888 331986
rect 119568 331718 119610 331954
rect 119846 331718 119888 331954
rect 119568 331634 119888 331718
rect 119568 331398 119610 331634
rect 119846 331398 119888 331634
rect 119568 331366 119888 331398
rect 150288 331954 150608 331986
rect 150288 331718 150330 331954
rect 150566 331718 150608 331954
rect 150288 331634 150608 331718
rect 150288 331398 150330 331634
rect 150566 331398 150608 331634
rect 150288 331366 150608 331398
rect 104208 327454 104528 327486
rect 104208 327218 104250 327454
rect 104486 327218 104528 327454
rect 104208 327134 104528 327218
rect 104208 326898 104250 327134
rect 104486 326898 104528 327134
rect 104208 326866 104528 326898
rect 134928 327454 135248 327486
rect 134928 327218 134970 327454
rect 135206 327218 135248 327454
rect 134928 327134 135248 327218
rect 134928 326898 134970 327134
rect 135206 326898 135248 327134
rect 134928 326866 135248 326898
rect 165648 327454 165968 327486
rect 165648 327218 165690 327454
rect 165926 327218 165968 327454
rect 165648 327134 165968 327218
rect 165648 326898 165690 327134
rect 165926 326898 165968 327134
rect 165648 326866 165968 326898
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 169155 301204 169221 301205
rect 169155 301140 169156 301204
rect 169220 301140 169221 301204
rect 169155 301139 169221 301140
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 241954 96914 277398
rect 96294 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 96914 241954
rect 96294 241634 96914 241718
rect 96294 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 96914 241634
rect 96294 205954 96914 241398
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5456 96914 25398
rect 96294 -5692 96326 -5456
rect 96562 -5692 96646 -5456
rect 96882 -5692 96914 -5456
rect 96294 -5776 96914 -5692
rect 96294 -6012 96326 -5776
rect 96562 -6012 96646 -5776
rect 96882 -6012 96914 -5776
rect 96294 -7964 96914 -6012
rect 100794 282454 101414 298000
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 246454 101414 281898
rect 100794 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 101414 246454
rect 100794 246134 101414 246218
rect 100794 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 101414 246134
rect 100794 210454 101414 245898
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 100794 174454 101414 209898
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 138454 101414 173898
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6416 101414 29898
rect 100794 -6652 100826 -6416
rect 101062 -6652 101146 -6416
rect 101382 -6652 101414 -6416
rect 100794 -6736 101414 -6652
rect 100794 -6972 100826 -6736
rect 101062 -6972 101146 -6736
rect 101382 -6972 101414 -6736
rect 100794 -7964 101414 -6972
rect 105294 286954 105914 298000
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 214954 105914 250398
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 105294 142954 105914 178398
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7376 105914 34398
rect 105294 -7612 105326 -7376
rect 105562 -7612 105646 -7376
rect 105882 -7612 105914 -7376
rect 105294 -7696 105914 -7612
rect 105294 -7932 105326 -7696
rect 105562 -7932 105646 -7696
rect 105882 -7932 105914 -7696
rect 105294 -7964 105914 -7932
rect 109794 291454 110414 298000
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -656 110414 2898
rect 109794 -892 109826 -656
rect 110062 -892 110146 -656
rect 110382 -892 110414 -656
rect 109794 -976 110414 -892
rect 109794 -1212 109826 -976
rect 110062 -1212 110146 -976
rect 110382 -1212 110414 -976
rect 109794 -7964 110414 -1212
rect 114294 295954 114914 298000
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 259954 114914 295398
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 223954 114914 259398
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 151954 114914 187398
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114294 115954 114914 151398
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1616 114914 7398
rect 114294 -1852 114326 -1616
rect 114562 -1852 114646 -1616
rect 114882 -1852 114914 -1616
rect 114294 -1936 114914 -1852
rect 114294 -2172 114326 -1936
rect 114562 -2172 114646 -1936
rect 114882 -2172 114914 -1936
rect 114294 -7964 114914 -2172
rect 118794 264454 119414 298000
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118794 228454 119414 263898
rect 118794 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 119414 228454
rect 118794 228134 119414 228218
rect 118794 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 119414 228134
rect 118794 192454 119414 227898
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 120454 119414 155898
rect 118794 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 119414 120454
rect 118794 120134 119414 120218
rect 118794 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 119414 120134
rect 118794 84454 119414 119898
rect 118794 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 119414 84454
rect 118794 84134 119414 84218
rect 118794 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 119414 84134
rect 118794 48454 119414 83898
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2576 119414 11898
rect 118794 -2812 118826 -2576
rect 119062 -2812 119146 -2576
rect 119382 -2812 119414 -2576
rect 118794 -2896 119414 -2812
rect 118794 -3132 118826 -2896
rect 119062 -3132 119146 -2896
rect 119382 -3132 119414 -2896
rect 118794 -7964 119414 -3132
rect 123294 268954 123914 298000
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 232954 123914 268398
rect 123294 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 123914 232954
rect 123294 232634 123914 232718
rect 123294 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 123914 232634
rect 123294 196954 123914 232398
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 123294 124954 123914 160398
rect 123294 124718 123326 124954
rect 123562 124718 123646 124954
rect 123882 124718 123914 124954
rect 123294 124634 123914 124718
rect 123294 124398 123326 124634
rect 123562 124398 123646 124634
rect 123882 124398 123914 124634
rect 123294 88954 123914 124398
rect 123294 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 123914 88954
rect 123294 88634 123914 88718
rect 123294 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 123914 88634
rect 123294 52954 123914 88398
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3536 123914 16398
rect 123294 -3772 123326 -3536
rect 123562 -3772 123646 -3536
rect 123882 -3772 123914 -3536
rect 123294 -3856 123914 -3772
rect 123294 -4092 123326 -3856
rect 123562 -4092 123646 -3856
rect 123882 -4092 123914 -3856
rect 123294 -7964 123914 -4092
rect 127794 273454 128414 298000
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4496 128414 20898
rect 127794 -4732 127826 -4496
rect 128062 -4732 128146 -4496
rect 128382 -4732 128414 -4496
rect 127794 -4816 128414 -4732
rect 127794 -5052 127826 -4816
rect 128062 -5052 128146 -4816
rect 128382 -5052 128414 -4816
rect 127794 -7964 128414 -5052
rect 132294 277954 132914 298000
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 241954 132914 277398
rect 132294 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 132914 241954
rect 132294 241634 132914 241718
rect 132294 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 132914 241634
rect 132294 205954 132914 241398
rect 132294 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 132914 205954
rect 132294 205634 132914 205718
rect 132294 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 132914 205634
rect 132294 169954 132914 205398
rect 132294 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 132914 169954
rect 132294 169634 132914 169718
rect 132294 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 132914 169634
rect 132294 133954 132914 169398
rect 132294 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 132914 133954
rect 132294 133634 132914 133718
rect 132294 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 132914 133634
rect 132294 97954 132914 133398
rect 132294 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 132914 97954
rect 132294 97634 132914 97718
rect 132294 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 132914 97634
rect 132294 61954 132914 97398
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5456 132914 25398
rect 132294 -5692 132326 -5456
rect 132562 -5692 132646 -5456
rect 132882 -5692 132914 -5456
rect 132294 -5776 132914 -5692
rect 132294 -6012 132326 -5776
rect 132562 -6012 132646 -5776
rect 132882 -6012 132914 -5776
rect 132294 -7964 132914 -6012
rect 136794 282454 137414 298000
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 246454 137414 281898
rect 136794 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 137414 246454
rect 136794 246134 137414 246218
rect 136794 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 137414 246134
rect 136794 210454 137414 245898
rect 136794 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 137414 210454
rect 136794 210134 137414 210218
rect 136794 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 137414 210134
rect 136794 174454 137414 209898
rect 136794 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 137414 174454
rect 136794 174134 137414 174218
rect 136794 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 137414 174134
rect 136794 138454 137414 173898
rect 136794 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 137414 138454
rect 136794 138134 137414 138218
rect 136794 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 137414 138134
rect 136794 102454 137414 137898
rect 136794 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 137414 102454
rect 136794 102134 137414 102218
rect 136794 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 137414 102134
rect 136794 66454 137414 101898
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6416 137414 29898
rect 136794 -6652 136826 -6416
rect 137062 -6652 137146 -6416
rect 137382 -6652 137414 -6416
rect 136794 -6736 137414 -6652
rect 136794 -6972 136826 -6736
rect 137062 -6972 137146 -6736
rect 137382 -6972 137414 -6736
rect 136794 -7964 137414 -6972
rect 141294 286954 141914 298000
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 214954 141914 250398
rect 141294 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 141914 214954
rect 141294 214634 141914 214718
rect 141294 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 141914 214634
rect 141294 178954 141914 214398
rect 141294 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 141914 178954
rect 141294 178634 141914 178718
rect 141294 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 141914 178634
rect 141294 142954 141914 178398
rect 141294 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 141914 142954
rect 141294 142634 141914 142718
rect 141294 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 141914 142634
rect 141294 106954 141914 142398
rect 141294 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 141914 106954
rect 141294 106634 141914 106718
rect 141294 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 141914 106634
rect 141294 70954 141914 106398
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7376 141914 34398
rect 141294 -7612 141326 -7376
rect 141562 -7612 141646 -7376
rect 141882 -7612 141914 -7376
rect 141294 -7696 141914 -7612
rect 141294 -7932 141326 -7696
rect 141562 -7932 141646 -7696
rect 141882 -7932 141914 -7696
rect 141294 -7964 141914 -7932
rect 145794 291454 146414 298000
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -656 146414 2898
rect 145794 -892 145826 -656
rect 146062 -892 146146 -656
rect 146382 -892 146414 -656
rect 145794 -976 146414 -892
rect 145794 -1212 145826 -976
rect 146062 -1212 146146 -976
rect 146382 -1212 146414 -976
rect 145794 -7964 146414 -1212
rect 150294 295954 150914 298000
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 223954 150914 259398
rect 150294 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 150914 223954
rect 150294 223634 150914 223718
rect 150294 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 150914 223634
rect 150294 187954 150914 223398
rect 150294 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 150914 187954
rect 150294 187634 150914 187718
rect 150294 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 150914 187634
rect 150294 151954 150914 187398
rect 150294 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 150914 151954
rect 150294 151634 150914 151718
rect 150294 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 150914 151634
rect 150294 115954 150914 151398
rect 150294 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 150914 115954
rect 150294 115634 150914 115718
rect 150294 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 150914 115634
rect 150294 79954 150914 115398
rect 150294 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 150914 79954
rect 150294 79634 150914 79718
rect 150294 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 150914 79634
rect 150294 43954 150914 79398
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1616 150914 7398
rect 150294 -1852 150326 -1616
rect 150562 -1852 150646 -1616
rect 150882 -1852 150914 -1616
rect 150294 -1936 150914 -1852
rect 150294 -2172 150326 -1936
rect 150562 -2172 150646 -1936
rect 150882 -2172 150914 -1936
rect 150294 -7964 150914 -2172
rect 154794 264454 155414 298000
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 228454 155414 263898
rect 154794 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 155414 228454
rect 154794 228134 155414 228218
rect 154794 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 155414 228134
rect 154794 192454 155414 227898
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 154794 156454 155414 191898
rect 154794 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 155414 156454
rect 154794 156134 155414 156218
rect 154794 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 155414 156134
rect 154794 120454 155414 155898
rect 154794 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 155414 120454
rect 154794 120134 155414 120218
rect 154794 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 155414 120134
rect 154794 84454 155414 119898
rect 154794 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 155414 84454
rect 154794 84134 155414 84218
rect 154794 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 155414 84134
rect 154794 48454 155414 83898
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2576 155414 11898
rect 154794 -2812 154826 -2576
rect 155062 -2812 155146 -2576
rect 155382 -2812 155414 -2576
rect 154794 -2896 155414 -2812
rect 154794 -3132 154826 -2896
rect 155062 -3132 155146 -2896
rect 155382 -3132 155414 -2896
rect 154794 -7964 155414 -3132
rect 159294 268954 159914 298000
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 232954 159914 268398
rect 159294 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 159914 232954
rect 159294 232634 159914 232718
rect 159294 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 159914 232634
rect 159294 196954 159914 232398
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 159294 160954 159914 196398
rect 159294 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 159914 160954
rect 159294 160634 159914 160718
rect 159294 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 159914 160634
rect 159294 124954 159914 160398
rect 159294 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 159914 124954
rect 159294 124634 159914 124718
rect 159294 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 159914 124634
rect 159294 88954 159914 124398
rect 159294 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 159914 88954
rect 159294 88634 159914 88718
rect 159294 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 159914 88634
rect 159294 52954 159914 88398
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3536 159914 16398
rect 159294 -3772 159326 -3536
rect 159562 -3772 159646 -3536
rect 159882 -3772 159914 -3536
rect 159294 -3856 159914 -3772
rect 159294 -4092 159326 -3856
rect 159562 -4092 159646 -3856
rect 159882 -4092 159914 -3856
rect 159294 -7964 159914 -4092
rect 163794 273454 164414 298000
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4496 164414 20898
rect 163794 -4732 163826 -4496
rect 164062 -4732 164146 -4496
rect 164382 -4732 164414 -4496
rect 163794 -4816 164414 -4732
rect 163794 -5052 163826 -4816
rect 164062 -5052 164146 -4816
rect 164382 -5052 164414 -4816
rect 163794 -7964 164414 -5052
rect 168294 277954 168914 298000
rect 169158 297941 169218 301139
rect 169155 297940 169221 297941
rect 169155 297876 169156 297940
rect 169220 297876 169221 297940
rect 169155 297875 169221 297876
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 241954 168914 277398
rect 168294 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 168914 241954
rect 168294 241634 168914 241718
rect 168294 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 168914 241634
rect 168294 205954 168914 241398
rect 168294 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 168914 205954
rect 168294 205634 168914 205718
rect 168294 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 168914 205634
rect 168294 169954 168914 205398
rect 168294 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 168914 169954
rect 168294 169634 168914 169718
rect 168294 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 168914 169634
rect 168294 133954 168914 169398
rect 168294 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 168914 133954
rect 168294 133634 168914 133718
rect 168294 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 168914 133634
rect 168294 97954 168914 133398
rect 168294 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 168914 97954
rect 168294 97634 168914 97718
rect 168294 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 168914 97634
rect 168294 61954 168914 97398
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5456 168914 25398
rect 168294 -5692 168326 -5456
rect 168562 -5692 168646 -5456
rect 168882 -5692 168914 -5456
rect 168294 -5776 168914 -5692
rect 168294 -6012 168326 -5776
rect 168562 -6012 168646 -5776
rect 168882 -6012 168914 -5776
rect 168294 -7964 168914 -6012
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 246454 173414 281898
rect 172794 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 173414 246454
rect 172794 246134 173414 246218
rect 172794 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 173414 246134
rect 172794 210454 173414 245898
rect 172794 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 173414 210454
rect 172794 210134 173414 210218
rect 172794 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 173414 210134
rect 172794 174454 173414 209898
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 172794 138454 173414 173898
rect 172794 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 173414 138454
rect 172794 138134 173414 138218
rect 172794 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 173414 138134
rect 172794 102454 173414 137898
rect 172794 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 173414 102454
rect 172794 102134 173414 102218
rect 172794 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 173414 102134
rect 172794 66454 173414 101898
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6416 173414 29898
rect 172794 -6652 172826 -6416
rect 173062 -6652 173146 -6416
rect 173382 -6652 173414 -6416
rect 172794 -6736 173414 -6652
rect 172794 -6972 172826 -6736
rect 173062 -6972 173146 -6736
rect 173382 -6972 173414 -6736
rect 172794 -7964 173414 -6972
rect 177294 711868 177914 711900
rect 177294 711632 177326 711868
rect 177562 711632 177646 711868
rect 177882 711632 177914 711868
rect 177294 711548 177914 711632
rect 177294 711312 177326 711548
rect 177562 711312 177646 711548
rect 177882 711312 177914 711548
rect 177294 682954 177914 711312
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 214954 177914 250398
rect 177294 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 177914 214954
rect 177294 214634 177914 214718
rect 177294 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 177914 214634
rect 177294 178954 177914 214398
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 106954 177914 142398
rect 177294 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 177914 106954
rect 177294 106634 177914 106718
rect 177294 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 177914 106634
rect 177294 70954 177914 106398
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7376 177914 34398
rect 177294 -7612 177326 -7376
rect 177562 -7612 177646 -7376
rect 177882 -7612 177914 -7376
rect 177294 -7696 177914 -7612
rect 177294 -7932 177326 -7696
rect 177562 -7932 177646 -7696
rect 177882 -7932 177914 -7696
rect 177294 -7964 177914 -7932
rect 181794 705148 182414 711900
rect 181794 704912 181826 705148
rect 182062 704912 182146 705148
rect 182382 704912 182414 705148
rect 181794 704828 182414 704912
rect 181794 704592 181826 704828
rect 182062 704592 182146 704828
rect 182382 704592 182414 704828
rect 181794 687454 182414 704592
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -656 182414 2898
rect 181794 -892 181826 -656
rect 182062 -892 182146 -656
rect 182382 -892 182414 -656
rect 181794 -976 182414 -892
rect 181794 -1212 181826 -976
rect 182062 -1212 182146 -976
rect 182382 -1212 182414 -976
rect 181794 -7964 182414 -1212
rect 186294 706108 186914 711900
rect 186294 705872 186326 706108
rect 186562 705872 186646 706108
rect 186882 705872 186914 706108
rect 186294 705788 186914 705872
rect 186294 705552 186326 705788
rect 186562 705552 186646 705788
rect 186882 705552 186914 705788
rect 186294 691954 186914 705552
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 259954 186914 295398
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 223954 186914 259398
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 187954 186914 223398
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 115954 186914 151398
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 186294 79954 186914 115398
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 186294 79634 186914 79718
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1616 186914 7398
rect 186294 -1852 186326 -1616
rect 186562 -1852 186646 -1616
rect 186882 -1852 186914 -1616
rect 186294 -1936 186914 -1852
rect 186294 -2172 186326 -1936
rect 186562 -2172 186646 -1936
rect 186882 -2172 186914 -1936
rect 186294 -7964 186914 -2172
rect 190794 707068 191414 711900
rect 190794 706832 190826 707068
rect 191062 706832 191146 707068
rect 191382 706832 191414 707068
rect 190794 706748 191414 706832
rect 190794 706512 190826 706748
rect 191062 706512 191146 706748
rect 191382 706512 191414 706748
rect 190794 696454 191414 706512
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 228454 191414 263898
rect 190794 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 191414 228454
rect 190794 228134 191414 228218
rect 190794 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 191414 228134
rect 190794 192454 191414 227898
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 120454 191414 155898
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 84454 191414 119898
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2576 191414 11898
rect 190794 -2812 190826 -2576
rect 191062 -2812 191146 -2576
rect 191382 -2812 191414 -2576
rect 190794 -2896 191414 -2812
rect 190794 -3132 190826 -2896
rect 191062 -3132 191146 -2896
rect 191382 -3132 191414 -2896
rect 190794 -7964 191414 -3132
rect 195294 708028 195914 711900
rect 195294 707792 195326 708028
rect 195562 707792 195646 708028
rect 195882 707792 195914 708028
rect 195294 707708 195914 707792
rect 195294 707472 195326 707708
rect 195562 707472 195646 707708
rect 195882 707472 195914 707708
rect 195294 700954 195914 707472
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 195294 232954 195914 268398
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 196954 195914 232398
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3536 195914 16398
rect 195294 -3772 195326 -3536
rect 195562 -3772 195646 -3536
rect 195882 -3772 195914 -3536
rect 195294 -3856 195914 -3772
rect 195294 -4092 195326 -3856
rect 195562 -4092 195646 -3856
rect 195882 -4092 195914 -3856
rect 195294 -7964 195914 -4092
rect 199794 708988 200414 711900
rect 199794 708752 199826 708988
rect 200062 708752 200146 708988
rect 200382 708752 200414 708988
rect 199794 708668 200414 708752
rect 199794 708432 199826 708668
rect 200062 708432 200146 708668
rect 200382 708432 200414 708668
rect 199794 669454 200414 708432
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4496 200414 20898
rect 199794 -4732 199826 -4496
rect 200062 -4732 200146 -4496
rect 200382 -4732 200414 -4496
rect 199794 -4816 200414 -4732
rect 199794 -5052 199826 -4816
rect 200062 -5052 200146 -4816
rect 200382 -5052 200414 -4816
rect 199794 -7964 200414 -5052
rect 204294 709948 204914 711900
rect 204294 709712 204326 709948
rect 204562 709712 204646 709948
rect 204882 709712 204914 709948
rect 204294 709628 204914 709712
rect 204294 709392 204326 709628
rect 204562 709392 204646 709628
rect 204882 709392 204914 709628
rect 204294 673954 204914 709392
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 241954 204914 277398
rect 204294 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 204914 241954
rect 204294 241634 204914 241718
rect 204294 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 204914 241634
rect 204294 205954 204914 241398
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5456 204914 25398
rect 204294 -5692 204326 -5456
rect 204562 -5692 204646 -5456
rect 204882 -5692 204914 -5456
rect 204294 -5776 204914 -5692
rect 204294 -6012 204326 -5776
rect 204562 -6012 204646 -5776
rect 204882 -6012 204914 -5776
rect 204294 -7964 204914 -6012
rect 208794 710908 209414 711900
rect 208794 710672 208826 710908
rect 209062 710672 209146 710908
rect 209382 710672 209414 710908
rect 208794 710588 209414 710672
rect 208794 710352 208826 710588
rect 209062 710352 209146 710588
rect 209382 710352 209414 710588
rect 208794 678454 209414 710352
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 213294 711868 213914 711900
rect 213294 711632 213326 711868
rect 213562 711632 213646 711868
rect 213882 711632 213914 711868
rect 213294 711548 213914 711632
rect 213294 711312 213326 711548
rect 213562 711312 213646 711548
rect 213882 711312 213914 711548
rect 213294 682954 213914 711312
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 217794 705148 218414 711900
rect 217794 704912 217826 705148
rect 218062 704912 218146 705148
rect 218382 704912 218414 705148
rect 217794 704828 218414 704912
rect 217794 704592 217826 704828
rect 218062 704592 218146 704828
rect 218382 704592 218414 704828
rect 217794 687454 218414 704592
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 565308 218414 578898
rect 222294 706108 222914 711900
rect 222294 705872 222326 706108
rect 222562 705872 222646 706108
rect 222882 705872 222914 706108
rect 222294 705788 222914 705872
rect 222294 705552 222326 705788
rect 222562 705552 222646 705788
rect 222882 705552 222914 705788
rect 222294 691954 222914 705552
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 565308 222914 583398
rect 226794 707068 227414 711900
rect 226794 706832 226826 707068
rect 227062 706832 227146 707068
rect 227382 706832 227414 707068
rect 226794 706748 227414 706832
rect 226794 706512 226826 706748
rect 227062 706512 227146 706748
rect 227382 706512 227414 706748
rect 226794 696454 227414 706512
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 565308 227414 587898
rect 231294 708028 231914 711900
rect 231294 707792 231326 708028
rect 231562 707792 231646 708028
rect 231882 707792 231914 708028
rect 231294 707708 231914 707792
rect 231294 707472 231326 707708
rect 231562 707472 231646 707708
rect 231882 707472 231914 707708
rect 231294 700954 231914 707472
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 565308 231914 592398
rect 235794 708988 236414 711900
rect 235794 708752 235826 708988
rect 236062 708752 236146 708988
rect 236382 708752 236414 708988
rect 235794 708668 236414 708752
rect 235794 708432 235826 708668
rect 236062 708432 236146 708668
rect 236382 708432 236414 708668
rect 235794 669454 236414 708432
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 565308 236414 596898
rect 240294 709948 240914 711900
rect 240294 709712 240326 709948
rect 240562 709712 240646 709948
rect 240882 709712 240914 709948
rect 240294 709628 240914 709712
rect 240294 709392 240326 709628
rect 240562 709392 240646 709628
rect 240882 709392 240914 709628
rect 240294 673954 240914 709392
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 565308 240914 565398
rect 244794 710908 245414 711900
rect 244794 710672 244826 710908
rect 245062 710672 245146 710908
rect 245382 710672 245414 710908
rect 244794 710588 245414 710672
rect 244794 710352 244826 710588
rect 245062 710352 245146 710588
rect 245382 710352 245414 710588
rect 244794 678454 245414 710352
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 565308 245414 569898
rect 249294 711868 249914 711900
rect 249294 711632 249326 711868
rect 249562 711632 249646 711868
rect 249882 711632 249914 711868
rect 249294 711548 249914 711632
rect 249294 711312 249326 711548
rect 249562 711312 249646 711548
rect 249882 711312 249914 711548
rect 249294 682954 249914 711312
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 565308 249914 574398
rect 253794 705148 254414 711900
rect 253794 704912 253826 705148
rect 254062 704912 254146 705148
rect 254382 704912 254414 705148
rect 253794 704828 254414 704912
rect 253794 704592 253826 704828
rect 254062 704592 254146 704828
rect 254382 704592 254414 704828
rect 253794 687454 254414 704592
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 565308 254414 578898
rect 258294 706108 258914 711900
rect 258294 705872 258326 706108
rect 258562 705872 258646 706108
rect 258882 705872 258914 706108
rect 258294 705788 258914 705872
rect 258294 705552 258326 705788
rect 258562 705552 258646 705788
rect 258882 705552 258914 705788
rect 258294 691954 258914 705552
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 565308 258914 583398
rect 262794 707068 263414 711900
rect 262794 706832 262826 707068
rect 263062 706832 263146 707068
rect 263382 706832 263414 707068
rect 262794 706748 263414 706832
rect 262794 706512 262826 706748
rect 263062 706512 263146 706748
rect 263382 706512 263414 706748
rect 262794 696454 263414 706512
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 565308 263414 587898
rect 267294 708028 267914 711900
rect 267294 707792 267326 708028
rect 267562 707792 267646 708028
rect 267882 707792 267914 708028
rect 267294 707708 267914 707792
rect 267294 707472 267326 707708
rect 267562 707472 267646 707708
rect 267882 707472 267914 707708
rect 267294 700954 267914 707472
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 565308 267914 592398
rect 271794 708988 272414 711900
rect 271794 708752 271826 708988
rect 272062 708752 272146 708988
rect 272382 708752 272414 708988
rect 271794 708668 272414 708752
rect 271794 708432 271826 708668
rect 272062 708432 272146 708668
rect 272382 708432 272414 708668
rect 271794 669454 272414 708432
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 565308 272414 596898
rect 276294 709948 276914 711900
rect 276294 709712 276326 709948
rect 276562 709712 276646 709948
rect 276882 709712 276914 709948
rect 276294 709628 276914 709712
rect 276294 709392 276326 709628
rect 276562 709392 276646 709628
rect 276882 709392 276914 709628
rect 276294 673954 276914 709392
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 565308 276914 565398
rect 280794 710908 281414 711900
rect 280794 710672 280826 710908
rect 281062 710672 281146 710908
rect 281382 710672 281414 710908
rect 280794 710588 281414 710672
rect 280794 710352 280826 710588
rect 281062 710352 281146 710588
rect 281382 710352 281414 710588
rect 280794 678454 281414 710352
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 565308 281414 569898
rect 285294 711868 285914 711900
rect 285294 711632 285326 711868
rect 285562 711632 285646 711868
rect 285882 711632 285914 711868
rect 285294 711548 285914 711632
rect 285294 711312 285326 711548
rect 285562 711312 285646 711548
rect 285882 711312 285914 711548
rect 285294 682954 285914 711312
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 565308 285914 574398
rect 289794 705148 290414 711900
rect 289794 704912 289826 705148
rect 290062 704912 290146 705148
rect 290382 704912 290414 705148
rect 289794 704828 290414 704912
rect 289794 704592 289826 704828
rect 290062 704592 290146 704828
rect 290382 704592 290414 704828
rect 289794 687454 290414 704592
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 565308 290414 578898
rect 294294 706108 294914 711900
rect 294294 705872 294326 706108
rect 294562 705872 294646 706108
rect 294882 705872 294914 706108
rect 294294 705788 294914 705872
rect 294294 705552 294326 705788
rect 294562 705552 294646 705788
rect 294882 705552 294914 705788
rect 294294 691954 294914 705552
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 565308 294914 583398
rect 298794 707068 299414 711900
rect 298794 706832 298826 707068
rect 299062 706832 299146 707068
rect 299382 706832 299414 707068
rect 298794 706748 299414 706832
rect 298794 706512 298826 706748
rect 299062 706512 299146 706748
rect 299382 706512 299414 706748
rect 298794 696454 299414 706512
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 565308 299414 587898
rect 303294 708028 303914 711900
rect 303294 707792 303326 708028
rect 303562 707792 303646 708028
rect 303882 707792 303914 708028
rect 303294 707708 303914 707792
rect 303294 707472 303326 707708
rect 303562 707472 303646 707708
rect 303882 707472 303914 707708
rect 303294 700954 303914 707472
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 565308 303914 592398
rect 307794 708988 308414 711900
rect 307794 708752 307826 708988
rect 308062 708752 308146 708988
rect 308382 708752 308414 708988
rect 307794 708668 308414 708752
rect 307794 708432 307826 708668
rect 308062 708432 308146 708668
rect 308382 708432 308414 708668
rect 307794 669454 308414 708432
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 565308 308414 596898
rect 312294 709948 312914 711900
rect 312294 709712 312326 709948
rect 312562 709712 312646 709948
rect 312882 709712 312914 709948
rect 312294 709628 312914 709712
rect 312294 709392 312326 709628
rect 312562 709392 312646 709628
rect 312882 709392 312914 709628
rect 312294 673954 312914 709392
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 565308 312914 565398
rect 316794 710908 317414 711900
rect 316794 710672 316826 710908
rect 317062 710672 317146 710908
rect 317382 710672 317414 710908
rect 316794 710588 317414 710672
rect 316794 710352 316826 710588
rect 317062 710352 317146 710588
rect 317382 710352 317414 710588
rect 316794 678454 317414 710352
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 565308 317414 569898
rect 321294 711868 321914 711900
rect 321294 711632 321326 711868
rect 321562 711632 321646 711868
rect 321882 711632 321914 711868
rect 321294 711548 321914 711632
rect 321294 711312 321326 711548
rect 321562 711312 321646 711548
rect 321882 711312 321914 711548
rect 321294 682954 321914 711312
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 565308 321914 574398
rect 325794 705148 326414 711900
rect 325794 704912 325826 705148
rect 326062 704912 326146 705148
rect 326382 704912 326414 705148
rect 325794 704828 326414 704912
rect 325794 704592 325826 704828
rect 326062 704592 326146 704828
rect 326382 704592 326414 704828
rect 325794 687454 326414 704592
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 565308 326414 578898
rect 330294 706108 330914 711900
rect 330294 705872 330326 706108
rect 330562 705872 330646 706108
rect 330882 705872 330914 706108
rect 330294 705788 330914 705872
rect 330294 705552 330326 705788
rect 330562 705552 330646 705788
rect 330882 705552 330914 705788
rect 330294 691954 330914 705552
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 565308 330914 583398
rect 334794 707068 335414 711900
rect 334794 706832 334826 707068
rect 335062 706832 335146 707068
rect 335382 706832 335414 707068
rect 334794 706748 335414 706832
rect 334794 706512 334826 706748
rect 335062 706512 335146 706748
rect 335382 706512 335414 706748
rect 334794 696454 335414 706512
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 565308 335414 587898
rect 339294 708028 339914 711900
rect 339294 707792 339326 708028
rect 339562 707792 339646 708028
rect 339882 707792 339914 708028
rect 339294 707708 339914 707792
rect 339294 707472 339326 707708
rect 339562 707472 339646 707708
rect 339882 707472 339914 707708
rect 339294 700954 339914 707472
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 565308 339914 592398
rect 343794 708988 344414 711900
rect 343794 708752 343826 708988
rect 344062 708752 344146 708988
rect 344382 708752 344414 708988
rect 343794 708668 344414 708752
rect 343794 708432 343826 708668
rect 344062 708432 344146 708668
rect 344382 708432 344414 708668
rect 343794 669454 344414 708432
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 565308 344414 596898
rect 348294 709948 348914 711900
rect 348294 709712 348326 709948
rect 348562 709712 348646 709948
rect 348882 709712 348914 709948
rect 348294 709628 348914 709712
rect 348294 709392 348326 709628
rect 348562 709392 348646 709628
rect 348882 709392 348914 709628
rect 348294 673954 348914 709392
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 565308 348914 565398
rect 352794 710908 353414 711900
rect 352794 710672 352826 710908
rect 353062 710672 353146 710908
rect 353382 710672 353414 710908
rect 352794 710588 353414 710672
rect 352794 710352 352826 710588
rect 353062 710352 353146 710588
rect 353382 710352 353414 710588
rect 352794 678454 353414 710352
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 565308 353414 569898
rect 357294 711868 357914 711900
rect 357294 711632 357326 711868
rect 357562 711632 357646 711868
rect 357882 711632 357914 711868
rect 357294 711548 357914 711632
rect 357294 711312 357326 711548
rect 357562 711312 357646 711548
rect 357882 711312 357914 711548
rect 357294 682954 357914 711312
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 565308 357914 574398
rect 361794 705148 362414 711900
rect 361794 704912 361826 705148
rect 362062 704912 362146 705148
rect 362382 704912 362414 705148
rect 361794 704828 362414 704912
rect 361794 704592 361826 704828
rect 362062 704592 362146 704828
rect 362382 704592 362414 704828
rect 361794 687454 362414 704592
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 220272 547954 220620 547986
rect 220272 547718 220328 547954
rect 220564 547718 220620 547954
rect 220272 547634 220620 547718
rect 220272 547398 220328 547634
rect 220564 547398 220620 547634
rect 220272 547366 220620 547398
rect 356000 547954 356348 547986
rect 356000 547718 356056 547954
rect 356292 547718 356348 547954
rect 356000 547634 356348 547718
rect 356000 547398 356056 547634
rect 356292 547398 356348 547634
rect 356000 547366 356348 547398
rect 220952 543454 221300 543486
rect 220952 543218 221008 543454
rect 221244 543218 221300 543454
rect 220952 543134 221300 543218
rect 220952 542898 221008 543134
rect 221244 542898 221300 543134
rect 220952 542866 221300 542898
rect 355320 543454 355668 543486
rect 355320 543218 355376 543454
rect 355612 543218 355668 543454
rect 355320 543134 355668 543218
rect 355320 542898 355376 543134
rect 355612 542898 355668 543134
rect 355320 542866 355668 542898
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 220272 511954 220620 511986
rect 220272 511718 220328 511954
rect 220564 511718 220620 511954
rect 220272 511634 220620 511718
rect 220272 511398 220328 511634
rect 220564 511398 220620 511634
rect 220272 511366 220620 511398
rect 356000 511954 356348 511986
rect 356000 511718 356056 511954
rect 356292 511718 356348 511954
rect 356000 511634 356348 511718
rect 356000 511398 356056 511634
rect 356292 511398 356348 511634
rect 356000 511366 356348 511398
rect 220952 507454 221300 507486
rect 220952 507218 221008 507454
rect 221244 507218 221300 507454
rect 220952 507134 221300 507218
rect 220952 506898 221008 507134
rect 221244 506898 221300 507134
rect 220952 506866 221300 506898
rect 355320 507454 355668 507486
rect 355320 507218 355376 507454
rect 355612 507218 355668 507454
rect 355320 507134 355668 507218
rect 355320 506898 355376 507134
rect 355612 506898 355668 507134
rect 355320 506866 355668 506898
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 236056 479770 236116 480080
rect 237144 479770 237204 480080
rect 238232 479770 238292 480080
rect 239592 479770 239652 480080
rect 240544 479770 240604 480080
rect 241768 479770 241828 480080
rect 243128 479770 243188 480080
rect 236056 479710 236194 479770
rect 237144 479710 237298 479770
rect 238232 479710 238402 479770
rect 239592 479710 239690 479770
rect 240544 479710 240610 479770
rect 241768 479710 241898 479770
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 211659 435028 211725 435029
rect 211659 434964 211660 435028
rect 211724 434964 211725 435028
rect 211659 434963 211725 434964
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 246454 209414 281898
rect 208794 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 209414 246454
rect 208794 246134 209414 246218
rect 208794 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 209414 246134
rect 208794 210454 209414 245898
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 211662 110533 211722 434963
rect 213294 430954 213914 466398
rect 217794 471454 218414 478000
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 214419 435300 214485 435301
rect 214419 435236 214420 435300
rect 214484 435236 214485 435300
rect 214419 435235 214485 435236
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 212395 265572 212461 265573
rect 212395 265508 212396 265572
rect 212460 265508 212461 265572
rect 212395 265507 212461 265508
rect 211659 110532 211725 110533
rect 211659 110468 211660 110532
rect 211724 110468 211725 110532
rect 211659 110467 211725 110468
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6416 209414 29898
rect 212398 3501 212458 265507
rect 213131 262852 213197 262853
rect 213131 262788 213132 262852
rect 213196 262788 213197 262852
rect 213131 262787 213197 262788
rect 213134 3501 213194 262787
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 214954 213914 250398
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 214422 162893 214482 435235
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 215891 435164 215957 435165
rect 215891 435100 215892 435164
rect 215956 435100 215957 435164
rect 215891 435099 215957 435100
rect 217794 435134 218414 435218
rect 214787 303244 214853 303245
rect 214787 303180 214788 303244
rect 214852 303180 214853 303244
rect 214787 303179 214853 303180
rect 214419 162892 214485 162893
rect 214419 162828 214420 162892
rect 214484 162828 214485 162892
rect 214419 162827 214485 162828
rect 214790 157861 214850 303179
rect 215155 302972 215221 302973
rect 215155 302908 215156 302972
rect 215220 302908 215221 302972
rect 215155 302907 215221 302908
rect 214971 301748 215037 301749
rect 214971 301684 214972 301748
rect 215036 301684 215037 301748
rect 214971 301683 215037 301684
rect 214787 157860 214853 157861
rect 214787 157796 214788 157860
rect 214852 157796 214853 157860
rect 214787 157795 214853 157796
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 212395 3500 212461 3501
rect 212395 3436 212396 3500
rect 212460 3436 212461 3500
rect 212395 3435 212461 3436
rect 213131 3500 213197 3501
rect 213131 3436 213132 3500
rect 213196 3436 213197 3500
rect 213131 3435 213197 3436
rect 208794 -6652 208826 -6416
rect 209062 -6652 209146 -6416
rect 209382 -6652 209414 -6416
rect 208794 -6736 209414 -6652
rect 208794 -6972 208826 -6736
rect 209062 -6972 209146 -6736
rect 209382 -6972 209414 -6736
rect 208794 -7964 209414 -6972
rect 213294 -7376 213914 34398
rect 214974 3501 215034 301683
rect 215158 3909 215218 302907
rect 215894 31789 215954 435099
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217547 305964 217613 305965
rect 217547 305900 217548 305964
rect 217612 305900 217613 305964
rect 217547 305899 217613 305900
rect 217363 305828 217429 305829
rect 217363 305764 217364 305828
rect 217428 305764 217429 305828
rect 217363 305763 217429 305764
rect 216443 303380 216509 303381
rect 216443 303316 216444 303380
rect 216508 303316 216509 303380
rect 216443 303315 216509 303316
rect 216075 303108 216141 303109
rect 216075 303044 216076 303108
rect 216140 303044 216141 303108
rect 216075 303043 216141 303044
rect 216078 158405 216138 303043
rect 216259 284884 216325 284885
rect 216259 284820 216260 284884
rect 216324 284820 216325 284884
rect 216259 284819 216325 284820
rect 216075 158404 216141 158405
rect 216075 158340 216076 158404
rect 216140 158340 216141 158404
rect 216075 158339 216141 158340
rect 215891 31788 215957 31789
rect 215891 31724 215892 31788
rect 215956 31724 215957 31788
rect 215891 31723 215957 31724
rect 215155 3908 215221 3909
rect 215155 3844 215156 3908
rect 215220 3844 215221 3908
rect 215155 3843 215221 3844
rect 216262 3501 216322 284819
rect 216446 3773 216506 303315
rect 216995 302836 217061 302837
rect 216995 302772 216996 302836
rect 217060 302772 217061 302836
rect 216995 302771 217061 302772
rect 216998 157997 217058 302771
rect 217179 301476 217245 301477
rect 217179 301412 217180 301476
rect 217244 301412 217245 301476
rect 217179 301411 217245 301412
rect 216995 157996 217061 157997
rect 216995 157932 216996 157996
rect 217060 157932 217061 157996
rect 216995 157931 217061 157932
rect 217182 155277 217242 301411
rect 217366 158269 217426 305763
rect 217363 158268 217429 158269
rect 217363 158204 217364 158268
rect 217428 158204 217429 158268
rect 217363 158203 217429 158204
rect 217550 158133 217610 305899
rect 217794 291454 218414 326898
rect 222294 475954 222914 478000
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 219019 306236 219085 306237
rect 219019 306172 219020 306236
rect 219084 306172 219085 306236
rect 219019 306171 219085 306172
rect 218835 306100 218901 306101
rect 218835 306036 218836 306100
rect 218900 306036 218901 306100
rect 218835 306035 218901 306036
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 245308 218414 254898
rect 218651 243540 218717 243541
rect 218651 243476 218652 243540
rect 218716 243476 218717 243540
rect 218651 243475 218717 243476
rect 217547 158132 217613 158133
rect 217547 158068 217548 158132
rect 217612 158068 217613 158132
rect 217547 158067 217613 158068
rect 217179 155276 217245 155277
rect 217179 155212 217180 155276
rect 217244 155212 217245 155276
rect 217179 155211 217245 155212
rect 217794 147454 218414 158000
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 216443 3772 216509 3773
rect 216443 3708 216444 3772
rect 216508 3708 216509 3772
rect 216443 3707 216509 3708
rect 214971 3500 215037 3501
rect 214971 3436 214972 3500
rect 215036 3436 215037 3500
rect 214971 3435 215037 3436
rect 216259 3500 216325 3501
rect 216259 3436 216260 3500
rect 216324 3436 216325 3500
rect 216259 3435 216325 3436
rect 217794 3454 218414 38898
rect 218654 3501 218714 243475
rect 218838 158677 218898 306035
rect 218835 158676 218901 158677
rect 218835 158612 218836 158676
rect 218900 158612 218901 158676
rect 218835 158611 218901 158612
rect 219022 158541 219082 306171
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 219203 293180 219269 293181
rect 219203 293116 219204 293180
rect 219268 293116 219269 293180
rect 219203 293115 219269 293116
rect 219019 158540 219085 158541
rect 219019 158476 219020 158540
rect 219084 158476 219085 158540
rect 219019 158475 219085 158476
rect 219206 3637 219266 293115
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 245308 222914 259398
rect 226794 444454 227414 478000
rect 236134 476373 236194 479710
rect 236131 476372 236197 476373
rect 236131 476308 236132 476372
rect 236196 476308 236197 476372
rect 236131 476307 236197 476308
rect 237238 476237 237298 479710
rect 238342 477325 238402 479710
rect 238339 477324 238405 477325
rect 238339 477260 238340 477324
rect 238404 477260 238405 477324
rect 238339 477259 238405 477260
rect 239630 476917 239690 479710
rect 240550 476917 240610 479710
rect 241838 477189 241898 479710
rect 243126 479710 243188 479770
rect 244216 479770 244276 480080
rect 245440 479770 245500 480080
rect 246528 479770 246588 480080
rect 247616 479770 247676 480080
rect 248296 479770 248356 480080
rect 248704 479770 248764 480080
rect 244216 479710 244290 479770
rect 245440 479710 245578 479770
rect 246528 479710 246682 479770
rect 247616 479710 247786 479770
rect 241835 477188 241901 477189
rect 241835 477124 241836 477188
rect 241900 477124 241901 477188
rect 241835 477123 241901 477124
rect 239627 476916 239693 476917
rect 239627 476852 239628 476916
rect 239692 476852 239693 476916
rect 239627 476851 239693 476852
rect 240547 476916 240613 476917
rect 240547 476852 240548 476916
rect 240612 476852 240613 476916
rect 240547 476851 240613 476852
rect 243126 476237 243186 479710
rect 244230 476373 244290 479710
rect 244227 476372 244293 476373
rect 244227 476308 244228 476372
rect 244292 476308 244293 476372
rect 244227 476307 244293 476308
rect 245518 476237 245578 479710
rect 246622 476373 246682 479710
rect 246619 476372 246685 476373
rect 246619 476308 246620 476372
rect 246684 476308 246685 476372
rect 246619 476307 246685 476308
rect 247726 476237 247786 479710
rect 248278 479710 248356 479770
rect 248646 479710 248764 479770
rect 250064 479770 250124 480080
rect 250744 479770 250804 480080
rect 251288 479770 251348 480080
rect 252376 479770 252436 480080
rect 253464 479770 253524 480080
rect 250064 479710 250178 479770
rect 250744 479710 250914 479770
rect 251288 479710 251466 479770
rect 248278 476645 248338 479710
rect 248275 476644 248341 476645
rect 248275 476580 248276 476644
rect 248340 476580 248341 476644
rect 248275 476579 248341 476580
rect 248646 476237 248706 479710
rect 250118 476373 250178 479710
rect 250115 476372 250181 476373
rect 250115 476308 250116 476372
rect 250180 476308 250181 476372
rect 250115 476307 250181 476308
rect 250854 476237 250914 479710
rect 251406 476373 251466 479710
rect 252326 479710 252436 479770
rect 253430 479710 253524 479770
rect 253600 479770 253660 480080
rect 254552 479770 254612 480080
rect 255912 479770 255972 480080
rect 253600 479710 253674 479770
rect 251403 476372 251469 476373
rect 251403 476308 251404 476372
rect 251468 476308 251469 476372
rect 251403 476307 251469 476308
rect 252326 476237 252386 479710
rect 253430 476237 253490 479710
rect 253614 476509 253674 479710
rect 254534 479710 254612 479770
rect 255822 479710 255972 479770
rect 256048 479770 256108 480080
rect 257000 479770 257060 480080
rect 258088 479770 258148 480080
rect 256048 479710 256250 479770
rect 257000 479710 257170 479770
rect 253611 476508 253677 476509
rect 253611 476444 253612 476508
rect 253676 476444 253677 476508
rect 253611 476443 253677 476444
rect 237235 476236 237301 476237
rect 237235 476172 237236 476236
rect 237300 476172 237301 476236
rect 237235 476171 237301 476172
rect 243123 476236 243189 476237
rect 243123 476172 243124 476236
rect 243188 476172 243189 476236
rect 243123 476171 243189 476172
rect 245515 476236 245581 476237
rect 245515 476172 245516 476236
rect 245580 476172 245581 476236
rect 245515 476171 245581 476172
rect 247723 476236 247789 476237
rect 247723 476172 247724 476236
rect 247788 476172 247789 476236
rect 247723 476171 247789 476172
rect 248643 476236 248709 476237
rect 248643 476172 248644 476236
rect 248708 476172 248709 476236
rect 248643 476171 248709 476172
rect 250851 476236 250917 476237
rect 250851 476172 250852 476236
rect 250916 476172 250917 476236
rect 250851 476171 250917 476172
rect 252323 476236 252389 476237
rect 252323 476172 252324 476236
rect 252388 476172 252389 476236
rect 252323 476171 252389 476172
rect 253427 476236 253493 476237
rect 253427 476172 253428 476236
rect 253492 476172 253493 476236
rect 253427 476171 253493 476172
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 253794 471454 254414 478000
rect 254534 476237 254594 479710
rect 255822 476373 255882 479710
rect 255819 476372 255885 476373
rect 255819 476308 255820 476372
rect 255884 476308 255885 476372
rect 255819 476307 255885 476308
rect 256190 476237 256250 479710
rect 257110 476237 257170 479710
rect 257846 479710 258148 479770
rect 258496 479770 258556 480080
rect 259448 479770 259508 480080
rect 260672 479770 260732 480080
rect 258496 479710 259194 479770
rect 259448 479710 259562 479770
rect 257846 476642 257906 479710
rect 258027 476644 258093 476645
rect 258027 476642 258028 476644
rect 257846 476582 258028 476642
rect 258027 476580 258028 476582
rect 258092 476580 258093 476644
rect 258027 476579 258093 476580
rect 254531 476236 254597 476237
rect 254531 476172 254532 476236
rect 254596 476172 254597 476236
rect 254531 476171 254597 476172
rect 256187 476236 256253 476237
rect 256187 476172 256188 476236
rect 256252 476172 256253 476236
rect 256187 476171 256253 476172
rect 257107 476236 257173 476237
rect 257107 476172 257108 476236
rect 257172 476172 257173 476236
rect 257107 476171 257173 476172
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 434302 254414 434898
rect 258294 475954 258914 478000
rect 259134 476509 259194 479710
rect 259131 476508 259197 476509
rect 259131 476444 259132 476508
rect 259196 476444 259197 476508
rect 259131 476443 259197 476444
rect 259502 476373 259562 479710
rect 260606 479710 260732 479770
rect 261080 479770 261140 480080
rect 261760 479770 261820 480080
rect 262848 479770 262908 480080
rect 261080 479710 261218 479770
rect 259499 476372 259565 476373
rect 259499 476308 259500 476372
rect 259564 476308 259565 476372
rect 259499 476307 259565 476308
rect 260606 476237 260666 479710
rect 261158 476373 261218 479710
rect 261710 479710 261820 479770
rect 262814 479710 262908 479770
rect 263528 479770 263588 480080
rect 263936 479770 263996 480080
rect 263528 479710 263610 479770
rect 261155 476372 261221 476373
rect 261155 476308 261156 476372
rect 261220 476308 261221 476372
rect 261155 476307 261221 476308
rect 261710 476237 261770 479710
rect 262814 476237 262874 479710
rect 263550 476645 263610 479710
rect 263918 479710 263996 479770
rect 265296 479770 265356 480080
rect 265976 479770 266036 480080
rect 265296 479710 265450 479770
rect 263547 476644 263613 476645
rect 263547 476580 263548 476644
rect 263612 476580 263613 476644
rect 263547 476579 263613 476580
rect 263918 476237 263978 479710
rect 265390 476373 265450 479710
rect 265942 479710 266036 479770
rect 266384 479770 266444 480080
rect 267608 479770 267668 480080
rect 266384 479710 266554 479770
rect 265387 476372 265453 476373
rect 265387 476308 265388 476372
rect 265452 476308 265453 476372
rect 265387 476307 265453 476308
rect 265942 476237 266002 479710
rect 266494 476373 266554 479710
rect 267598 479710 267668 479770
rect 268288 479770 268348 480080
rect 268696 479770 268756 480080
rect 269784 479770 269844 480080
rect 271008 479770 271068 480080
rect 268288 479710 268394 479770
rect 268696 479710 268762 479770
rect 269784 479710 269866 479770
rect 266491 476372 266557 476373
rect 266491 476308 266492 476372
rect 266556 476308 266557 476372
rect 266491 476307 266557 476308
rect 267598 476237 267658 479710
rect 268334 477325 268394 479710
rect 268331 477324 268397 477325
rect 268331 477260 268332 477324
rect 268396 477260 268397 477324
rect 268331 477259 268397 477260
rect 268702 476237 268762 479710
rect 269806 476237 269866 479710
rect 270910 479710 271068 479770
rect 271144 479770 271204 480080
rect 272232 479770 272292 480080
rect 273320 479770 273380 480080
rect 271144 479710 271338 479770
rect 270910 476373 270970 479710
rect 270907 476372 270973 476373
rect 270907 476308 270908 476372
rect 270972 476308 270973 476372
rect 270907 476307 270973 476308
rect 271278 476237 271338 479710
rect 272198 479710 272292 479770
rect 273302 479710 273380 479770
rect 273592 479770 273652 480080
rect 274408 479770 274468 480080
rect 273592 479710 273730 479770
rect 272198 476237 272258 479710
rect 273302 476373 273362 479710
rect 273670 476509 273730 479710
rect 274406 479710 274468 479770
rect 275768 479770 275828 480080
rect 276040 479770 276100 480080
rect 276992 479770 277052 480080
rect 275768 479710 275938 479770
rect 276040 479710 276122 479770
rect 273667 476508 273733 476509
rect 273667 476444 273668 476508
rect 273732 476444 273733 476508
rect 273667 476443 273733 476444
rect 273299 476372 273365 476373
rect 273299 476308 273300 476372
rect 273364 476308 273365 476372
rect 273299 476307 273365 476308
rect 274406 476237 274466 479710
rect 275878 476237 275938 479710
rect 276062 476373 276122 479710
rect 276982 479710 277052 479770
rect 278080 479770 278140 480080
rect 278488 479770 278548 480080
rect 278080 479710 278146 479770
rect 276059 476372 276125 476373
rect 276059 476308 276060 476372
rect 276124 476308 276125 476372
rect 276059 476307 276125 476308
rect 276982 476237 277042 479710
rect 278086 476373 278146 479710
rect 278454 479710 278548 479770
rect 279168 479770 279228 480080
rect 280936 479770 280996 480080
rect 283520 479770 283580 480080
rect 285968 479770 286028 480080
rect 288280 479770 288340 480080
rect 291000 479770 291060 480080
rect 279168 479710 279250 479770
rect 280936 479710 281090 479770
rect 283520 479710 283666 479770
rect 285968 479710 286058 479770
rect 278083 476372 278149 476373
rect 278083 476308 278084 476372
rect 278148 476308 278149 476372
rect 278083 476307 278149 476308
rect 278454 476237 278514 479710
rect 279190 476237 279250 479710
rect 281030 476917 281090 479710
rect 281027 476916 281093 476917
rect 281027 476852 281028 476916
rect 281092 476852 281093 476916
rect 281027 476851 281093 476852
rect 283606 476237 283666 479710
rect 285998 476237 286058 479710
rect 288206 479710 288340 479770
rect 290966 479710 291060 479770
rect 293448 479770 293508 480080
rect 295896 479770 295956 480080
rect 298480 479770 298540 480080
rect 300928 479770 300988 480080
rect 303512 479770 303572 480080
rect 293448 479710 293602 479770
rect 295896 479710 295994 479770
rect 298480 479710 298570 479770
rect 288206 476237 288266 479710
rect 260603 476236 260669 476237
rect 260603 476172 260604 476236
rect 260668 476172 260669 476236
rect 260603 476171 260669 476172
rect 261707 476236 261773 476237
rect 261707 476172 261708 476236
rect 261772 476172 261773 476236
rect 261707 476171 261773 476172
rect 262811 476236 262877 476237
rect 262811 476172 262812 476236
rect 262876 476172 262877 476236
rect 262811 476171 262877 476172
rect 263915 476236 263981 476237
rect 263915 476172 263916 476236
rect 263980 476172 263981 476236
rect 263915 476171 263981 476172
rect 265939 476236 266005 476237
rect 265939 476172 265940 476236
rect 266004 476172 266005 476236
rect 265939 476171 266005 476172
rect 267595 476236 267661 476237
rect 267595 476172 267596 476236
rect 267660 476172 267661 476236
rect 267595 476171 267661 476172
rect 268699 476236 268765 476237
rect 268699 476172 268700 476236
rect 268764 476172 268765 476236
rect 268699 476171 268765 476172
rect 269803 476236 269869 476237
rect 269803 476172 269804 476236
rect 269868 476172 269869 476236
rect 269803 476171 269869 476172
rect 271275 476236 271341 476237
rect 271275 476172 271276 476236
rect 271340 476172 271341 476236
rect 271275 476171 271341 476172
rect 272195 476236 272261 476237
rect 272195 476172 272196 476236
rect 272260 476172 272261 476236
rect 272195 476171 272261 476172
rect 274403 476236 274469 476237
rect 274403 476172 274404 476236
rect 274468 476172 274469 476236
rect 274403 476171 274469 476172
rect 275875 476236 275941 476237
rect 275875 476172 275876 476236
rect 275940 476172 275941 476236
rect 275875 476171 275941 476172
rect 276979 476236 277045 476237
rect 276979 476172 276980 476236
rect 277044 476172 277045 476236
rect 276979 476171 277045 476172
rect 278451 476236 278517 476237
rect 278451 476172 278452 476236
rect 278516 476172 278517 476236
rect 278451 476171 278517 476172
rect 279187 476236 279253 476237
rect 279187 476172 279188 476236
rect 279252 476172 279253 476236
rect 279187 476171 279253 476172
rect 283603 476236 283669 476237
rect 283603 476172 283604 476236
rect 283668 476172 283669 476236
rect 283603 476171 283669 476172
rect 285995 476236 286061 476237
rect 285995 476172 285996 476236
rect 286060 476172 286061 476236
rect 285995 476171 286061 476172
rect 288203 476236 288269 476237
rect 288203 476172 288204 476236
rect 288268 476172 288269 476236
rect 288203 476171 288269 476172
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 434302 258914 439398
rect 289794 471454 290414 478000
rect 290966 476237 291026 479710
rect 293542 476237 293602 479710
rect 290963 476236 291029 476237
rect 290963 476172 290964 476236
rect 291028 476172 291029 476236
rect 290963 476171 291029 476172
rect 293539 476236 293605 476237
rect 293539 476172 293540 476236
rect 293604 476172 293605 476236
rect 293539 476171 293605 476172
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 434302 290414 434898
rect 294294 475954 294914 478000
rect 295934 476237 295994 479710
rect 298510 476237 298570 479710
rect 300902 479710 300988 479770
rect 303478 479710 303572 479770
rect 305960 479770 306020 480080
rect 308544 479770 308604 480080
rect 310992 479770 311052 480080
rect 313440 479770 313500 480080
rect 315888 479770 315948 480080
rect 305960 479710 306114 479770
rect 308544 479710 308690 479770
rect 310992 479710 311082 479770
rect 300902 476237 300962 479710
rect 303478 476373 303538 479710
rect 306054 477053 306114 479710
rect 306051 477052 306117 477053
rect 306051 476988 306052 477052
rect 306116 476988 306117 477052
rect 306051 476987 306117 476988
rect 308630 476781 308690 479710
rect 308627 476780 308693 476781
rect 308627 476716 308628 476780
rect 308692 476716 308693 476780
rect 308627 476715 308693 476716
rect 303475 476372 303541 476373
rect 303475 476308 303476 476372
rect 303540 476308 303541 476372
rect 303475 476307 303541 476308
rect 311022 476237 311082 479710
rect 313414 479710 313500 479770
rect 315806 479710 315948 479770
rect 318472 479770 318532 480080
rect 320920 479770 320980 480080
rect 323368 479770 323428 480080
rect 318472 479710 318626 479770
rect 320920 479710 321018 479770
rect 313414 476645 313474 479710
rect 313411 476644 313477 476645
rect 313411 476580 313412 476644
rect 313476 476580 313477 476644
rect 313411 476579 313477 476580
rect 315806 476237 315866 479710
rect 318566 476509 318626 479710
rect 320958 477053 321018 479710
rect 323350 479710 323428 479770
rect 325952 479770 326012 480080
rect 325952 479710 326722 479770
rect 320955 477052 321021 477053
rect 320955 476988 320956 477052
rect 321020 476988 321021 477052
rect 320955 476987 321021 476988
rect 318563 476508 318629 476509
rect 318563 476444 318564 476508
rect 318628 476444 318629 476508
rect 318563 476443 318629 476444
rect 323350 476373 323410 479710
rect 323347 476372 323413 476373
rect 323347 476308 323348 476372
rect 323412 476308 323413 476372
rect 323347 476307 323413 476308
rect 295931 476236 295997 476237
rect 295931 476172 295932 476236
rect 295996 476172 295997 476236
rect 295931 476171 295997 476172
rect 298507 476236 298573 476237
rect 298507 476172 298508 476236
rect 298572 476172 298573 476236
rect 298507 476171 298573 476172
rect 300899 476236 300965 476237
rect 300899 476172 300900 476236
rect 300964 476172 300965 476236
rect 300899 476171 300965 476172
rect 311019 476236 311085 476237
rect 311019 476172 311020 476236
rect 311084 476172 311085 476236
rect 311019 476171 311085 476172
rect 315803 476236 315869 476237
rect 315803 476172 315804 476236
rect 315868 476172 315869 476236
rect 315803 476171 315869 476172
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 434302 294914 439398
rect 325794 471454 326414 478000
rect 326662 476237 326722 479710
rect 326659 476236 326725 476237
rect 326659 476172 326660 476236
rect 326724 476172 326725 476236
rect 326659 476171 326725 476172
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 434302 326414 434898
rect 330294 475954 330914 478000
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 439954 330914 475398
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 434302 330914 439398
rect 357294 466954 357914 478000
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 245699 431764 245765 431765
rect 245699 431700 245700 431764
rect 245764 431700 245765 431764
rect 245699 431699 245765 431700
rect 245702 430677 245762 431699
rect 357294 430954 357914 466398
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 360699 434892 360765 434893
rect 360699 434828 360700 434892
rect 360764 434828 360765 434892
rect 360699 434827 360765 434828
rect 359411 434756 359477 434757
rect 359411 434692 359412 434756
rect 359476 434692 359477 434756
rect 359411 434691 359477 434692
rect 358491 432308 358557 432309
rect 358491 432244 358492 432308
rect 358556 432244 358557 432308
rect 358491 432243 358557 432244
rect 358307 432172 358373 432173
rect 358307 432108 358308 432172
rect 358372 432108 358373 432172
rect 358307 432107 358373 432108
rect 358123 432036 358189 432037
rect 358123 431972 358124 432036
rect 358188 431972 358189 432036
rect 358123 431971 358189 431972
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 245699 430676 245765 430677
rect 245699 430612 245700 430676
rect 245764 430612 245765 430676
rect 245699 430611 245765 430612
rect 357294 430634 357914 430718
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 251968 403954 252288 403986
rect 251968 403718 252010 403954
rect 252246 403718 252288 403954
rect 251968 403634 252288 403718
rect 251968 403398 252010 403634
rect 252246 403398 252288 403634
rect 251968 403366 252288 403398
rect 282688 403954 283008 403986
rect 282688 403718 282730 403954
rect 282966 403718 283008 403954
rect 282688 403634 283008 403718
rect 282688 403398 282730 403634
rect 282966 403398 283008 403634
rect 282688 403366 283008 403398
rect 313408 403954 313728 403986
rect 313408 403718 313450 403954
rect 313686 403718 313728 403954
rect 313408 403634 313728 403718
rect 313408 403398 313450 403634
rect 313686 403398 313728 403634
rect 313408 403366 313728 403398
rect 344128 403954 344448 403986
rect 344128 403718 344170 403954
rect 344406 403718 344448 403954
rect 344128 403634 344448 403718
rect 344128 403398 344170 403634
rect 344406 403398 344448 403634
rect 344128 403366 344448 403398
rect 236608 399454 236928 399486
rect 236608 399218 236650 399454
rect 236886 399218 236928 399454
rect 236608 399134 236928 399218
rect 236608 398898 236650 399134
rect 236886 398898 236928 399134
rect 236608 398866 236928 398898
rect 267328 399454 267648 399486
rect 267328 399218 267370 399454
rect 267606 399218 267648 399454
rect 267328 399134 267648 399218
rect 267328 398898 267370 399134
rect 267606 398898 267648 399134
rect 267328 398866 267648 398898
rect 298048 399454 298368 399486
rect 298048 399218 298090 399454
rect 298326 399218 298368 399454
rect 298048 399134 298368 399218
rect 298048 398898 298090 399134
rect 298326 398898 298368 399134
rect 298048 398866 298368 398898
rect 328768 399454 329088 399486
rect 328768 399218 328810 399454
rect 329046 399218 329088 399454
rect 328768 399134 329088 399218
rect 328768 398898 328810 399134
rect 329046 398898 329088 399134
rect 328768 398866 329088 398898
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 232083 374100 232149 374101
rect 232083 374036 232084 374100
rect 232148 374036 232149 374100
rect 232083 374035 232149 374036
rect 232086 373010 232146 374035
rect 232086 372950 232698 373010
rect 232083 372740 232149 372741
rect 232083 372676 232084 372740
rect 232148 372676 232149 372740
rect 232083 372675 232149 372676
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 232086 364350 232146 372675
rect 232086 364290 232514 364350
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 245308 227414 263898
rect 231294 304954 231914 308400
rect 232454 308277 232514 364290
rect 232638 309909 232698 372950
rect 251968 367954 252288 367986
rect 251968 367718 252010 367954
rect 252246 367718 252288 367954
rect 251968 367634 252288 367718
rect 251968 367398 252010 367634
rect 252246 367398 252288 367634
rect 251968 367366 252288 367398
rect 282688 367954 283008 367986
rect 282688 367718 282730 367954
rect 282966 367718 283008 367954
rect 282688 367634 283008 367718
rect 282688 367398 282730 367634
rect 282966 367398 283008 367634
rect 282688 367366 283008 367398
rect 313408 367954 313728 367986
rect 313408 367718 313450 367954
rect 313686 367718 313728 367954
rect 313408 367634 313728 367718
rect 313408 367398 313450 367634
rect 313686 367398 313728 367634
rect 313408 367366 313728 367398
rect 344128 367954 344448 367986
rect 344128 367718 344170 367954
rect 344406 367718 344448 367954
rect 344128 367634 344448 367718
rect 344128 367398 344170 367634
rect 344406 367398 344448 367634
rect 344128 367366 344448 367398
rect 236608 363454 236928 363486
rect 236608 363218 236650 363454
rect 236886 363218 236928 363454
rect 236608 363134 236928 363218
rect 236608 362898 236650 363134
rect 236886 362898 236928 363134
rect 236608 362866 236928 362898
rect 267328 363454 267648 363486
rect 267328 363218 267370 363454
rect 267606 363218 267648 363454
rect 267328 363134 267648 363218
rect 267328 362898 267370 363134
rect 267606 362898 267648 363134
rect 267328 362866 267648 362898
rect 298048 363454 298368 363486
rect 298048 363218 298090 363454
rect 298326 363218 298368 363454
rect 298048 363134 298368 363218
rect 298048 362898 298090 363134
rect 298326 362898 298368 363134
rect 298048 362866 298368 362898
rect 328768 363454 329088 363486
rect 328768 363218 328810 363454
rect 329046 363218 329088 363454
rect 328768 363134 329088 363218
rect 328768 362898 328810 363134
rect 329046 362898 329088 363134
rect 328768 362866 329088 362898
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 251968 331954 252288 331986
rect 251968 331718 252010 331954
rect 252246 331718 252288 331954
rect 251968 331634 252288 331718
rect 251968 331398 252010 331634
rect 252246 331398 252288 331634
rect 251968 331366 252288 331398
rect 282688 331954 283008 331986
rect 282688 331718 282730 331954
rect 282966 331718 283008 331954
rect 282688 331634 283008 331718
rect 282688 331398 282730 331634
rect 282966 331398 283008 331634
rect 282688 331366 283008 331398
rect 313408 331954 313728 331986
rect 313408 331718 313450 331954
rect 313686 331718 313728 331954
rect 313408 331634 313728 331718
rect 313408 331398 313450 331634
rect 313686 331398 313728 331634
rect 313408 331366 313728 331398
rect 344128 331954 344448 331986
rect 344128 331718 344170 331954
rect 344406 331718 344448 331954
rect 344128 331634 344448 331718
rect 344128 331398 344170 331634
rect 344406 331398 344448 331634
rect 344128 331366 344448 331398
rect 236608 327454 236928 327486
rect 236608 327218 236650 327454
rect 236886 327218 236928 327454
rect 236608 327134 236928 327218
rect 236608 326898 236650 327134
rect 236886 326898 236928 327134
rect 236608 326866 236928 326898
rect 267328 327454 267648 327486
rect 267328 327218 267370 327454
rect 267606 327218 267648 327454
rect 267328 327134 267648 327218
rect 267328 326898 267370 327134
rect 267606 326898 267648 327134
rect 267328 326866 267648 326898
rect 298048 327454 298368 327486
rect 298048 327218 298090 327454
rect 298326 327218 298368 327454
rect 298048 327134 298368 327218
rect 298048 326898 298090 327134
rect 298326 326898 298368 327134
rect 298048 326866 298368 326898
rect 328768 327454 329088 327486
rect 328768 327218 328810 327454
rect 329046 327218 329088 327454
rect 328768 327134 329088 327218
rect 328768 326898 328810 327134
rect 329046 326898 329088 327134
rect 328768 326866 329088 326898
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 232635 309908 232701 309909
rect 232635 309844 232636 309908
rect 232700 309844 232701 309908
rect 232635 309843 232701 309844
rect 234475 309092 234541 309093
rect 234475 309028 234476 309092
rect 234540 309028 234541 309092
rect 234475 309027 234541 309028
rect 234478 308685 234538 309027
rect 234475 308684 234541 308685
rect 234475 308620 234476 308684
rect 234540 308620 234541 308684
rect 234475 308619 234541 308620
rect 232451 308276 232517 308277
rect 232451 308212 232452 308276
rect 232516 308212 232517 308276
rect 232451 308211 232517 308212
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 245308 231914 268398
rect 244794 282454 245414 308400
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 246454 245414 281898
rect 244794 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 245414 246454
rect 244794 246134 245414 246218
rect 244794 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 245414 246134
rect 244794 245308 245414 245898
rect 249294 286954 249914 308400
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 245308 249914 250398
rect 253794 291454 254414 308400
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 245308 254414 254898
rect 258294 295954 258914 308400
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 245308 258914 259398
rect 262794 300454 263414 308400
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 245308 263414 263898
rect 267294 304954 267914 308400
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 245308 267914 268398
rect 280794 282454 281414 308400
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 246454 281414 281898
rect 280794 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 281414 246454
rect 280794 246134 281414 246218
rect 280794 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 281414 246134
rect 280794 245308 281414 245898
rect 285294 286954 285914 308400
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 245308 285914 250398
rect 289794 291454 290414 308400
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 245308 290414 254898
rect 294294 295954 294914 308400
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 245308 294914 259398
rect 298794 300454 299414 308400
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 245308 299414 263898
rect 303294 304954 303914 308400
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 245308 303914 268398
rect 316794 282454 317414 308400
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 246454 317414 281898
rect 316794 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 317414 246454
rect 316794 246134 317414 246218
rect 316794 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 317414 246134
rect 316794 245308 317414 245898
rect 321294 286954 321914 308400
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 245308 321914 250398
rect 325794 291454 326414 308400
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 245308 326414 254898
rect 330294 295954 330914 308400
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 245308 330914 259398
rect 334794 300454 335414 308400
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 245308 335414 263898
rect 339294 304954 339914 308400
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 245308 339914 268398
rect 352794 282454 353414 308400
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 245308 353414 245898
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 245308 357914 250398
rect 220272 223954 220620 223986
rect 220272 223718 220328 223954
rect 220564 223718 220620 223954
rect 220272 223634 220620 223718
rect 220272 223398 220328 223634
rect 220564 223398 220620 223634
rect 220272 223366 220620 223398
rect 356000 223954 356348 223986
rect 356000 223718 356056 223954
rect 356292 223718 356348 223954
rect 356000 223634 356348 223718
rect 356000 223398 356056 223634
rect 356292 223398 356348 223634
rect 356000 223366 356348 223398
rect 220952 219454 221300 219486
rect 220952 219218 221008 219454
rect 221244 219218 221300 219454
rect 220952 219134 221300 219218
rect 220952 218898 221008 219134
rect 221244 218898 221300 219134
rect 220952 218866 221300 218898
rect 355320 219454 355668 219486
rect 355320 219218 355376 219454
rect 355612 219218 355668 219454
rect 355320 219134 355668 219218
rect 355320 218898 355376 219134
rect 355612 218898 355668 219134
rect 355320 218866 355668 218898
rect 220272 187954 220620 187986
rect 220272 187718 220328 187954
rect 220564 187718 220620 187954
rect 220272 187634 220620 187718
rect 220272 187398 220328 187634
rect 220564 187398 220620 187634
rect 220272 187366 220620 187398
rect 356000 187954 356348 187986
rect 356000 187718 356056 187954
rect 356292 187718 356348 187954
rect 356000 187634 356348 187718
rect 356000 187398 356056 187634
rect 356292 187398 356348 187634
rect 356000 187366 356348 187398
rect 220952 183454 221300 183486
rect 220952 183218 221008 183454
rect 221244 183218 221300 183454
rect 220952 183134 221300 183218
rect 220952 182898 221008 183134
rect 221244 182898 221300 183134
rect 220952 182866 221300 182898
rect 355320 183454 355668 183486
rect 355320 183218 355376 183454
rect 355612 183218 355668 183454
rect 355320 183134 355668 183218
rect 355320 182898 355376 183134
rect 355612 182898 355668 183134
rect 355320 182866 355668 182898
rect 236056 159490 236116 160106
rect 237144 159490 237204 160106
rect 238232 159901 238292 160106
rect 239592 159901 239652 160106
rect 238229 159900 238295 159901
rect 238229 159836 238230 159900
rect 238294 159836 238295 159900
rect 238229 159835 238295 159836
rect 239589 159900 239655 159901
rect 239589 159836 239590 159900
rect 239654 159836 239655 159900
rect 239589 159835 239655 159836
rect 240544 159490 240604 160106
rect 241768 159901 241828 160106
rect 241765 159900 241831 159901
rect 241765 159836 241766 159900
rect 241830 159836 241831 159900
rect 241765 159835 241831 159836
rect 243128 159490 243188 160106
rect 236056 159430 236194 159490
rect 237144 159430 237298 159490
rect 240544 159430 240610 159490
rect 236134 158541 236194 159430
rect 236131 158540 236197 158541
rect 236131 158476 236132 158540
rect 236196 158476 236197 158540
rect 236131 158475 236197 158476
rect 222294 151954 222914 158000
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 219203 3636 219269 3637
rect 219203 3572 219204 3636
rect 219268 3572 219269 3636
rect 219203 3571 219269 3572
rect 213294 -7612 213326 -7376
rect 213562 -7612 213646 -7376
rect 213882 -7612 213914 -7376
rect 213294 -7696 213914 -7612
rect 213294 -7932 213326 -7696
rect 213562 -7932 213646 -7696
rect 213882 -7932 213914 -7696
rect 213294 -7964 213914 -7932
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 218651 3500 218717 3501
rect 218651 3436 218652 3500
rect 218716 3436 218717 3500
rect 218651 3435 218717 3436
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -656 218414 2898
rect 217794 -892 217826 -656
rect 218062 -892 218146 -656
rect 218382 -892 218414 -656
rect 217794 -976 218414 -892
rect 217794 -1212 217826 -976
rect 218062 -1212 218146 -976
rect 218382 -1212 218414 -976
rect 217794 -7964 218414 -1212
rect 222294 -1616 222914 7398
rect 222294 -1852 222326 -1616
rect 222562 -1852 222646 -1616
rect 222882 -1852 222914 -1616
rect 222294 -1936 222914 -1852
rect 222294 -2172 222326 -1936
rect 222562 -2172 222646 -1936
rect 222882 -2172 222914 -1936
rect 222294 -7964 222914 -2172
rect 226794 156454 227414 158000
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2576 227414 11898
rect 226794 -2812 226826 -2576
rect 227062 -2812 227146 -2576
rect 227382 -2812 227414 -2576
rect 226794 -2896 227414 -2812
rect 226794 -3132 226826 -2896
rect 227062 -3132 227146 -2896
rect 227382 -3132 227414 -2896
rect 226794 -7964 227414 -3132
rect 231294 124954 231914 158000
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3536 231914 16398
rect 231294 -3772 231326 -3536
rect 231562 -3772 231646 -3536
rect 231882 -3772 231914 -3536
rect 231294 -3856 231914 -3772
rect 231294 -4092 231326 -3856
rect 231562 -4092 231646 -3856
rect 231882 -4092 231914 -3856
rect 231294 -7964 231914 -4092
rect 235794 129454 236414 158000
rect 237238 157589 237298 159430
rect 240550 158677 240610 159430
rect 243126 159430 243188 159490
rect 244216 159490 244276 160106
rect 245440 159490 245500 160106
rect 246528 159490 246588 160106
rect 247616 159490 247676 160106
rect 248296 159490 248356 160106
rect 248704 159490 248764 160106
rect 244216 159430 244290 159490
rect 245440 159430 245578 159490
rect 246528 159430 246682 159490
rect 247616 159430 247786 159490
rect 240547 158676 240613 158677
rect 240547 158612 240548 158676
rect 240612 158612 240613 158676
rect 240547 158611 240613 158612
rect 243126 158269 243186 159430
rect 244230 158813 244290 159430
rect 244227 158812 244293 158813
rect 244227 158748 244228 158812
rect 244292 158748 244293 158812
rect 244227 158747 244293 158748
rect 243123 158268 243189 158269
rect 243123 158204 243124 158268
rect 243188 158204 243189 158268
rect 243123 158203 243189 158204
rect 237235 157588 237301 157589
rect 237235 157524 237236 157588
rect 237300 157524 237301 157588
rect 237235 157523 237301 157524
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4496 236414 20898
rect 235794 -4732 235826 -4496
rect 236062 -4732 236146 -4496
rect 236382 -4732 236414 -4496
rect 235794 -4816 236414 -4732
rect 235794 -5052 235826 -4816
rect 236062 -5052 236146 -4816
rect 236382 -5052 236414 -4816
rect 235794 -7964 236414 -5052
rect 240294 133954 240914 158000
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5456 240914 25398
rect 240294 -5692 240326 -5456
rect 240562 -5692 240646 -5456
rect 240882 -5692 240914 -5456
rect 240294 -5776 240914 -5692
rect 240294 -6012 240326 -5776
rect 240562 -6012 240646 -5776
rect 240882 -6012 240914 -5776
rect 240294 -7964 240914 -6012
rect 244794 138454 245414 158000
rect 245518 157453 245578 159430
rect 246622 157453 246682 159430
rect 247726 157453 247786 159430
rect 248278 159430 248356 159490
rect 248646 159430 248764 159490
rect 250064 159490 250124 160106
rect 250744 159490 250804 160106
rect 251288 159490 251348 160106
rect 252376 159490 252436 160106
rect 253464 159490 253524 160106
rect 250064 159430 250178 159490
rect 250744 159430 250914 159490
rect 251288 159430 251466 159490
rect 248278 158677 248338 159430
rect 248275 158676 248341 158677
rect 248275 158612 248276 158676
rect 248340 158612 248341 158676
rect 248275 158611 248341 158612
rect 248646 158405 248706 159430
rect 250118 158677 250178 159430
rect 250115 158676 250181 158677
rect 250115 158612 250116 158676
rect 250180 158612 250181 158676
rect 250115 158611 250181 158612
rect 248643 158404 248709 158405
rect 248643 158340 248644 158404
rect 248708 158340 248709 158404
rect 248643 158339 248709 158340
rect 250854 158133 250914 159430
rect 251406 158677 251466 159430
rect 252326 159430 252436 159490
rect 253430 159430 253524 159490
rect 253600 159490 253660 160106
rect 254552 159490 254612 160106
rect 255912 159629 255972 160106
rect 255909 159628 255975 159629
rect 255909 159564 255910 159628
rect 255974 159564 255975 159628
rect 255909 159563 255975 159564
rect 256048 159490 256108 160106
rect 253600 159430 253674 159490
rect 251403 158676 251469 158677
rect 251403 158612 251404 158676
rect 251468 158612 251469 158676
rect 251403 158611 251469 158612
rect 250851 158132 250917 158133
rect 250851 158068 250852 158132
rect 250916 158068 250917 158132
rect 250851 158067 250917 158068
rect 245515 157452 245581 157453
rect 245515 157388 245516 157452
rect 245580 157388 245581 157452
rect 245515 157387 245581 157388
rect 246619 157452 246685 157453
rect 246619 157388 246620 157452
rect 246684 157388 246685 157452
rect 246619 157387 246685 157388
rect 247723 157452 247789 157453
rect 247723 157388 247724 157452
rect 247788 157388 247789 157452
rect 247723 157387 247789 157388
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6416 245414 29898
rect 244794 -6652 244826 -6416
rect 245062 -6652 245146 -6416
rect 245382 -6652 245414 -6416
rect 244794 -6736 245414 -6652
rect 244794 -6972 244826 -6736
rect 245062 -6972 245146 -6736
rect 245382 -6972 245414 -6736
rect 244794 -7964 245414 -6972
rect 249294 142954 249914 158000
rect 252326 157997 252386 159430
rect 253430 157997 253490 159430
rect 252323 157996 252389 157997
rect 252323 157932 252324 157996
rect 252388 157932 252389 157996
rect 252323 157931 252389 157932
rect 253427 157996 253493 157997
rect 253427 157932 253428 157996
rect 253492 157932 253493 157996
rect 253427 157931 253493 157932
rect 253614 157453 253674 159430
rect 254534 159430 254612 159490
rect 256006 159430 256108 159490
rect 257000 159490 257060 160106
rect 258088 159490 258148 160106
rect 258496 159490 258556 160106
rect 259448 159490 259508 160106
rect 260672 159490 260732 160106
rect 261080 159490 261140 160106
rect 261760 159490 261820 160106
rect 262848 159490 262908 160106
rect 257000 159430 257170 159490
rect 258088 159430 258274 159490
rect 258496 159430 258642 159490
rect 259448 159430 259562 159490
rect 260672 159430 260850 159490
rect 261080 159430 261218 159490
rect 254534 158677 254594 159430
rect 256006 158677 256066 159430
rect 257110 158677 257170 159430
rect 258214 158677 258274 159430
rect 258582 158677 258642 159430
rect 259502 158677 259562 159430
rect 260790 158949 260850 159430
rect 260787 158948 260853 158949
rect 260787 158884 260788 158948
rect 260852 158884 260853 158948
rect 260787 158883 260853 158884
rect 261158 158677 261218 159430
rect 261710 159430 261820 159490
rect 262814 159430 262908 159490
rect 263528 159490 263588 160106
rect 263936 159490 263996 160106
rect 265296 159629 265356 160106
rect 265293 159628 265359 159629
rect 265293 159564 265294 159628
rect 265358 159564 265359 159628
rect 265293 159563 265359 159564
rect 265976 159490 266036 160106
rect 263528 159430 263610 159490
rect 261710 159085 261770 159430
rect 261707 159084 261773 159085
rect 261707 159020 261708 159084
rect 261772 159020 261773 159084
rect 261707 159019 261773 159020
rect 262814 158677 262874 159430
rect 254531 158676 254597 158677
rect 254531 158612 254532 158676
rect 254596 158612 254597 158676
rect 254531 158611 254597 158612
rect 256003 158676 256069 158677
rect 256003 158612 256004 158676
rect 256068 158612 256069 158676
rect 256003 158611 256069 158612
rect 257107 158676 257173 158677
rect 257107 158612 257108 158676
rect 257172 158612 257173 158676
rect 257107 158611 257173 158612
rect 258211 158676 258277 158677
rect 258211 158612 258212 158676
rect 258276 158612 258277 158676
rect 258211 158611 258277 158612
rect 258579 158676 258645 158677
rect 258579 158612 258580 158676
rect 258644 158612 258645 158676
rect 258579 158611 258645 158612
rect 259499 158676 259565 158677
rect 259499 158612 259500 158676
rect 259564 158612 259565 158676
rect 259499 158611 259565 158612
rect 261155 158676 261221 158677
rect 261155 158612 261156 158676
rect 261220 158612 261221 158676
rect 261155 158611 261221 158612
rect 262811 158676 262877 158677
rect 262811 158612 262812 158676
rect 262876 158612 262877 158676
rect 262811 158611 262877 158612
rect 253611 157452 253677 157453
rect 253611 157388 253612 157452
rect 253676 157388 253677 157452
rect 253611 157387 253677 157388
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7376 249914 34398
rect 249294 -7612 249326 -7376
rect 249562 -7612 249646 -7376
rect 249882 -7612 249914 -7376
rect 249294 -7696 249914 -7612
rect 249294 -7932 249326 -7696
rect 249562 -7932 249646 -7696
rect 249882 -7932 249914 -7696
rect 249294 -7964 249914 -7932
rect 253794 147454 254414 158000
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -656 254414 2898
rect 253794 -892 253826 -656
rect 254062 -892 254146 -656
rect 254382 -892 254414 -656
rect 253794 -976 254414 -892
rect 253794 -1212 253826 -976
rect 254062 -1212 254146 -976
rect 254382 -1212 254414 -976
rect 253794 -7964 254414 -1212
rect 258294 151954 258914 158000
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1616 258914 7398
rect 258294 -1852 258326 -1616
rect 258562 -1852 258646 -1616
rect 258882 -1852 258914 -1616
rect 258294 -1936 258914 -1852
rect 258294 -2172 258326 -1936
rect 258562 -2172 258646 -1936
rect 258882 -2172 258914 -1936
rect 258294 -7964 258914 -2172
rect 262794 156454 263414 158000
rect 263550 157453 263610 159430
rect 263918 159430 263996 159490
rect 265942 159430 266036 159490
rect 266384 159490 266444 160106
rect 267608 159490 267668 160106
rect 266384 159430 266554 159490
rect 263918 158677 263978 159430
rect 265942 158677 266002 159430
rect 266494 158677 266554 159430
rect 267598 159430 267668 159490
rect 268288 159490 268348 160106
rect 268696 159490 268756 160106
rect 269784 159490 269844 160106
rect 271008 159629 271068 160106
rect 271005 159628 271071 159629
rect 271005 159564 271006 159628
rect 271070 159564 271071 159628
rect 271005 159563 271071 159564
rect 271144 159490 271204 160106
rect 272232 159490 272292 160106
rect 273320 159490 273380 160106
rect 273592 159901 273652 160106
rect 273589 159900 273655 159901
rect 273589 159836 273590 159900
rect 273654 159836 273655 159900
rect 273589 159835 273655 159836
rect 274408 159490 274468 160106
rect 268288 159430 268394 159490
rect 268696 159430 268762 159490
rect 269784 159430 269866 159490
rect 267598 158677 267658 159430
rect 263915 158676 263981 158677
rect 263915 158612 263916 158676
rect 263980 158612 263981 158676
rect 263915 158611 263981 158612
rect 265939 158676 266005 158677
rect 265939 158612 265940 158676
rect 266004 158612 266005 158676
rect 265939 158611 266005 158612
rect 266491 158676 266557 158677
rect 266491 158612 266492 158676
rect 266556 158612 266557 158676
rect 266491 158611 266557 158612
rect 267595 158676 267661 158677
rect 267595 158612 267596 158676
rect 267660 158612 267661 158676
rect 267595 158611 267661 158612
rect 263547 157452 263613 157453
rect 263547 157388 263548 157452
rect 263612 157388 263613 157452
rect 263547 157387 263613 157388
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2576 263414 11898
rect 262794 -2812 262826 -2576
rect 263062 -2812 263146 -2576
rect 263382 -2812 263414 -2576
rect 262794 -2896 263414 -2812
rect 262794 -3132 262826 -2896
rect 263062 -3132 263146 -2896
rect 263382 -3132 263414 -2896
rect 262794 -7964 263414 -3132
rect 267294 124954 267914 158000
rect 268334 157997 268394 159430
rect 268702 158677 268762 159430
rect 269806 158677 269866 159430
rect 271094 159430 271204 159490
rect 272198 159430 272292 159490
rect 273302 159430 273380 159490
rect 274406 159430 274468 159490
rect 275768 159490 275828 160106
rect 276040 159901 276100 160106
rect 276037 159900 276103 159901
rect 276037 159836 276038 159900
rect 276102 159836 276103 159900
rect 276037 159835 276103 159836
rect 276992 159490 277052 160106
rect 275768 159430 275938 159490
rect 271094 158677 271154 159430
rect 272198 158677 272258 159430
rect 273302 158677 273362 159430
rect 274406 158677 274466 159430
rect 275878 158677 275938 159430
rect 276982 159430 277052 159490
rect 278080 159490 278140 160106
rect 278488 159901 278548 160106
rect 278485 159900 278551 159901
rect 278485 159836 278486 159900
rect 278550 159836 278551 159900
rect 278485 159835 278551 159836
rect 279168 159490 279228 160106
rect 280936 159490 280996 160106
rect 283520 159490 283580 160106
rect 285968 159490 286028 160106
rect 288280 159490 288340 160106
rect 291000 159490 291060 160106
rect 293448 159901 293508 160106
rect 295896 159901 295956 160106
rect 293445 159900 293511 159901
rect 293445 159836 293446 159900
rect 293510 159836 293511 159900
rect 293445 159835 293511 159836
rect 295893 159900 295959 159901
rect 295893 159836 295894 159900
rect 295958 159836 295959 159900
rect 295893 159835 295959 159836
rect 298480 159765 298540 160106
rect 298477 159764 298543 159765
rect 298477 159700 298478 159764
rect 298542 159700 298543 159764
rect 298477 159699 298543 159700
rect 300928 159490 300988 160106
rect 303512 159901 303572 160106
rect 303509 159900 303575 159901
rect 303509 159836 303510 159900
rect 303574 159836 303575 159900
rect 303509 159835 303575 159836
rect 278080 159430 278146 159490
rect 279168 159430 279250 159490
rect 280936 159430 281090 159490
rect 283520 159430 283666 159490
rect 285968 159430 286058 159490
rect 268699 158676 268765 158677
rect 268699 158612 268700 158676
rect 268764 158612 268765 158676
rect 268699 158611 268765 158612
rect 269803 158676 269869 158677
rect 269803 158612 269804 158676
rect 269868 158612 269869 158676
rect 269803 158611 269869 158612
rect 271091 158676 271157 158677
rect 271091 158612 271092 158676
rect 271156 158612 271157 158676
rect 271091 158611 271157 158612
rect 272195 158676 272261 158677
rect 272195 158612 272196 158676
rect 272260 158612 272261 158676
rect 272195 158611 272261 158612
rect 273299 158676 273365 158677
rect 273299 158612 273300 158676
rect 273364 158612 273365 158676
rect 273299 158611 273365 158612
rect 274403 158676 274469 158677
rect 274403 158612 274404 158676
rect 274468 158612 274469 158676
rect 274403 158611 274469 158612
rect 275875 158676 275941 158677
rect 275875 158612 275876 158676
rect 275940 158612 275941 158676
rect 275875 158611 275941 158612
rect 276982 158133 277042 159430
rect 278086 158133 278146 159430
rect 279190 158133 279250 159430
rect 281030 158677 281090 159430
rect 281027 158676 281093 158677
rect 281027 158612 281028 158676
rect 281092 158612 281093 158676
rect 281027 158611 281093 158612
rect 276979 158132 277045 158133
rect 276979 158068 276980 158132
rect 277044 158068 277045 158132
rect 276979 158067 277045 158068
rect 278083 158132 278149 158133
rect 278083 158068 278084 158132
rect 278148 158068 278149 158132
rect 278083 158067 278149 158068
rect 279187 158132 279253 158133
rect 279187 158068 279188 158132
rect 279252 158068 279253 158132
rect 279187 158067 279253 158068
rect 268331 157996 268397 157997
rect 268331 157932 268332 157996
rect 268396 157932 268397 157996
rect 268331 157931 268397 157932
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3536 267914 16398
rect 267294 -3772 267326 -3536
rect 267562 -3772 267646 -3536
rect 267882 -3772 267914 -3536
rect 267294 -3856 267914 -3772
rect 267294 -4092 267326 -3856
rect 267562 -4092 267646 -3856
rect 267882 -4092 267914 -3856
rect 267294 -7964 267914 -4092
rect 271794 129454 272414 158000
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4496 272414 20898
rect 271794 -4732 271826 -4496
rect 272062 -4732 272146 -4496
rect 272382 -4732 272414 -4496
rect 271794 -4816 272414 -4732
rect 271794 -5052 271826 -4816
rect 272062 -5052 272146 -4816
rect 272382 -5052 272414 -4816
rect 271794 -7964 272414 -5052
rect 276294 133954 276914 158000
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5456 276914 25398
rect 276294 -5692 276326 -5456
rect 276562 -5692 276646 -5456
rect 276882 -5692 276914 -5456
rect 276294 -5776 276914 -5692
rect 276294 -6012 276326 -5776
rect 276562 -6012 276646 -5776
rect 276882 -6012 276914 -5776
rect 276294 -7964 276914 -6012
rect 280794 138454 281414 158000
rect 283606 157861 283666 159430
rect 283603 157860 283669 157861
rect 283603 157796 283604 157860
rect 283668 157796 283669 157860
rect 283603 157795 283669 157796
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6416 281414 29898
rect 280794 -6652 280826 -6416
rect 281062 -6652 281146 -6416
rect 281382 -6652 281414 -6416
rect 280794 -6736 281414 -6652
rect 280794 -6972 280826 -6736
rect 281062 -6972 281146 -6736
rect 281382 -6972 281414 -6736
rect 280794 -7964 281414 -6972
rect 285294 142954 285914 158000
rect 285998 157861 286058 159430
rect 288206 159430 288340 159490
rect 290966 159430 291060 159490
rect 300902 159430 300988 159490
rect 305960 159490 306020 160106
rect 308544 159490 308604 160106
rect 310992 159901 311052 160106
rect 313440 159901 313500 160106
rect 310989 159900 311055 159901
rect 310989 159836 310990 159900
rect 311054 159836 311055 159900
rect 310989 159835 311055 159836
rect 313437 159900 313503 159901
rect 313437 159836 313438 159900
rect 313502 159836 313503 159900
rect 313437 159835 313503 159836
rect 315888 159490 315948 160106
rect 305960 159430 306114 159490
rect 308544 159430 308690 159490
rect 285995 157860 286061 157861
rect 285995 157796 285996 157860
rect 286060 157796 286061 157860
rect 285995 157795 286061 157796
rect 288206 157453 288266 159430
rect 290966 158677 291026 159430
rect 300902 158677 300962 159430
rect 290963 158676 291029 158677
rect 290963 158612 290964 158676
rect 291028 158612 291029 158676
rect 290963 158611 291029 158612
rect 300899 158676 300965 158677
rect 300899 158612 300900 158676
rect 300964 158612 300965 158676
rect 300899 158611 300965 158612
rect 288203 157452 288269 157453
rect 288203 157388 288204 157452
rect 288268 157388 288269 157452
rect 288203 157387 288269 157388
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7376 285914 34398
rect 285294 -7612 285326 -7376
rect 285562 -7612 285646 -7376
rect 285882 -7612 285914 -7376
rect 285294 -7696 285914 -7612
rect 285294 -7932 285326 -7696
rect 285562 -7932 285646 -7696
rect 285882 -7932 285914 -7696
rect 285294 -7964 285914 -7932
rect 289794 147454 290414 158000
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -656 290414 2898
rect 289794 -892 289826 -656
rect 290062 -892 290146 -656
rect 290382 -892 290414 -656
rect 289794 -976 290414 -892
rect 289794 -1212 289826 -976
rect 290062 -1212 290146 -976
rect 290382 -1212 290414 -976
rect 289794 -7964 290414 -1212
rect 294294 151954 294914 158000
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1616 294914 7398
rect 294294 -1852 294326 -1616
rect 294562 -1852 294646 -1616
rect 294882 -1852 294914 -1616
rect 294294 -1936 294914 -1852
rect 294294 -2172 294326 -1936
rect 294562 -2172 294646 -1936
rect 294882 -2172 294914 -1936
rect 294294 -7964 294914 -2172
rect 298794 156454 299414 158000
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2576 299414 11898
rect 298794 -2812 298826 -2576
rect 299062 -2812 299146 -2576
rect 299382 -2812 299414 -2576
rect 298794 -2896 299414 -2812
rect 298794 -3132 298826 -2896
rect 299062 -3132 299146 -2896
rect 299382 -3132 299414 -2896
rect 298794 -7964 299414 -3132
rect 303294 124954 303914 158000
rect 306054 157453 306114 159430
rect 308630 158677 308690 159430
rect 315806 159430 315948 159490
rect 318472 159490 318532 160106
rect 320920 159490 320980 160106
rect 323368 159490 323428 160106
rect 325952 159490 326012 160106
rect 318472 159430 318626 159490
rect 320920 159430 321018 159490
rect 308627 158676 308693 158677
rect 308627 158612 308628 158676
rect 308692 158612 308693 158676
rect 308627 158611 308693 158612
rect 306051 157452 306117 157453
rect 306051 157388 306052 157452
rect 306116 157388 306117 157452
rect 306051 157387 306117 157388
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3536 303914 16398
rect 303294 -3772 303326 -3536
rect 303562 -3772 303646 -3536
rect 303882 -3772 303914 -3536
rect 303294 -3856 303914 -3772
rect 303294 -4092 303326 -3856
rect 303562 -4092 303646 -3856
rect 303882 -4092 303914 -3856
rect 303294 -7964 303914 -4092
rect 307794 129454 308414 158000
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4496 308414 20898
rect 307794 -4732 307826 -4496
rect 308062 -4732 308146 -4496
rect 308382 -4732 308414 -4496
rect 307794 -4816 308414 -4732
rect 307794 -5052 307826 -4816
rect 308062 -5052 308146 -4816
rect 308382 -5052 308414 -4816
rect 307794 -7964 308414 -5052
rect 312294 133954 312914 158000
rect 315806 157453 315866 159430
rect 315803 157452 315869 157453
rect 315803 157388 315804 157452
rect 315868 157388 315869 157452
rect 315803 157387 315869 157388
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5456 312914 25398
rect 312294 -5692 312326 -5456
rect 312562 -5692 312646 -5456
rect 312882 -5692 312914 -5456
rect 312294 -5776 312914 -5692
rect 312294 -6012 312326 -5776
rect 312562 -6012 312646 -5776
rect 312882 -6012 312914 -5776
rect 312294 -7964 312914 -6012
rect 316794 138454 317414 158000
rect 318566 157453 318626 159430
rect 320958 158677 321018 159430
rect 323350 159430 323428 159490
rect 325926 159430 326012 159490
rect 323350 158677 323410 159430
rect 325926 158677 325986 159430
rect 320955 158676 321021 158677
rect 320955 158612 320956 158676
rect 321020 158612 321021 158676
rect 320955 158611 321021 158612
rect 323347 158676 323413 158677
rect 323347 158612 323348 158676
rect 323412 158612 323413 158676
rect 323347 158611 323413 158612
rect 325923 158676 325989 158677
rect 325923 158612 325924 158676
rect 325988 158612 325989 158676
rect 325923 158611 325989 158612
rect 318563 157452 318629 157453
rect 318563 157388 318564 157452
rect 318628 157388 318629 157452
rect 318563 157387 318629 157388
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6416 317414 29898
rect 316794 -6652 316826 -6416
rect 317062 -6652 317146 -6416
rect 317382 -6652 317414 -6416
rect 316794 -6736 317414 -6652
rect 316794 -6972 316826 -6736
rect 317062 -6972 317146 -6736
rect 317382 -6972 317414 -6736
rect 316794 -7964 317414 -6972
rect 321294 142954 321914 158000
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7376 321914 34398
rect 321294 -7612 321326 -7376
rect 321562 -7612 321646 -7376
rect 321882 -7612 321914 -7376
rect 321294 -7696 321914 -7612
rect 321294 -7932 321326 -7696
rect 321562 -7932 321646 -7696
rect 321882 -7932 321914 -7696
rect 321294 -7964 321914 -7932
rect 325794 147454 326414 158000
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -656 326414 2898
rect 325794 -892 325826 -656
rect 326062 -892 326146 -656
rect 326382 -892 326414 -656
rect 325794 -976 326414 -892
rect 325794 -1212 325826 -976
rect 326062 -1212 326146 -976
rect 326382 -1212 326414 -976
rect 325794 -7964 326414 -1212
rect 330294 151954 330914 158000
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1616 330914 7398
rect 330294 -1852 330326 -1616
rect 330562 -1852 330646 -1616
rect 330882 -1852 330914 -1616
rect 330294 -1936 330914 -1852
rect 330294 -2172 330326 -1936
rect 330562 -2172 330646 -1936
rect 330882 -2172 330914 -1936
rect 330294 -7964 330914 -2172
rect 334794 156454 335414 158000
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2576 335414 11898
rect 334794 -2812 334826 -2576
rect 335062 -2812 335146 -2576
rect 335382 -2812 335414 -2576
rect 334794 -2896 335414 -2812
rect 334794 -3132 334826 -2896
rect 335062 -3132 335146 -2896
rect 335382 -3132 335414 -2896
rect 334794 -7964 335414 -3132
rect 339294 124954 339914 158000
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3536 339914 16398
rect 339294 -3772 339326 -3536
rect 339562 -3772 339646 -3536
rect 339882 -3772 339914 -3536
rect 339294 -3856 339914 -3772
rect 339294 -4092 339326 -3856
rect 339562 -4092 339646 -3856
rect 339882 -4092 339914 -3856
rect 339294 -7964 339914 -4092
rect 343794 129454 344414 158000
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4496 344414 20898
rect 343794 -4732 343826 -4496
rect 344062 -4732 344146 -4496
rect 344382 -4732 344414 -4496
rect 343794 -4816 344414 -4732
rect 343794 -5052 343826 -4816
rect 344062 -5052 344146 -4816
rect 344382 -5052 344414 -4816
rect 343794 -7964 344414 -5052
rect 348294 133954 348914 158000
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5456 348914 25398
rect 348294 -5692 348326 -5456
rect 348562 -5692 348646 -5456
rect 348882 -5692 348914 -5456
rect 348294 -5776 348914 -5692
rect 348294 -6012 348326 -5776
rect 348562 -6012 348646 -5776
rect 348882 -6012 348914 -5776
rect 348294 -7964 348914 -6012
rect 352794 138454 353414 158000
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6416 353414 29898
rect 352794 -6652 352826 -6416
rect 353062 -6652 353146 -6416
rect 353382 -6652 353414 -6416
rect 352794 -6736 353414 -6652
rect 352794 -6972 352826 -6736
rect 353062 -6972 353146 -6736
rect 353382 -6972 353414 -6736
rect 352794 -7964 353414 -6972
rect 357294 142954 357914 158000
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 358126 71909 358186 431971
rect 358310 111893 358370 432107
rect 358494 165749 358554 432243
rect 358859 300660 358925 300661
rect 358859 300596 358860 300660
rect 358924 300596 358925 300660
rect 358859 300595 358925 300596
rect 358675 244356 358741 244357
rect 358675 244292 358676 244356
rect 358740 244292 358741 244356
rect 358675 244291 358741 244292
rect 358491 165748 358557 165749
rect 358491 165684 358492 165748
rect 358556 165684 358557 165748
rect 358491 165683 358557 165684
rect 358307 111892 358373 111893
rect 358307 111828 358308 111892
rect 358372 111828 358373 111892
rect 358307 111827 358373 111828
rect 358123 71908 358189 71909
rect 358123 71844 358124 71908
rect 358188 71844 358189 71908
rect 358123 71843 358189 71844
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7376 357914 34398
rect 358678 19413 358738 244291
rect 358675 19412 358741 19413
rect 358675 19348 358676 19412
rect 358740 19348 358741 19412
rect 358675 19347 358741 19348
rect 358862 3501 358922 300595
rect 359227 245580 359293 245581
rect 359227 245516 359228 245580
rect 359292 245516 359293 245580
rect 359227 245515 359293 245516
rect 359043 245444 359109 245445
rect 359043 245380 359044 245444
rect 359108 245380 359109 245444
rect 359043 245379 359109 245380
rect 359046 3773 359106 245379
rect 359230 3909 359290 245515
rect 359414 45661 359474 434691
rect 360147 296036 360213 296037
rect 360147 295972 360148 296036
rect 360212 295972 360213 296036
rect 360147 295971 360213 295972
rect 359411 45660 359477 45661
rect 359411 45596 359412 45660
rect 359476 45596 359477 45660
rect 359411 45595 359477 45596
rect 359227 3908 359293 3909
rect 359227 3844 359228 3908
rect 359292 3844 359293 3908
rect 359227 3843 359293 3844
rect 359043 3772 359109 3773
rect 359043 3708 359044 3772
rect 359108 3708 359109 3772
rect 359043 3707 359109 3708
rect 360150 3501 360210 295971
rect 360331 248300 360397 248301
rect 360331 248236 360332 248300
rect 360396 248236 360397 248300
rect 360331 248235 360397 248236
rect 360334 157453 360394 248235
rect 360331 157452 360397 157453
rect 360331 157388 360332 157452
rect 360396 157388 360397 157452
rect 360331 157387 360397 157388
rect 360702 85645 360762 434827
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 360883 294540 360949 294541
rect 360883 294476 360884 294540
rect 360948 294476 360949 294540
rect 360883 294475 360949 294476
rect 360699 85644 360765 85645
rect 360699 85580 360700 85644
rect 360764 85580 360765 85644
rect 360699 85579 360765 85580
rect 360886 3909 360946 294475
rect 361794 291454 362414 326898
rect 366294 706108 366914 711900
rect 366294 705872 366326 706108
rect 366562 705872 366646 706108
rect 366882 705872 366914 706108
rect 366294 705788 366914 705872
rect 366294 705552 366326 705788
rect 366562 705552 366646 705788
rect 366882 705552 366914 705788
rect 366294 691954 366914 705552
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 370794 707068 371414 711900
rect 370794 706832 370826 707068
rect 371062 706832 371146 707068
rect 371382 706832 371414 707068
rect 370794 706748 371414 706832
rect 370794 706512 370826 706748
rect 371062 706512 371146 706748
rect 371382 706512 371414 706748
rect 370794 696454 371414 706512
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 368979 436252 369045 436253
rect 368979 436188 368980 436252
rect 369044 436188 369045 436252
rect 368979 436187 369045 436188
rect 367691 436116 367757 436117
rect 367691 436052 367692 436116
rect 367756 436052 367757 436116
rect 367691 436051 367757 436052
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 362907 302972 362973 302973
rect 362907 302908 362908 302972
rect 362972 302908 362973 302972
rect 362907 302907 362973 302908
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361619 280804 361685 280805
rect 361619 280740 361620 280804
rect 361684 280740 361685 280804
rect 361619 280739 361685 280740
rect 360883 3908 360949 3909
rect 360883 3844 360884 3908
rect 360948 3844 360949 3908
rect 360883 3843 360949 3844
rect 361622 3501 361682 280739
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 362539 250884 362605 250885
rect 362539 250820 362540 250884
rect 362604 250820 362605 250884
rect 362539 250819 362605 250820
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 362542 157453 362602 250819
rect 362539 157452 362605 157453
rect 362539 157388 362540 157452
rect 362604 157388 362605 157452
rect 362539 157387 362605 157388
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 358859 3500 358925 3501
rect 358859 3436 358860 3500
rect 358924 3436 358925 3500
rect 358859 3435 358925 3436
rect 360147 3500 360213 3501
rect 360147 3436 360148 3500
rect 360212 3436 360213 3500
rect 360147 3435 360213 3436
rect 361619 3500 361685 3501
rect 361619 3436 361620 3500
rect 361684 3436 361685 3500
rect 361619 3435 361685 3436
rect 361794 3454 362414 38898
rect 362910 3501 362970 302907
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 365667 283524 365733 283525
rect 365667 283460 365668 283524
rect 365732 283460 365733 283524
rect 365667 283459 365733 283460
rect 364379 267068 364445 267069
rect 364379 267004 364380 267068
rect 364444 267004 364445 267068
rect 364379 267003 364445 267004
rect 363091 250748 363157 250749
rect 363091 250684 363092 250748
rect 363156 250684 363157 250748
rect 363091 250683 363157 250684
rect 363094 6901 363154 250683
rect 363275 250612 363341 250613
rect 363275 250548 363276 250612
rect 363340 250548 363341 250612
rect 363275 250547 363341 250548
rect 363091 6900 363157 6901
rect 363091 6836 363092 6900
rect 363156 6836 363157 6900
rect 363091 6835 363157 6836
rect 363278 6629 363338 250547
rect 363459 250476 363525 250477
rect 363459 250412 363460 250476
rect 363524 250412 363525 250476
rect 363459 250411 363525 250412
rect 363462 6765 363522 250411
rect 363459 6764 363525 6765
rect 363459 6700 363460 6764
rect 363524 6700 363525 6764
rect 363459 6699 363525 6700
rect 363275 6628 363341 6629
rect 363275 6564 363276 6628
rect 363340 6564 363341 6628
rect 363275 6563 363341 6564
rect 364382 3501 364442 267003
rect 364747 248164 364813 248165
rect 364747 248100 364748 248164
rect 364812 248100 364813 248164
rect 364747 248099 364813 248100
rect 364563 248028 364629 248029
rect 364563 247964 364564 248028
rect 364628 247964 364629 248028
rect 364563 247963 364629 247964
rect 364566 8941 364626 247963
rect 364750 9077 364810 248099
rect 364931 243540 364997 243541
rect 364931 243476 364932 243540
rect 364996 243476 364997 243540
rect 364931 243475 364997 243476
rect 364934 205597 364994 243475
rect 364931 205596 364997 205597
rect 364931 205532 364932 205596
rect 364996 205532 364997 205596
rect 364931 205531 364997 205532
rect 364747 9076 364813 9077
rect 364747 9012 364748 9076
rect 364812 9012 364813 9076
rect 364747 9011 364813 9012
rect 364563 8940 364629 8941
rect 364563 8876 364564 8940
rect 364628 8876 364629 8940
rect 364563 8875 364629 8876
rect 365670 3501 365730 283459
rect 366294 259954 366914 295398
rect 367139 265572 367205 265573
rect 367139 265508 367140 265572
rect 367204 265508 367205 265572
rect 367139 265507 367205 265508
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 357294 -7612 357326 -7376
rect 357562 -7612 357646 -7376
rect 357882 -7612 357914 -7376
rect 357294 -7696 357914 -7612
rect 357294 -7932 357326 -7696
rect 357562 -7932 357646 -7696
rect 357882 -7932 357914 -7696
rect 357294 -7964 357914 -7932
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 362907 3500 362973 3501
rect 362907 3436 362908 3500
rect 362972 3436 362973 3500
rect 362907 3435 362973 3436
rect 364379 3500 364445 3501
rect 364379 3436 364380 3500
rect 364444 3436 364445 3500
rect 364379 3435 364445 3436
rect 365667 3500 365733 3501
rect 365667 3436 365668 3500
rect 365732 3436 365733 3500
rect 365667 3435 365733 3436
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -656 362414 2898
rect 361794 -892 361826 -656
rect 362062 -892 362146 -656
rect 362382 -892 362414 -656
rect 361794 -976 362414 -892
rect 361794 -1212 361826 -976
rect 362062 -1212 362146 -976
rect 362382 -1212 362414 -976
rect 361794 -7964 362414 -1212
rect 366294 -1616 366914 7398
rect 367142 3501 367202 265507
rect 367694 59397 367754 436051
rect 368427 272508 368493 272509
rect 368427 272444 368428 272508
rect 368492 272444 368493 272508
rect 368427 272443 368493 272444
rect 367691 59396 367757 59397
rect 367691 59332 367692 59396
rect 367756 59332 367757 59396
rect 367691 59331 367757 59332
rect 368430 3501 368490 272443
rect 368611 246260 368677 246261
rect 368611 246196 368612 246260
rect 368676 246196 368677 246260
rect 368611 246195 368677 246196
rect 368614 158813 368674 246195
rect 368611 158812 368677 158813
rect 368611 158748 368612 158812
rect 368676 158748 368677 158812
rect 368611 158747 368677 158748
rect 368982 99517 369042 436187
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 369899 262852 369965 262853
rect 369899 262788 369900 262852
rect 369964 262788 369965 262852
rect 369899 262787 369965 262788
rect 368979 99516 369045 99517
rect 368979 99452 368980 99516
rect 369044 99452 369045 99516
rect 368979 99451 369045 99452
rect 369902 3501 369962 262787
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 367139 3500 367205 3501
rect 367139 3436 367140 3500
rect 367204 3436 367205 3500
rect 367139 3435 367205 3436
rect 368427 3500 368493 3501
rect 368427 3436 368428 3500
rect 368492 3436 368493 3500
rect 368427 3435 368493 3436
rect 369899 3500 369965 3501
rect 369899 3436 369900 3500
rect 369964 3436 369965 3500
rect 369899 3435 369965 3436
rect 366294 -1852 366326 -1616
rect 366562 -1852 366646 -1616
rect 366882 -1852 366914 -1616
rect 366294 -1936 366914 -1852
rect 366294 -2172 366326 -1936
rect 366562 -2172 366646 -1936
rect 366882 -2172 366914 -1936
rect 366294 -7964 366914 -2172
rect 370794 -2576 371414 11898
rect 370794 -2812 370826 -2576
rect 371062 -2812 371146 -2576
rect 371382 -2812 371414 -2576
rect 370794 -2896 371414 -2812
rect 370794 -3132 370826 -2896
rect 371062 -3132 371146 -2896
rect 371382 -3132 371414 -2896
rect 370794 -7964 371414 -3132
rect 375294 708028 375914 711900
rect 375294 707792 375326 708028
rect 375562 707792 375646 708028
rect 375882 707792 375914 708028
rect 375294 707708 375914 707792
rect 375294 707472 375326 707708
rect 375562 707472 375646 707708
rect 375882 707472 375914 707708
rect 375294 700954 375914 707472
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3536 375914 16398
rect 375294 -3772 375326 -3536
rect 375562 -3772 375646 -3536
rect 375882 -3772 375914 -3536
rect 375294 -3856 375914 -3772
rect 375294 -4092 375326 -3856
rect 375562 -4092 375646 -3856
rect 375882 -4092 375914 -3856
rect 375294 -7964 375914 -4092
rect 379794 708988 380414 711900
rect 379794 708752 379826 708988
rect 380062 708752 380146 708988
rect 380382 708752 380414 708988
rect 379794 708668 380414 708752
rect 379794 708432 379826 708668
rect 380062 708432 380146 708668
rect 380382 708432 380414 708668
rect 379794 669454 380414 708432
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4496 380414 20898
rect 379794 -4732 379826 -4496
rect 380062 -4732 380146 -4496
rect 380382 -4732 380414 -4496
rect 379794 -4816 380414 -4732
rect 379794 -5052 379826 -4816
rect 380062 -5052 380146 -4816
rect 380382 -5052 380414 -4816
rect 379794 -7964 380414 -5052
rect 384294 709948 384914 711900
rect 384294 709712 384326 709948
rect 384562 709712 384646 709948
rect 384882 709712 384914 709948
rect 384294 709628 384914 709712
rect 384294 709392 384326 709628
rect 384562 709392 384646 709628
rect 384882 709392 384914 709628
rect 384294 673954 384914 709392
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5456 384914 25398
rect 384294 -5692 384326 -5456
rect 384562 -5692 384646 -5456
rect 384882 -5692 384914 -5456
rect 384294 -5776 384914 -5692
rect 384294 -6012 384326 -5776
rect 384562 -6012 384646 -5776
rect 384882 -6012 384914 -5776
rect 384294 -7964 384914 -6012
rect 388794 710908 389414 711900
rect 388794 710672 388826 710908
rect 389062 710672 389146 710908
rect 389382 710672 389414 710908
rect 388794 710588 389414 710672
rect 388794 710352 388826 710588
rect 389062 710352 389146 710588
rect 389382 710352 389414 710588
rect 388794 678454 389414 710352
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 210454 389414 245898
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6416 389414 29898
rect 388794 -6652 388826 -6416
rect 389062 -6652 389146 -6416
rect 389382 -6652 389414 -6416
rect 388794 -6736 389414 -6652
rect 388794 -6972 388826 -6736
rect 389062 -6972 389146 -6736
rect 389382 -6972 389414 -6736
rect 388794 -7964 389414 -6972
rect 393294 711868 393914 711900
rect 393294 711632 393326 711868
rect 393562 711632 393646 711868
rect 393882 711632 393914 711868
rect 393294 711548 393914 711632
rect 393294 711312 393326 711548
rect 393562 711312 393646 711548
rect 393882 711312 393914 711548
rect 393294 682954 393914 711312
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 214954 393914 250398
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7376 393914 34398
rect 393294 -7612 393326 -7376
rect 393562 -7612 393646 -7376
rect 393882 -7612 393914 -7376
rect 393294 -7696 393914 -7612
rect 393294 -7932 393326 -7696
rect 393562 -7932 393646 -7696
rect 393882 -7932 393914 -7696
rect 393294 -7964 393914 -7932
rect 397794 705148 398414 711900
rect 397794 704912 397826 705148
rect 398062 704912 398146 705148
rect 398382 704912 398414 705148
rect 397794 704828 398414 704912
rect 397794 704592 397826 704828
rect 398062 704592 398146 704828
rect 398382 704592 398414 704828
rect 397794 687454 398414 704592
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -656 398414 2898
rect 397794 -892 397826 -656
rect 398062 -892 398146 -656
rect 398382 -892 398414 -656
rect 397794 -976 398414 -892
rect 397794 -1212 397826 -976
rect 398062 -1212 398146 -976
rect 398382 -1212 398414 -976
rect 397794 -7964 398414 -1212
rect 402294 706108 402914 711900
rect 402294 705872 402326 706108
rect 402562 705872 402646 706108
rect 402882 705872 402914 706108
rect 402294 705788 402914 705872
rect 402294 705552 402326 705788
rect 402562 705552 402646 705788
rect 402882 705552 402914 705788
rect 402294 691954 402914 705552
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1616 402914 7398
rect 402294 -1852 402326 -1616
rect 402562 -1852 402646 -1616
rect 402882 -1852 402914 -1616
rect 402294 -1936 402914 -1852
rect 402294 -2172 402326 -1936
rect 402562 -2172 402646 -1936
rect 402882 -2172 402914 -1936
rect 402294 -7964 402914 -2172
rect 406794 707068 407414 711900
rect 406794 706832 406826 707068
rect 407062 706832 407146 707068
rect 407382 706832 407414 707068
rect 406794 706748 407414 706832
rect 406794 706512 406826 706748
rect 407062 706512 407146 706748
rect 407382 706512 407414 706748
rect 406794 696454 407414 706512
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2576 407414 11898
rect 406794 -2812 406826 -2576
rect 407062 -2812 407146 -2576
rect 407382 -2812 407414 -2576
rect 406794 -2896 407414 -2812
rect 406794 -3132 406826 -2896
rect 407062 -3132 407146 -2896
rect 407382 -3132 407414 -2896
rect 406794 -7964 407414 -3132
rect 411294 708028 411914 711900
rect 411294 707792 411326 708028
rect 411562 707792 411646 708028
rect 411882 707792 411914 708028
rect 411294 707708 411914 707792
rect 411294 707472 411326 707708
rect 411562 707472 411646 707708
rect 411882 707472 411914 707708
rect 411294 700954 411914 707472
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3536 411914 16398
rect 411294 -3772 411326 -3536
rect 411562 -3772 411646 -3536
rect 411882 -3772 411914 -3536
rect 411294 -3856 411914 -3772
rect 411294 -4092 411326 -3856
rect 411562 -4092 411646 -3856
rect 411882 -4092 411914 -3856
rect 411294 -7964 411914 -4092
rect 415794 708988 416414 711900
rect 415794 708752 415826 708988
rect 416062 708752 416146 708988
rect 416382 708752 416414 708988
rect 415794 708668 416414 708752
rect 415794 708432 415826 708668
rect 416062 708432 416146 708668
rect 416382 708432 416414 708668
rect 415794 669454 416414 708432
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4496 416414 20898
rect 415794 -4732 415826 -4496
rect 416062 -4732 416146 -4496
rect 416382 -4732 416414 -4496
rect 415794 -4816 416414 -4732
rect 415794 -5052 415826 -4816
rect 416062 -5052 416146 -4816
rect 416382 -5052 416414 -4816
rect 415794 -7964 416414 -5052
rect 420294 709948 420914 711900
rect 420294 709712 420326 709948
rect 420562 709712 420646 709948
rect 420882 709712 420914 709948
rect 420294 709628 420914 709712
rect 420294 709392 420326 709628
rect 420562 709392 420646 709628
rect 420882 709392 420914 709628
rect 420294 673954 420914 709392
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5456 420914 25398
rect 420294 -5692 420326 -5456
rect 420562 -5692 420646 -5456
rect 420882 -5692 420914 -5456
rect 420294 -5776 420914 -5692
rect 420294 -6012 420326 -5776
rect 420562 -6012 420646 -5776
rect 420882 -6012 420914 -5776
rect 420294 -7964 420914 -6012
rect 424794 710908 425414 711900
rect 424794 710672 424826 710908
rect 425062 710672 425146 710908
rect 425382 710672 425414 710908
rect 424794 710588 425414 710672
rect 424794 710352 424826 710588
rect 425062 710352 425146 710588
rect 425382 710352 425414 710588
rect 424794 678454 425414 710352
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6416 425414 29898
rect 424794 -6652 424826 -6416
rect 425062 -6652 425146 -6416
rect 425382 -6652 425414 -6416
rect 424794 -6736 425414 -6652
rect 424794 -6972 424826 -6736
rect 425062 -6972 425146 -6736
rect 425382 -6972 425414 -6736
rect 424794 -7964 425414 -6972
rect 429294 711868 429914 711900
rect 429294 711632 429326 711868
rect 429562 711632 429646 711868
rect 429882 711632 429914 711868
rect 429294 711548 429914 711632
rect 429294 711312 429326 711548
rect 429562 711312 429646 711548
rect 429882 711312 429914 711548
rect 429294 682954 429914 711312
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7376 429914 34398
rect 429294 -7612 429326 -7376
rect 429562 -7612 429646 -7376
rect 429882 -7612 429914 -7376
rect 429294 -7696 429914 -7612
rect 429294 -7932 429326 -7696
rect 429562 -7932 429646 -7696
rect 429882 -7932 429914 -7696
rect 429294 -7964 429914 -7932
rect 433794 705148 434414 711900
rect 433794 704912 433826 705148
rect 434062 704912 434146 705148
rect 434382 704912 434414 705148
rect 433794 704828 434414 704912
rect 433794 704592 433826 704828
rect 434062 704592 434146 704828
rect 434382 704592 434414 704828
rect 433794 687454 434414 704592
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -656 434414 2898
rect 433794 -892 433826 -656
rect 434062 -892 434146 -656
rect 434382 -892 434414 -656
rect 433794 -976 434414 -892
rect 433794 -1212 433826 -976
rect 434062 -1212 434146 -976
rect 434382 -1212 434414 -976
rect 433794 -7964 434414 -1212
rect 438294 706108 438914 711900
rect 438294 705872 438326 706108
rect 438562 705872 438646 706108
rect 438882 705872 438914 706108
rect 438294 705788 438914 705872
rect 438294 705552 438326 705788
rect 438562 705552 438646 705788
rect 438882 705552 438914 705788
rect 438294 691954 438914 705552
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1616 438914 7398
rect 438294 -1852 438326 -1616
rect 438562 -1852 438646 -1616
rect 438882 -1852 438914 -1616
rect 438294 -1936 438914 -1852
rect 438294 -2172 438326 -1936
rect 438562 -2172 438646 -1936
rect 438882 -2172 438914 -1936
rect 438294 -7964 438914 -2172
rect 442794 707068 443414 711900
rect 442794 706832 442826 707068
rect 443062 706832 443146 707068
rect 443382 706832 443414 707068
rect 442794 706748 443414 706832
rect 442794 706512 442826 706748
rect 443062 706512 443146 706748
rect 443382 706512 443414 706748
rect 442794 696454 443414 706512
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2576 443414 11898
rect 442794 -2812 442826 -2576
rect 443062 -2812 443146 -2576
rect 443382 -2812 443414 -2576
rect 442794 -2896 443414 -2812
rect 442794 -3132 442826 -2896
rect 443062 -3132 443146 -2896
rect 443382 -3132 443414 -2896
rect 442794 -7964 443414 -3132
rect 447294 708028 447914 711900
rect 447294 707792 447326 708028
rect 447562 707792 447646 708028
rect 447882 707792 447914 708028
rect 447294 707708 447914 707792
rect 447294 707472 447326 707708
rect 447562 707472 447646 707708
rect 447882 707472 447914 707708
rect 447294 700954 447914 707472
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3536 447914 16398
rect 447294 -3772 447326 -3536
rect 447562 -3772 447646 -3536
rect 447882 -3772 447914 -3536
rect 447294 -3856 447914 -3772
rect 447294 -4092 447326 -3856
rect 447562 -4092 447646 -3856
rect 447882 -4092 447914 -3856
rect 447294 -7964 447914 -4092
rect 451794 708988 452414 711900
rect 451794 708752 451826 708988
rect 452062 708752 452146 708988
rect 452382 708752 452414 708988
rect 451794 708668 452414 708752
rect 451794 708432 451826 708668
rect 452062 708432 452146 708668
rect 452382 708432 452414 708668
rect 451794 669454 452414 708432
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4496 452414 20898
rect 451794 -4732 451826 -4496
rect 452062 -4732 452146 -4496
rect 452382 -4732 452414 -4496
rect 451794 -4816 452414 -4732
rect 451794 -5052 451826 -4816
rect 452062 -5052 452146 -4816
rect 452382 -5052 452414 -4816
rect 451794 -7964 452414 -5052
rect 456294 709948 456914 711900
rect 456294 709712 456326 709948
rect 456562 709712 456646 709948
rect 456882 709712 456914 709948
rect 456294 709628 456914 709712
rect 456294 709392 456326 709628
rect 456562 709392 456646 709628
rect 456882 709392 456914 709628
rect 456294 673954 456914 709392
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5456 456914 25398
rect 456294 -5692 456326 -5456
rect 456562 -5692 456646 -5456
rect 456882 -5692 456914 -5456
rect 456294 -5776 456914 -5692
rect 456294 -6012 456326 -5776
rect 456562 -6012 456646 -5776
rect 456882 -6012 456914 -5776
rect 456294 -7964 456914 -6012
rect 460794 710908 461414 711900
rect 460794 710672 460826 710908
rect 461062 710672 461146 710908
rect 461382 710672 461414 710908
rect 460794 710588 461414 710672
rect 460794 710352 460826 710588
rect 461062 710352 461146 710588
rect 461382 710352 461414 710588
rect 460794 678454 461414 710352
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6416 461414 29898
rect 460794 -6652 460826 -6416
rect 461062 -6652 461146 -6416
rect 461382 -6652 461414 -6416
rect 460794 -6736 461414 -6652
rect 460794 -6972 460826 -6736
rect 461062 -6972 461146 -6736
rect 461382 -6972 461414 -6736
rect 460794 -7964 461414 -6972
rect 465294 711868 465914 711900
rect 465294 711632 465326 711868
rect 465562 711632 465646 711868
rect 465882 711632 465914 711868
rect 465294 711548 465914 711632
rect 465294 711312 465326 711548
rect 465562 711312 465646 711548
rect 465882 711312 465914 711548
rect 465294 682954 465914 711312
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7376 465914 34398
rect 465294 -7612 465326 -7376
rect 465562 -7612 465646 -7376
rect 465882 -7612 465914 -7376
rect 465294 -7696 465914 -7612
rect 465294 -7932 465326 -7696
rect 465562 -7932 465646 -7696
rect 465882 -7932 465914 -7696
rect 465294 -7964 465914 -7932
rect 469794 705148 470414 711900
rect 469794 704912 469826 705148
rect 470062 704912 470146 705148
rect 470382 704912 470414 705148
rect 469794 704828 470414 704912
rect 469794 704592 469826 704828
rect 470062 704592 470146 704828
rect 470382 704592 470414 704828
rect 469794 687454 470414 704592
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -656 470414 2898
rect 469794 -892 469826 -656
rect 470062 -892 470146 -656
rect 470382 -892 470414 -656
rect 469794 -976 470414 -892
rect 469794 -1212 469826 -976
rect 470062 -1212 470146 -976
rect 470382 -1212 470414 -976
rect 469794 -7964 470414 -1212
rect 474294 706108 474914 711900
rect 474294 705872 474326 706108
rect 474562 705872 474646 706108
rect 474882 705872 474914 706108
rect 474294 705788 474914 705872
rect 474294 705552 474326 705788
rect 474562 705552 474646 705788
rect 474882 705552 474914 705788
rect 474294 691954 474914 705552
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1616 474914 7398
rect 474294 -1852 474326 -1616
rect 474562 -1852 474646 -1616
rect 474882 -1852 474914 -1616
rect 474294 -1936 474914 -1852
rect 474294 -2172 474326 -1936
rect 474562 -2172 474646 -1936
rect 474882 -2172 474914 -1936
rect 474294 -7964 474914 -2172
rect 478794 707068 479414 711900
rect 478794 706832 478826 707068
rect 479062 706832 479146 707068
rect 479382 706832 479414 707068
rect 478794 706748 479414 706832
rect 478794 706512 478826 706748
rect 479062 706512 479146 706748
rect 479382 706512 479414 706748
rect 478794 696454 479414 706512
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2576 479414 11898
rect 478794 -2812 478826 -2576
rect 479062 -2812 479146 -2576
rect 479382 -2812 479414 -2576
rect 478794 -2896 479414 -2812
rect 478794 -3132 478826 -2896
rect 479062 -3132 479146 -2896
rect 479382 -3132 479414 -2896
rect 478794 -7964 479414 -3132
rect 483294 708028 483914 711900
rect 483294 707792 483326 708028
rect 483562 707792 483646 708028
rect 483882 707792 483914 708028
rect 483294 707708 483914 707792
rect 483294 707472 483326 707708
rect 483562 707472 483646 707708
rect 483882 707472 483914 707708
rect 483294 700954 483914 707472
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3536 483914 16398
rect 483294 -3772 483326 -3536
rect 483562 -3772 483646 -3536
rect 483882 -3772 483914 -3536
rect 483294 -3856 483914 -3772
rect 483294 -4092 483326 -3856
rect 483562 -4092 483646 -3856
rect 483882 -4092 483914 -3856
rect 483294 -7964 483914 -4092
rect 487794 708988 488414 711900
rect 487794 708752 487826 708988
rect 488062 708752 488146 708988
rect 488382 708752 488414 708988
rect 487794 708668 488414 708752
rect 487794 708432 487826 708668
rect 488062 708432 488146 708668
rect 488382 708432 488414 708668
rect 487794 669454 488414 708432
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4496 488414 20898
rect 487794 -4732 487826 -4496
rect 488062 -4732 488146 -4496
rect 488382 -4732 488414 -4496
rect 487794 -4816 488414 -4732
rect 487794 -5052 487826 -4816
rect 488062 -5052 488146 -4816
rect 488382 -5052 488414 -4816
rect 487794 -7964 488414 -5052
rect 492294 709948 492914 711900
rect 492294 709712 492326 709948
rect 492562 709712 492646 709948
rect 492882 709712 492914 709948
rect 492294 709628 492914 709712
rect 492294 709392 492326 709628
rect 492562 709392 492646 709628
rect 492882 709392 492914 709628
rect 492294 673954 492914 709392
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5456 492914 25398
rect 492294 -5692 492326 -5456
rect 492562 -5692 492646 -5456
rect 492882 -5692 492914 -5456
rect 492294 -5776 492914 -5692
rect 492294 -6012 492326 -5776
rect 492562 -6012 492646 -5776
rect 492882 -6012 492914 -5776
rect 492294 -7964 492914 -6012
rect 496794 710908 497414 711900
rect 496794 710672 496826 710908
rect 497062 710672 497146 710908
rect 497382 710672 497414 710908
rect 496794 710588 497414 710672
rect 496794 710352 496826 710588
rect 497062 710352 497146 710588
rect 497382 710352 497414 710588
rect 496794 678454 497414 710352
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6416 497414 29898
rect 496794 -6652 496826 -6416
rect 497062 -6652 497146 -6416
rect 497382 -6652 497414 -6416
rect 496794 -6736 497414 -6652
rect 496794 -6972 496826 -6736
rect 497062 -6972 497146 -6736
rect 497382 -6972 497414 -6736
rect 496794 -7964 497414 -6972
rect 501294 711868 501914 711900
rect 501294 711632 501326 711868
rect 501562 711632 501646 711868
rect 501882 711632 501914 711868
rect 501294 711548 501914 711632
rect 501294 711312 501326 711548
rect 501562 711312 501646 711548
rect 501882 711312 501914 711548
rect 501294 682954 501914 711312
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7376 501914 34398
rect 501294 -7612 501326 -7376
rect 501562 -7612 501646 -7376
rect 501882 -7612 501914 -7376
rect 501294 -7696 501914 -7612
rect 501294 -7932 501326 -7696
rect 501562 -7932 501646 -7696
rect 501882 -7932 501914 -7696
rect 501294 -7964 501914 -7932
rect 505794 705148 506414 711900
rect 505794 704912 505826 705148
rect 506062 704912 506146 705148
rect 506382 704912 506414 705148
rect 505794 704828 506414 704912
rect 505794 704592 505826 704828
rect 506062 704592 506146 704828
rect 506382 704592 506414 704828
rect 505794 687454 506414 704592
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -656 506414 2898
rect 505794 -892 505826 -656
rect 506062 -892 506146 -656
rect 506382 -892 506414 -656
rect 505794 -976 506414 -892
rect 505794 -1212 505826 -976
rect 506062 -1212 506146 -976
rect 506382 -1212 506414 -976
rect 505794 -7964 506414 -1212
rect 510294 706108 510914 711900
rect 510294 705872 510326 706108
rect 510562 705872 510646 706108
rect 510882 705872 510914 706108
rect 510294 705788 510914 705872
rect 510294 705552 510326 705788
rect 510562 705552 510646 705788
rect 510882 705552 510914 705788
rect 510294 691954 510914 705552
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1616 510914 7398
rect 510294 -1852 510326 -1616
rect 510562 -1852 510646 -1616
rect 510882 -1852 510914 -1616
rect 510294 -1936 510914 -1852
rect 510294 -2172 510326 -1936
rect 510562 -2172 510646 -1936
rect 510882 -2172 510914 -1936
rect 510294 -7964 510914 -2172
rect 514794 707068 515414 711900
rect 514794 706832 514826 707068
rect 515062 706832 515146 707068
rect 515382 706832 515414 707068
rect 514794 706748 515414 706832
rect 514794 706512 514826 706748
rect 515062 706512 515146 706748
rect 515382 706512 515414 706748
rect 514794 696454 515414 706512
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2576 515414 11898
rect 514794 -2812 514826 -2576
rect 515062 -2812 515146 -2576
rect 515382 -2812 515414 -2576
rect 514794 -2896 515414 -2812
rect 514794 -3132 514826 -2896
rect 515062 -3132 515146 -2896
rect 515382 -3132 515414 -2896
rect 514794 -7964 515414 -3132
rect 519294 708028 519914 711900
rect 519294 707792 519326 708028
rect 519562 707792 519646 708028
rect 519882 707792 519914 708028
rect 519294 707708 519914 707792
rect 519294 707472 519326 707708
rect 519562 707472 519646 707708
rect 519882 707472 519914 707708
rect 519294 700954 519914 707472
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3536 519914 16398
rect 519294 -3772 519326 -3536
rect 519562 -3772 519646 -3536
rect 519882 -3772 519914 -3536
rect 519294 -3856 519914 -3772
rect 519294 -4092 519326 -3856
rect 519562 -4092 519646 -3856
rect 519882 -4092 519914 -3856
rect 519294 -7964 519914 -4092
rect 523794 708988 524414 711900
rect 523794 708752 523826 708988
rect 524062 708752 524146 708988
rect 524382 708752 524414 708988
rect 523794 708668 524414 708752
rect 523794 708432 523826 708668
rect 524062 708432 524146 708668
rect 524382 708432 524414 708668
rect 523794 669454 524414 708432
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4496 524414 20898
rect 523794 -4732 523826 -4496
rect 524062 -4732 524146 -4496
rect 524382 -4732 524414 -4496
rect 523794 -4816 524414 -4732
rect 523794 -5052 523826 -4816
rect 524062 -5052 524146 -4816
rect 524382 -5052 524414 -4816
rect 523794 -7964 524414 -5052
rect 528294 709948 528914 711900
rect 528294 709712 528326 709948
rect 528562 709712 528646 709948
rect 528882 709712 528914 709948
rect 528294 709628 528914 709712
rect 528294 709392 528326 709628
rect 528562 709392 528646 709628
rect 528882 709392 528914 709628
rect 528294 673954 528914 709392
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5456 528914 25398
rect 528294 -5692 528326 -5456
rect 528562 -5692 528646 -5456
rect 528882 -5692 528914 -5456
rect 528294 -5776 528914 -5692
rect 528294 -6012 528326 -5776
rect 528562 -6012 528646 -5776
rect 528882 -6012 528914 -5776
rect 528294 -7964 528914 -6012
rect 532794 710908 533414 711900
rect 532794 710672 532826 710908
rect 533062 710672 533146 710908
rect 533382 710672 533414 710908
rect 532794 710588 533414 710672
rect 532794 710352 532826 710588
rect 533062 710352 533146 710588
rect 533382 710352 533414 710588
rect 532794 678454 533414 710352
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6416 533414 29898
rect 532794 -6652 532826 -6416
rect 533062 -6652 533146 -6416
rect 533382 -6652 533414 -6416
rect 532794 -6736 533414 -6652
rect 532794 -6972 532826 -6736
rect 533062 -6972 533146 -6736
rect 533382 -6972 533414 -6736
rect 532794 -7964 533414 -6972
rect 537294 711868 537914 711900
rect 537294 711632 537326 711868
rect 537562 711632 537646 711868
rect 537882 711632 537914 711868
rect 537294 711548 537914 711632
rect 537294 711312 537326 711548
rect 537562 711312 537646 711548
rect 537882 711312 537914 711548
rect 537294 682954 537914 711312
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7376 537914 34398
rect 537294 -7612 537326 -7376
rect 537562 -7612 537646 -7376
rect 537882 -7612 537914 -7376
rect 537294 -7696 537914 -7612
rect 537294 -7932 537326 -7696
rect 537562 -7932 537646 -7696
rect 537882 -7932 537914 -7696
rect 537294 -7964 537914 -7932
rect 541794 705148 542414 711900
rect 541794 704912 541826 705148
rect 542062 704912 542146 705148
rect 542382 704912 542414 705148
rect 541794 704828 542414 704912
rect 541794 704592 541826 704828
rect 542062 704592 542146 704828
rect 542382 704592 542414 704828
rect 541794 687454 542414 704592
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -656 542414 2898
rect 541794 -892 541826 -656
rect 542062 -892 542146 -656
rect 542382 -892 542414 -656
rect 541794 -976 542414 -892
rect 541794 -1212 541826 -976
rect 542062 -1212 542146 -976
rect 542382 -1212 542414 -976
rect 541794 -7964 542414 -1212
rect 546294 706108 546914 711900
rect 546294 705872 546326 706108
rect 546562 705872 546646 706108
rect 546882 705872 546914 706108
rect 546294 705788 546914 705872
rect 546294 705552 546326 705788
rect 546562 705552 546646 705788
rect 546882 705552 546914 705788
rect 546294 691954 546914 705552
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1616 546914 7398
rect 546294 -1852 546326 -1616
rect 546562 -1852 546646 -1616
rect 546882 -1852 546914 -1616
rect 546294 -1936 546914 -1852
rect 546294 -2172 546326 -1936
rect 546562 -2172 546646 -1936
rect 546882 -2172 546914 -1936
rect 546294 -7964 546914 -2172
rect 550794 707068 551414 711900
rect 550794 706832 550826 707068
rect 551062 706832 551146 707068
rect 551382 706832 551414 707068
rect 550794 706748 551414 706832
rect 550794 706512 550826 706748
rect 551062 706512 551146 706748
rect 551382 706512 551414 706748
rect 550794 696454 551414 706512
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2576 551414 11898
rect 550794 -2812 550826 -2576
rect 551062 -2812 551146 -2576
rect 551382 -2812 551414 -2576
rect 550794 -2896 551414 -2812
rect 550794 -3132 550826 -2896
rect 551062 -3132 551146 -2896
rect 551382 -3132 551414 -2896
rect 550794 -7964 551414 -3132
rect 555294 708028 555914 711900
rect 555294 707792 555326 708028
rect 555562 707792 555646 708028
rect 555882 707792 555914 708028
rect 555294 707708 555914 707792
rect 555294 707472 555326 707708
rect 555562 707472 555646 707708
rect 555882 707472 555914 707708
rect 555294 700954 555914 707472
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3536 555914 16398
rect 555294 -3772 555326 -3536
rect 555562 -3772 555646 -3536
rect 555882 -3772 555914 -3536
rect 555294 -3856 555914 -3772
rect 555294 -4092 555326 -3856
rect 555562 -4092 555646 -3856
rect 555882 -4092 555914 -3856
rect 555294 -7964 555914 -4092
rect 559794 708988 560414 711900
rect 559794 708752 559826 708988
rect 560062 708752 560146 708988
rect 560382 708752 560414 708988
rect 559794 708668 560414 708752
rect 559794 708432 559826 708668
rect 560062 708432 560146 708668
rect 560382 708432 560414 708668
rect 559794 669454 560414 708432
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4496 560414 20898
rect 559794 -4732 559826 -4496
rect 560062 -4732 560146 -4496
rect 560382 -4732 560414 -4496
rect 559794 -4816 560414 -4732
rect 559794 -5052 559826 -4816
rect 560062 -5052 560146 -4816
rect 560382 -5052 560414 -4816
rect 559794 -7964 560414 -5052
rect 564294 709948 564914 711900
rect 564294 709712 564326 709948
rect 564562 709712 564646 709948
rect 564882 709712 564914 709948
rect 564294 709628 564914 709712
rect 564294 709392 564326 709628
rect 564562 709392 564646 709628
rect 564882 709392 564914 709628
rect 564294 673954 564914 709392
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5456 564914 25398
rect 564294 -5692 564326 -5456
rect 564562 -5692 564646 -5456
rect 564882 -5692 564914 -5456
rect 564294 -5776 564914 -5692
rect 564294 -6012 564326 -5776
rect 564562 -6012 564646 -5776
rect 564882 -6012 564914 -5776
rect 564294 -7964 564914 -6012
rect 568794 710908 569414 711900
rect 568794 710672 568826 710908
rect 569062 710672 569146 710908
rect 569382 710672 569414 710908
rect 568794 710588 569414 710672
rect 568794 710352 568826 710588
rect 569062 710352 569146 710588
rect 569382 710352 569414 710588
rect 568794 678454 569414 710352
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6416 569414 29898
rect 568794 -6652 568826 -6416
rect 569062 -6652 569146 -6416
rect 569382 -6652 569414 -6416
rect 568794 -6736 569414 -6652
rect 568794 -6972 568826 -6736
rect 569062 -6972 569146 -6736
rect 569382 -6972 569414 -6736
rect 568794 -7964 569414 -6972
rect 573294 711868 573914 711900
rect 573294 711632 573326 711868
rect 573562 711632 573646 711868
rect 573882 711632 573914 711868
rect 573294 711548 573914 711632
rect 573294 711312 573326 711548
rect 573562 711312 573646 711548
rect 573882 711312 573914 711548
rect 573294 682954 573914 711312
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7376 573914 34398
rect 573294 -7612 573326 -7376
rect 573562 -7612 573646 -7376
rect 573882 -7612 573914 -7376
rect 573294 -7696 573914 -7612
rect 573294 -7932 573326 -7696
rect 573562 -7932 573646 -7696
rect 573882 -7932 573914 -7696
rect 573294 -7964 573914 -7932
rect 577794 705148 578414 711900
rect 577794 704912 577826 705148
rect 578062 704912 578146 705148
rect 578382 704912 578414 705148
rect 577794 704828 578414 704912
rect 577794 704592 577826 704828
rect 578062 704592 578146 704828
rect 578382 704592 578414 704828
rect 577794 687454 578414 704592
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -656 578414 2898
rect 577794 -892 577826 -656
rect 578062 -892 578146 -656
rect 578382 -892 578414 -656
rect 577794 -976 578414 -892
rect 577794 -1212 577826 -976
rect 578062 -1212 578146 -976
rect 578382 -1212 578414 -976
rect 577794 -7964 578414 -1212
rect 582294 706108 582914 711900
rect 592340 711868 592960 711900
rect 592340 711632 592372 711868
rect 592608 711632 592692 711868
rect 592928 711632 592960 711868
rect 592340 711548 592960 711632
rect 592340 711312 592372 711548
rect 592608 711312 592692 711548
rect 592928 711312 592960 711548
rect 591380 710908 592000 710940
rect 591380 710672 591412 710908
rect 591648 710672 591732 710908
rect 591968 710672 592000 710908
rect 591380 710588 592000 710672
rect 591380 710352 591412 710588
rect 591648 710352 591732 710588
rect 591968 710352 592000 710588
rect 590420 709948 591040 709980
rect 590420 709712 590452 709948
rect 590688 709712 590772 709948
rect 591008 709712 591040 709948
rect 590420 709628 591040 709712
rect 590420 709392 590452 709628
rect 590688 709392 590772 709628
rect 591008 709392 591040 709628
rect 589460 708988 590080 709020
rect 589460 708752 589492 708988
rect 589728 708752 589812 708988
rect 590048 708752 590080 708988
rect 589460 708668 590080 708752
rect 589460 708432 589492 708668
rect 589728 708432 589812 708668
rect 590048 708432 590080 708668
rect 588500 708028 589120 708060
rect 588500 707792 588532 708028
rect 588768 707792 588852 708028
rect 589088 707792 589120 708028
rect 588500 707708 589120 707792
rect 588500 707472 588532 707708
rect 588768 707472 588852 707708
rect 589088 707472 589120 707708
rect 587540 707068 588160 707100
rect 587540 706832 587572 707068
rect 587808 706832 587892 707068
rect 588128 706832 588160 707068
rect 587540 706748 588160 706832
rect 587540 706512 587572 706748
rect 587808 706512 587892 706748
rect 588128 706512 588160 706748
rect 582294 705872 582326 706108
rect 582562 705872 582646 706108
rect 582882 705872 582914 706108
rect 582294 705788 582914 705872
rect 582294 705552 582326 705788
rect 582562 705552 582646 705788
rect 582882 705552 582914 705788
rect 582294 691954 582914 705552
rect 586580 706108 587200 706140
rect 586580 705872 586612 706108
rect 586848 705872 586932 706108
rect 587168 705872 587200 706108
rect 586580 705788 587200 705872
rect 586580 705552 586612 705788
rect 586848 705552 586932 705788
rect 587168 705552 587200 705788
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1616 582914 7398
rect 585620 705148 586240 705180
rect 585620 704912 585652 705148
rect 585888 704912 585972 705148
rect 586208 704912 586240 705148
rect 585620 704828 586240 704912
rect 585620 704592 585652 704828
rect 585888 704592 585972 704828
rect 586208 704592 586240 704828
rect 585620 687454 586240 704592
rect 585620 687218 585652 687454
rect 585888 687218 585972 687454
rect 586208 687218 586240 687454
rect 585620 687134 586240 687218
rect 585620 686898 585652 687134
rect 585888 686898 585972 687134
rect 586208 686898 586240 687134
rect 585620 651454 586240 686898
rect 585620 651218 585652 651454
rect 585888 651218 585972 651454
rect 586208 651218 586240 651454
rect 585620 651134 586240 651218
rect 585620 650898 585652 651134
rect 585888 650898 585972 651134
rect 586208 650898 586240 651134
rect 585620 615454 586240 650898
rect 585620 615218 585652 615454
rect 585888 615218 585972 615454
rect 586208 615218 586240 615454
rect 585620 615134 586240 615218
rect 585620 614898 585652 615134
rect 585888 614898 585972 615134
rect 586208 614898 586240 615134
rect 585620 579454 586240 614898
rect 585620 579218 585652 579454
rect 585888 579218 585972 579454
rect 586208 579218 586240 579454
rect 585620 579134 586240 579218
rect 585620 578898 585652 579134
rect 585888 578898 585972 579134
rect 586208 578898 586240 579134
rect 585620 543454 586240 578898
rect 585620 543218 585652 543454
rect 585888 543218 585972 543454
rect 586208 543218 586240 543454
rect 585620 543134 586240 543218
rect 585620 542898 585652 543134
rect 585888 542898 585972 543134
rect 586208 542898 586240 543134
rect 585620 507454 586240 542898
rect 585620 507218 585652 507454
rect 585888 507218 585972 507454
rect 586208 507218 586240 507454
rect 585620 507134 586240 507218
rect 585620 506898 585652 507134
rect 585888 506898 585972 507134
rect 586208 506898 586240 507134
rect 585620 471454 586240 506898
rect 585620 471218 585652 471454
rect 585888 471218 585972 471454
rect 586208 471218 586240 471454
rect 585620 471134 586240 471218
rect 585620 470898 585652 471134
rect 585888 470898 585972 471134
rect 586208 470898 586240 471134
rect 585620 435454 586240 470898
rect 585620 435218 585652 435454
rect 585888 435218 585972 435454
rect 586208 435218 586240 435454
rect 585620 435134 586240 435218
rect 585620 434898 585652 435134
rect 585888 434898 585972 435134
rect 586208 434898 586240 435134
rect 585620 399454 586240 434898
rect 585620 399218 585652 399454
rect 585888 399218 585972 399454
rect 586208 399218 586240 399454
rect 585620 399134 586240 399218
rect 585620 398898 585652 399134
rect 585888 398898 585972 399134
rect 586208 398898 586240 399134
rect 585620 363454 586240 398898
rect 585620 363218 585652 363454
rect 585888 363218 585972 363454
rect 586208 363218 586240 363454
rect 585620 363134 586240 363218
rect 585620 362898 585652 363134
rect 585888 362898 585972 363134
rect 586208 362898 586240 363134
rect 585620 327454 586240 362898
rect 585620 327218 585652 327454
rect 585888 327218 585972 327454
rect 586208 327218 586240 327454
rect 585620 327134 586240 327218
rect 585620 326898 585652 327134
rect 585888 326898 585972 327134
rect 586208 326898 586240 327134
rect 585620 291454 586240 326898
rect 585620 291218 585652 291454
rect 585888 291218 585972 291454
rect 586208 291218 586240 291454
rect 585620 291134 586240 291218
rect 585620 290898 585652 291134
rect 585888 290898 585972 291134
rect 586208 290898 586240 291134
rect 585620 255454 586240 290898
rect 585620 255218 585652 255454
rect 585888 255218 585972 255454
rect 586208 255218 586240 255454
rect 585620 255134 586240 255218
rect 585620 254898 585652 255134
rect 585888 254898 585972 255134
rect 586208 254898 586240 255134
rect 585620 219454 586240 254898
rect 585620 219218 585652 219454
rect 585888 219218 585972 219454
rect 586208 219218 586240 219454
rect 585620 219134 586240 219218
rect 585620 218898 585652 219134
rect 585888 218898 585972 219134
rect 586208 218898 586240 219134
rect 585620 183454 586240 218898
rect 585620 183218 585652 183454
rect 585888 183218 585972 183454
rect 586208 183218 586240 183454
rect 585620 183134 586240 183218
rect 585620 182898 585652 183134
rect 585888 182898 585972 183134
rect 586208 182898 586240 183134
rect 585620 147454 586240 182898
rect 585620 147218 585652 147454
rect 585888 147218 585972 147454
rect 586208 147218 586240 147454
rect 585620 147134 586240 147218
rect 585620 146898 585652 147134
rect 585888 146898 585972 147134
rect 586208 146898 586240 147134
rect 585620 111454 586240 146898
rect 585620 111218 585652 111454
rect 585888 111218 585972 111454
rect 586208 111218 586240 111454
rect 585620 111134 586240 111218
rect 585620 110898 585652 111134
rect 585888 110898 585972 111134
rect 586208 110898 586240 111134
rect 585620 75454 586240 110898
rect 585620 75218 585652 75454
rect 585888 75218 585972 75454
rect 586208 75218 586240 75454
rect 585620 75134 586240 75218
rect 585620 74898 585652 75134
rect 585888 74898 585972 75134
rect 586208 74898 586240 75134
rect 585620 39454 586240 74898
rect 585620 39218 585652 39454
rect 585888 39218 585972 39454
rect 586208 39218 586240 39454
rect 585620 39134 586240 39218
rect 585620 38898 585652 39134
rect 585888 38898 585972 39134
rect 586208 38898 586240 39134
rect 585620 3454 586240 38898
rect 585620 3218 585652 3454
rect 585888 3218 585972 3454
rect 586208 3218 586240 3454
rect 585620 3134 586240 3218
rect 585620 2898 585652 3134
rect 585888 2898 585972 3134
rect 586208 2898 586240 3134
rect 585620 -656 586240 2898
rect 585620 -892 585652 -656
rect 585888 -892 585972 -656
rect 586208 -892 586240 -656
rect 585620 -976 586240 -892
rect 585620 -1212 585652 -976
rect 585888 -1212 585972 -976
rect 586208 -1212 586240 -976
rect 585620 -1244 586240 -1212
rect 586580 691954 587200 705552
rect 586580 691718 586612 691954
rect 586848 691718 586932 691954
rect 587168 691718 587200 691954
rect 586580 691634 587200 691718
rect 586580 691398 586612 691634
rect 586848 691398 586932 691634
rect 587168 691398 587200 691634
rect 586580 655954 587200 691398
rect 586580 655718 586612 655954
rect 586848 655718 586932 655954
rect 587168 655718 587200 655954
rect 586580 655634 587200 655718
rect 586580 655398 586612 655634
rect 586848 655398 586932 655634
rect 587168 655398 587200 655634
rect 586580 619954 587200 655398
rect 586580 619718 586612 619954
rect 586848 619718 586932 619954
rect 587168 619718 587200 619954
rect 586580 619634 587200 619718
rect 586580 619398 586612 619634
rect 586848 619398 586932 619634
rect 587168 619398 587200 619634
rect 586580 583954 587200 619398
rect 586580 583718 586612 583954
rect 586848 583718 586932 583954
rect 587168 583718 587200 583954
rect 586580 583634 587200 583718
rect 586580 583398 586612 583634
rect 586848 583398 586932 583634
rect 587168 583398 587200 583634
rect 586580 547954 587200 583398
rect 586580 547718 586612 547954
rect 586848 547718 586932 547954
rect 587168 547718 587200 547954
rect 586580 547634 587200 547718
rect 586580 547398 586612 547634
rect 586848 547398 586932 547634
rect 587168 547398 587200 547634
rect 586580 511954 587200 547398
rect 586580 511718 586612 511954
rect 586848 511718 586932 511954
rect 587168 511718 587200 511954
rect 586580 511634 587200 511718
rect 586580 511398 586612 511634
rect 586848 511398 586932 511634
rect 587168 511398 587200 511634
rect 586580 475954 587200 511398
rect 586580 475718 586612 475954
rect 586848 475718 586932 475954
rect 587168 475718 587200 475954
rect 586580 475634 587200 475718
rect 586580 475398 586612 475634
rect 586848 475398 586932 475634
rect 587168 475398 587200 475634
rect 586580 439954 587200 475398
rect 586580 439718 586612 439954
rect 586848 439718 586932 439954
rect 587168 439718 587200 439954
rect 586580 439634 587200 439718
rect 586580 439398 586612 439634
rect 586848 439398 586932 439634
rect 587168 439398 587200 439634
rect 586580 403954 587200 439398
rect 586580 403718 586612 403954
rect 586848 403718 586932 403954
rect 587168 403718 587200 403954
rect 586580 403634 587200 403718
rect 586580 403398 586612 403634
rect 586848 403398 586932 403634
rect 587168 403398 587200 403634
rect 586580 367954 587200 403398
rect 586580 367718 586612 367954
rect 586848 367718 586932 367954
rect 587168 367718 587200 367954
rect 586580 367634 587200 367718
rect 586580 367398 586612 367634
rect 586848 367398 586932 367634
rect 587168 367398 587200 367634
rect 586580 331954 587200 367398
rect 586580 331718 586612 331954
rect 586848 331718 586932 331954
rect 587168 331718 587200 331954
rect 586580 331634 587200 331718
rect 586580 331398 586612 331634
rect 586848 331398 586932 331634
rect 587168 331398 587200 331634
rect 586580 295954 587200 331398
rect 586580 295718 586612 295954
rect 586848 295718 586932 295954
rect 587168 295718 587200 295954
rect 586580 295634 587200 295718
rect 586580 295398 586612 295634
rect 586848 295398 586932 295634
rect 587168 295398 587200 295634
rect 586580 259954 587200 295398
rect 586580 259718 586612 259954
rect 586848 259718 586932 259954
rect 587168 259718 587200 259954
rect 586580 259634 587200 259718
rect 586580 259398 586612 259634
rect 586848 259398 586932 259634
rect 587168 259398 587200 259634
rect 586580 223954 587200 259398
rect 586580 223718 586612 223954
rect 586848 223718 586932 223954
rect 587168 223718 587200 223954
rect 586580 223634 587200 223718
rect 586580 223398 586612 223634
rect 586848 223398 586932 223634
rect 587168 223398 587200 223634
rect 586580 187954 587200 223398
rect 586580 187718 586612 187954
rect 586848 187718 586932 187954
rect 587168 187718 587200 187954
rect 586580 187634 587200 187718
rect 586580 187398 586612 187634
rect 586848 187398 586932 187634
rect 587168 187398 587200 187634
rect 586580 151954 587200 187398
rect 586580 151718 586612 151954
rect 586848 151718 586932 151954
rect 587168 151718 587200 151954
rect 586580 151634 587200 151718
rect 586580 151398 586612 151634
rect 586848 151398 586932 151634
rect 587168 151398 587200 151634
rect 586580 115954 587200 151398
rect 586580 115718 586612 115954
rect 586848 115718 586932 115954
rect 587168 115718 587200 115954
rect 586580 115634 587200 115718
rect 586580 115398 586612 115634
rect 586848 115398 586932 115634
rect 587168 115398 587200 115634
rect 586580 79954 587200 115398
rect 586580 79718 586612 79954
rect 586848 79718 586932 79954
rect 587168 79718 587200 79954
rect 586580 79634 587200 79718
rect 586580 79398 586612 79634
rect 586848 79398 586932 79634
rect 587168 79398 587200 79634
rect 586580 43954 587200 79398
rect 586580 43718 586612 43954
rect 586848 43718 586932 43954
rect 587168 43718 587200 43954
rect 586580 43634 587200 43718
rect 586580 43398 586612 43634
rect 586848 43398 586932 43634
rect 587168 43398 587200 43634
rect 586580 7954 587200 43398
rect 586580 7718 586612 7954
rect 586848 7718 586932 7954
rect 587168 7718 587200 7954
rect 586580 7634 587200 7718
rect 586580 7398 586612 7634
rect 586848 7398 586932 7634
rect 587168 7398 587200 7634
rect 582294 -1852 582326 -1616
rect 582562 -1852 582646 -1616
rect 582882 -1852 582914 -1616
rect 582294 -1936 582914 -1852
rect 582294 -2172 582326 -1936
rect 582562 -2172 582646 -1936
rect 582882 -2172 582914 -1936
rect 582294 -7964 582914 -2172
rect 586580 -1616 587200 7398
rect 586580 -1852 586612 -1616
rect 586848 -1852 586932 -1616
rect 587168 -1852 587200 -1616
rect 586580 -1936 587200 -1852
rect 586580 -2172 586612 -1936
rect 586848 -2172 586932 -1936
rect 587168 -2172 587200 -1936
rect 586580 -2204 587200 -2172
rect 587540 696454 588160 706512
rect 587540 696218 587572 696454
rect 587808 696218 587892 696454
rect 588128 696218 588160 696454
rect 587540 696134 588160 696218
rect 587540 695898 587572 696134
rect 587808 695898 587892 696134
rect 588128 695898 588160 696134
rect 587540 660454 588160 695898
rect 587540 660218 587572 660454
rect 587808 660218 587892 660454
rect 588128 660218 588160 660454
rect 587540 660134 588160 660218
rect 587540 659898 587572 660134
rect 587808 659898 587892 660134
rect 588128 659898 588160 660134
rect 587540 624454 588160 659898
rect 587540 624218 587572 624454
rect 587808 624218 587892 624454
rect 588128 624218 588160 624454
rect 587540 624134 588160 624218
rect 587540 623898 587572 624134
rect 587808 623898 587892 624134
rect 588128 623898 588160 624134
rect 587540 588454 588160 623898
rect 587540 588218 587572 588454
rect 587808 588218 587892 588454
rect 588128 588218 588160 588454
rect 587540 588134 588160 588218
rect 587540 587898 587572 588134
rect 587808 587898 587892 588134
rect 588128 587898 588160 588134
rect 587540 552454 588160 587898
rect 587540 552218 587572 552454
rect 587808 552218 587892 552454
rect 588128 552218 588160 552454
rect 587540 552134 588160 552218
rect 587540 551898 587572 552134
rect 587808 551898 587892 552134
rect 588128 551898 588160 552134
rect 587540 516454 588160 551898
rect 587540 516218 587572 516454
rect 587808 516218 587892 516454
rect 588128 516218 588160 516454
rect 587540 516134 588160 516218
rect 587540 515898 587572 516134
rect 587808 515898 587892 516134
rect 588128 515898 588160 516134
rect 587540 480454 588160 515898
rect 587540 480218 587572 480454
rect 587808 480218 587892 480454
rect 588128 480218 588160 480454
rect 587540 480134 588160 480218
rect 587540 479898 587572 480134
rect 587808 479898 587892 480134
rect 588128 479898 588160 480134
rect 587540 444454 588160 479898
rect 587540 444218 587572 444454
rect 587808 444218 587892 444454
rect 588128 444218 588160 444454
rect 587540 444134 588160 444218
rect 587540 443898 587572 444134
rect 587808 443898 587892 444134
rect 588128 443898 588160 444134
rect 587540 408454 588160 443898
rect 587540 408218 587572 408454
rect 587808 408218 587892 408454
rect 588128 408218 588160 408454
rect 587540 408134 588160 408218
rect 587540 407898 587572 408134
rect 587808 407898 587892 408134
rect 588128 407898 588160 408134
rect 587540 372454 588160 407898
rect 587540 372218 587572 372454
rect 587808 372218 587892 372454
rect 588128 372218 588160 372454
rect 587540 372134 588160 372218
rect 587540 371898 587572 372134
rect 587808 371898 587892 372134
rect 588128 371898 588160 372134
rect 587540 336454 588160 371898
rect 587540 336218 587572 336454
rect 587808 336218 587892 336454
rect 588128 336218 588160 336454
rect 587540 336134 588160 336218
rect 587540 335898 587572 336134
rect 587808 335898 587892 336134
rect 588128 335898 588160 336134
rect 587540 300454 588160 335898
rect 587540 300218 587572 300454
rect 587808 300218 587892 300454
rect 588128 300218 588160 300454
rect 587540 300134 588160 300218
rect 587540 299898 587572 300134
rect 587808 299898 587892 300134
rect 588128 299898 588160 300134
rect 587540 264454 588160 299898
rect 587540 264218 587572 264454
rect 587808 264218 587892 264454
rect 588128 264218 588160 264454
rect 587540 264134 588160 264218
rect 587540 263898 587572 264134
rect 587808 263898 587892 264134
rect 588128 263898 588160 264134
rect 587540 228454 588160 263898
rect 587540 228218 587572 228454
rect 587808 228218 587892 228454
rect 588128 228218 588160 228454
rect 587540 228134 588160 228218
rect 587540 227898 587572 228134
rect 587808 227898 587892 228134
rect 588128 227898 588160 228134
rect 587540 192454 588160 227898
rect 587540 192218 587572 192454
rect 587808 192218 587892 192454
rect 588128 192218 588160 192454
rect 587540 192134 588160 192218
rect 587540 191898 587572 192134
rect 587808 191898 587892 192134
rect 588128 191898 588160 192134
rect 587540 156454 588160 191898
rect 587540 156218 587572 156454
rect 587808 156218 587892 156454
rect 588128 156218 588160 156454
rect 587540 156134 588160 156218
rect 587540 155898 587572 156134
rect 587808 155898 587892 156134
rect 588128 155898 588160 156134
rect 587540 120454 588160 155898
rect 587540 120218 587572 120454
rect 587808 120218 587892 120454
rect 588128 120218 588160 120454
rect 587540 120134 588160 120218
rect 587540 119898 587572 120134
rect 587808 119898 587892 120134
rect 588128 119898 588160 120134
rect 587540 84454 588160 119898
rect 587540 84218 587572 84454
rect 587808 84218 587892 84454
rect 588128 84218 588160 84454
rect 587540 84134 588160 84218
rect 587540 83898 587572 84134
rect 587808 83898 587892 84134
rect 588128 83898 588160 84134
rect 587540 48454 588160 83898
rect 587540 48218 587572 48454
rect 587808 48218 587892 48454
rect 588128 48218 588160 48454
rect 587540 48134 588160 48218
rect 587540 47898 587572 48134
rect 587808 47898 587892 48134
rect 588128 47898 588160 48134
rect 587540 12454 588160 47898
rect 587540 12218 587572 12454
rect 587808 12218 587892 12454
rect 588128 12218 588160 12454
rect 587540 12134 588160 12218
rect 587540 11898 587572 12134
rect 587808 11898 587892 12134
rect 588128 11898 588160 12134
rect 587540 -2576 588160 11898
rect 587540 -2812 587572 -2576
rect 587808 -2812 587892 -2576
rect 588128 -2812 588160 -2576
rect 587540 -2896 588160 -2812
rect 587540 -3132 587572 -2896
rect 587808 -3132 587892 -2896
rect 588128 -3132 588160 -2896
rect 587540 -3164 588160 -3132
rect 588500 700954 589120 707472
rect 588500 700718 588532 700954
rect 588768 700718 588852 700954
rect 589088 700718 589120 700954
rect 588500 700634 589120 700718
rect 588500 700398 588532 700634
rect 588768 700398 588852 700634
rect 589088 700398 589120 700634
rect 588500 664954 589120 700398
rect 588500 664718 588532 664954
rect 588768 664718 588852 664954
rect 589088 664718 589120 664954
rect 588500 664634 589120 664718
rect 588500 664398 588532 664634
rect 588768 664398 588852 664634
rect 589088 664398 589120 664634
rect 588500 628954 589120 664398
rect 588500 628718 588532 628954
rect 588768 628718 588852 628954
rect 589088 628718 589120 628954
rect 588500 628634 589120 628718
rect 588500 628398 588532 628634
rect 588768 628398 588852 628634
rect 589088 628398 589120 628634
rect 588500 592954 589120 628398
rect 588500 592718 588532 592954
rect 588768 592718 588852 592954
rect 589088 592718 589120 592954
rect 588500 592634 589120 592718
rect 588500 592398 588532 592634
rect 588768 592398 588852 592634
rect 589088 592398 589120 592634
rect 588500 556954 589120 592398
rect 588500 556718 588532 556954
rect 588768 556718 588852 556954
rect 589088 556718 589120 556954
rect 588500 556634 589120 556718
rect 588500 556398 588532 556634
rect 588768 556398 588852 556634
rect 589088 556398 589120 556634
rect 588500 520954 589120 556398
rect 588500 520718 588532 520954
rect 588768 520718 588852 520954
rect 589088 520718 589120 520954
rect 588500 520634 589120 520718
rect 588500 520398 588532 520634
rect 588768 520398 588852 520634
rect 589088 520398 589120 520634
rect 588500 484954 589120 520398
rect 588500 484718 588532 484954
rect 588768 484718 588852 484954
rect 589088 484718 589120 484954
rect 588500 484634 589120 484718
rect 588500 484398 588532 484634
rect 588768 484398 588852 484634
rect 589088 484398 589120 484634
rect 588500 448954 589120 484398
rect 588500 448718 588532 448954
rect 588768 448718 588852 448954
rect 589088 448718 589120 448954
rect 588500 448634 589120 448718
rect 588500 448398 588532 448634
rect 588768 448398 588852 448634
rect 589088 448398 589120 448634
rect 588500 412954 589120 448398
rect 588500 412718 588532 412954
rect 588768 412718 588852 412954
rect 589088 412718 589120 412954
rect 588500 412634 589120 412718
rect 588500 412398 588532 412634
rect 588768 412398 588852 412634
rect 589088 412398 589120 412634
rect 588500 376954 589120 412398
rect 588500 376718 588532 376954
rect 588768 376718 588852 376954
rect 589088 376718 589120 376954
rect 588500 376634 589120 376718
rect 588500 376398 588532 376634
rect 588768 376398 588852 376634
rect 589088 376398 589120 376634
rect 588500 340954 589120 376398
rect 588500 340718 588532 340954
rect 588768 340718 588852 340954
rect 589088 340718 589120 340954
rect 588500 340634 589120 340718
rect 588500 340398 588532 340634
rect 588768 340398 588852 340634
rect 589088 340398 589120 340634
rect 588500 304954 589120 340398
rect 588500 304718 588532 304954
rect 588768 304718 588852 304954
rect 589088 304718 589120 304954
rect 588500 304634 589120 304718
rect 588500 304398 588532 304634
rect 588768 304398 588852 304634
rect 589088 304398 589120 304634
rect 588500 268954 589120 304398
rect 588500 268718 588532 268954
rect 588768 268718 588852 268954
rect 589088 268718 589120 268954
rect 588500 268634 589120 268718
rect 588500 268398 588532 268634
rect 588768 268398 588852 268634
rect 589088 268398 589120 268634
rect 588500 232954 589120 268398
rect 588500 232718 588532 232954
rect 588768 232718 588852 232954
rect 589088 232718 589120 232954
rect 588500 232634 589120 232718
rect 588500 232398 588532 232634
rect 588768 232398 588852 232634
rect 589088 232398 589120 232634
rect 588500 196954 589120 232398
rect 588500 196718 588532 196954
rect 588768 196718 588852 196954
rect 589088 196718 589120 196954
rect 588500 196634 589120 196718
rect 588500 196398 588532 196634
rect 588768 196398 588852 196634
rect 589088 196398 589120 196634
rect 588500 160954 589120 196398
rect 588500 160718 588532 160954
rect 588768 160718 588852 160954
rect 589088 160718 589120 160954
rect 588500 160634 589120 160718
rect 588500 160398 588532 160634
rect 588768 160398 588852 160634
rect 589088 160398 589120 160634
rect 588500 124954 589120 160398
rect 588500 124718 588532 124954
rect 588768 124718 588852 124954
rect 589088 124718 589120 124954
rect 588500 124634 589120 124718
rect 588500 124398 588532 124634
rect 588768 124398 588852 124634
rect 589088 124398 589120 124634
rect 588500 88954 589120 124398
rect 588500 88718 588532 88954
rect 588768 88718 588852 88954
rect 589088 88718 589120 88954
rect 588500 88634 589120 88718
rect 588500 88398 588532 88634
rect 588768 88398 588852 88634
rect 589088 88398 589120 88634
rect 588500 52954 589120 88398
rect 588500 52718 588532 52954
rect 588768 52718 588852 52954
rect 589088 52718 589120 52954
rect 588500 52634 589120 52718
rect 588500 52398 588532 52634
rect 588768 52398 588852 52634
rect 589088 52398 589120 52634
rect 588500 16954 589120 52398
rect 588500 16718 588532 16954
rect 588768 16718 588852 16954
rect 589088 16718 589120 16954
rect 588500 16634 589120 16718
rect 588500 16398 588532 16634
rect 588768 16398 588852 16634
rect 589088 16398 589120 16634
rect 588500 -3536 589120 16398
rect 588500 -3772 588532 -3536
rect 588768 -3772 588852 -3536
rect 589088 -3772 589120 -3536
rect 588500 -3856 589120 -3772
rect 588500 -4092 588532 -3856
rect 588768 -4092 588852 -3856
rect 589088 -4092 589120 -3856
rect 588500 -4124 589120 -4092
rect 589460 669454 590080 708432
rect 589460 669218 589492 669454
rect 589728 669218 589812 669454
rect 590048 669218 590080 669454
rect 589460 669134 590080 669218
rect 589460 668898 589492 669134
rect 589728 668898 589812 669134
rect 590048 668898 590080 669134
rect 589460 633454 590080 668898
rect 589460 633218 589492 633454
rect 589728 633218 589812 633454
rect 590048 633218 590080 633454
rect 589460 633134 590080 633218
rect 589460 632898 589492 633134
rect 589728 632898 589812 633134
rect 590048 632898 590080 633134
rect 589460 597454 590080 632898
rect 589460 597218 589492 597454
rect 589728 597218 589812 597454
rect 590048 597218 590080 597454
rect 589460 597134 590080 597218
rect 589460 596898 589492 597134
rect 589728 596898 589812 597134
rect 590048 596898 590080 597134
rect 589460 561454 590080 596898
rect 589460 561218 589492 561454
rect 589728 561218 589812 561454
rect 590048 561218 590080 561454
rect 589460 561134 590080 561218
rect 589460 560898 589492 561134
rect 589728 560898 589812 561134
rect 590048 560898 590080 561134
rect 589460 525454 590080 560898
rect 589460 525218 589492 525454
rect 589728 525218 589812 525454
rect 590048 525218 590080 525454
rect 589460 525134 590080 525218
rect 589460 524898 589492 525134
rect 589728 524898 589812 525134
rect 590048 524898 590080 525134
rect 589460 489454 590080 524898
rect 589460 489218 589492 489454
rect 589728 489218 589812 489454
rect 590048 489218 590080 489454
rect 589460 489134 590080 489218
rect 589460 488898 589492 489134
rect 589728 488898 589812 489134
rect 590048 488898 590080 489134
rect 589460 453454 590080 488898
rect 589460 453218 589492 453454
rect 589728 453218 589812 453454
rect 590048 453218 590080 453454
rect 589460 453134 590080 453218
rect 589460 452898 589492 453134
rect 589728 452898 589812 453134
rect 590048 452898 590080 453134
rect 589460 417454 590080 452898
rect 589460 417218 589492 417454
rect 589728 417218 589812 417454
rect 590048 417218 590080 417454
rect 589460 417134 590080 417218
rect 589460 416898 589492 417134
rect 589728 416898 589812 417134
rect 590048 416898 590080 417134
rect 589460 381454 590080 416898
rect 589460 381218 589492 381454
rect 589728 381218 589812 381454
rect 590048 381218 590080 381454
rect 589460 381134 590080 381218
rect 589460 380898 589492 381134
rect 589728 380898 589812 381134
rect 590048 380898 590080 381134
rect 589460 345454 590080 380898
rect 589460 345218 589492 345454
rect 589728 345218 589812 345454
rect 590048 345218 590080 345454
rect 589460 345134 590080 345218
rect 589460 344898 589492 345134
rect 589728 344898 589812 345134
rect 590048 344898 590080 345134
rect 589460 309454 590080 344898
rect 589460 309218 589492 309454
rect 589728 309218 589812 309454
rect 590048 309218 590080 309454
rect 589460 309134 590080 309218
rect 589460 308898 589492 309134
rect 589728 308898 589812 309134
rect 590048 308898 590080 309134
rect 589460 273454 590080 308898
rect 589460 273218 589492 273454
rect 589728 273218 589812 273454
rect 590048 273218 590080 273454
rect 589460 273134 590080 273218
rect 589460 272898 589492 273134
rect 589728 272898 589812 273134
rect 590048 272898 590080 273134
rect 589460 237454 590080 272898
rect 589460 237218 589492 237454
rect 589728 237218 589812 237454
rect 590048 237218 590080 237454
rect 589460 237134 590080 237218
rect 589460 236898 589492 237134
rect 589728 236898 589812 237134
rect 590048 236898 590080 237134
rect 589460 201454 590080 236898
rect 589460 201218 589492 201454
rect 589728 201218 589812 201454
rect 590048 201218 590080 201454
rect 589460 201134 590080 201218
rect 589460 200898 589492 201134
rect 589728 200898 589812 201134
rect 590048 200898 590080 201134
rect 589460 165454 590080 200898
rect 589460 165218 589492 165454
rect 589728 165218 589812 165454
rect 590048 165218 590080 165454
rect 589460 165134 590080 165218
rect 589460 164898 589492 165134
rect 589728 164898 589812 165134
rect 590048 164898 590080 165134
rect 589460 129454 590080 164898
rect 589460 129218 589492 129454
rect 589728 129218 589812 129454
rect 590048 129218 590080 129454
rect 589460 129134 590080 129218
rect 589460 128898 589492 129134
rect 589728 128898 589812 129134
rect 590048 128898 590080 129134
rect 589460 93454 590080 128898
rect 589460 93218 589492 93454
rect 589728 93218 589812 93454
rect 590048 93218 590080 93454
rect 589460 93134 590080 93218
rect 589460 92898 589492 93134
rect 589728 92898 589812 93134
rect 590048 92898 590080 93134
rect 589460 57454 590080 92898
rect 589460 57218 589492 57454
rect 589728 57218 589812 57454
rect 590048 57218 590080 57454
rect 589460 57134 590080 57218
rect 589460 56898 589492 57134
rect 589728 56898 589812 57134
rect 590048 56898 590080 57134
rect 589460 21454 590080 56898
rect 589460 21218 589492 21454
rect 589728 21218 589812 21454
rect 590048 21218 590080 21454
rect 589460 21134 590080 21218
rect 589460 20898 589492 21134
rect 589728 20898 589812 21134
rect 590048 20898 590080 21134
rect 589460 -4496 590080 20898
rect 589460 -4732 589492 -4496
rect 589728 -4732 589812 -4496
rect 590048 -4732 590080 -4496
rect 589460 -4816 590080 -4732
rect 589460 -5052 589492 -4816
rect 589728 -5052 589812 -4816
rect 590048 -5052 590080 -4816
rect 589460 -5084 590080 -5052
rect 590420 673954 591040 709392
rect 590420 673718 590452 673954
rect 590688 673718 590772 673954
rect 591008 673718 591040 673954
rect 590420 673634 591040 673718
rect 590420 673398 590452 673634
rect 590688 673398 590772 673634
rect 591008 673398 591040 673634
rect 590420 637954 591040 673398
rect 590420 637718 590452 637954
rect 590688 637718 590772 637954
rect 591008 637718 591040 637954
rect 590420 637634 591040 637718
rect 590420 637398 590452 637634
rect 590688 637398 590772 637634
rect 591008 637398 591040 637634
rect 590420 601954 591040 637398
rect 590420 601718 590452 601954
rect 590688 601718 590772 601954
rect 591008 601718 591040 601954
rect 590420 601634 591040 601718
rect 590420 601398 590452 601634
rect 590688 601398 590772 601634
rect 591008 601398 591040 601634
rect 590420 565954 591040 601398
rect 590420 565718 590452 565954
rect 590688 565718 590772 565954
rect 591008 565718 591040 565954
rect 590420 565634 591040 565718
rect 590420 565398 590452 565634
rect 590688 565398 590772 565634
rect 591008 565398 591040 565634
rect 590420 529954 591040 565398
rect 590420 529718 590452 529954
rect 590688 529718 590772 529954
rect 591008 529718 591040 529954
rect 590420 529634 591040 529718
rect 590420 529398 590452 529634
rect 590688 529398 590772 529634
rect 591008 529398 591040 529634
rect 590420 493954 591040 529398
rect 590420 493718 590452 493954
rect 590688 493718 590772 493954
rect 591008 493718 591040 493954
rect 590420 493634 591040 493718
rect 590420 493398 590452 493634
rect 590688 493398 590772 493634
rect 591008 493398 591040 493634
rect 590420 457954 591040 493398
rect 590420 457718 590452 457954
rect 590688 457718 590772 457954
rect 591008 457718 591040 457954
rect 590420 457634 591040 457718
rect 590420 457398 590452 457634
rect 590688 457398 590772 457634
rect 591008 457398 591040 457634
rect 590420 421954 591040 457398
rect 590420 421718 590452 421954
rect 590688 421718 590772 421954
rect 591008 421718 591040 421954
rect 590420 421634 591040 421718
rect 590420 421398 590452 421634
rect 590688 421398 590772 421634
rect 591008 421398 591040 421634
rect 590420 385954 591040 421398
rect 590420 385718 590452 385954
rect 590688 385718 590772 385954
rect 591008 385718 591040 385954
rect 590420 385634 591040 385718
rect 590420 385398 590452 385634
rect 590688 385398 590772 385634
rect 591008 385398 591040 385634
rect 590420 349954 591040 385398
rect 590420 349718 590452 349954
rect 590688 349718 590772 349954
rect 591008 349718 591040 349954
rect 590420 349634 591040 349718
rect 590420 349398 590452 349634
rect 590688 349398 590772 349634
rect 591008 349398 591040 349634
rect 590420 313954 591040 349398
rect 590420 313718 590452 313954
rect 590688 313718 590772 313954
rect 591008 313718 591040 313954
rect 590420 313634 591040 313718
rect 590420 313398 590452 313634
rect 590688 313398 590772 313634
rect 591008 313398 591040 313634
rect 590420 277954 591040 313398
rect 590420 277718 590452 277954
rect 590688 277718 590772 277954
rect 591008 277718 591040 277954
rect 590420 277634 591040 277718
rect 590420 277398 590452 277634
rect 590688 277398 590772 277634
rect 591008 277398 591040 277634
rect 590420 241954 591040 277398
rect 590420 241718 590452 241954
rect 590688 241718 590772 241954
rect 591008 241718 591040 241954
rect 590420 241634 591040 241718
rect 590420 241398 590452 241634
rect 590688 241398 590772 241634
rect 591008 241398 591040 241634
rect 590420 205954 591040 241398
rect 590420 205718 590452 205954
rect 590688 205718 590772 205954
rect 591008 205718 591040 205954
rect 590420 205634 591040 205718
rect 590420 205398 590452 205634
rect 590688 205398 590772 205634
rect 591008 205398 591040 205634
rect 590420 169954 591040 205398
rect 590420 169718 590452 169954
rect 590688 169718 590772 169954
rect 591008 169718 591040 169954
rect 590420 169634 591040 169718
rect 590420 169398 590452 169634
rect 590688 169398 590772 169634
rect 591008 169398 591040 169634
rect 590420 133954 591040 169398
rect 590420 133718 590452 133954
rect 590688 133718 590772 133954
rect 591008 133718 591040 133954
rect 590420 133634 591040 133718
rect 590420 133398 590452 133634
rect 590688 133398 590772 133634
rect 591008 133398 591040 133634
rect 590420 97954 591040 133398
rect 590420 97718 590452 97954
rect 590688 97718 590772 97954
rect 591008 97718 591040 97954
rect 590420 97634 591040 97718
rect 590420 97398 590452 97634
rect 590688 97398 590772 97634
rect 591008 97398 591040 97634
rect 590420 61954 591040 97398
rect 590420 61718 590452 61954
rect 590688 61718 590772 61954
rect 591008 61718 591040 61954
rect 590420 61634 591040 61718
rect 590420 61398 590452 61634
rect 590688 61398 590772 61634
rect 591008 61398 591040 61634
rect 590420 25954 591040 61398
rect 590420 25718 590452 25954
rect 590688 25718 590772 25954
rect 591008 25718 591040 25954
rect 590420 25634 591040 25718
rect 590420 25398 590452 25634
rect 590688 25398 590772 25634
rect 591008 25398 591040 25634
rect 590420 -5456 591040 25398
rect 590420 -5692 590452 -5456
rect 590688 -5692 590772 -5456
rect 591008 -5692 591040 -5456
rect 590420 -5776 591040 -5692
rect 590420 -6012 590452 -5776
rect 590688 -6012 590772 -5776
rect 591008 -6012 591040 -5776
rect 590420 -6044 591040 -6012
rect 591380 678454 592000 710352
rect 591380 678218 591412 678454
rect 591648 678218 591732 678454
rect 591968 678218 592000 678454
rect 591380 678134 592000 678218
rect 591380 677898 591412 678134
rect 591648 677898 591732 678134
rect 591968 677898 592000 678134
rect 591380 642454 592000 677898
rect 591380 642218 591412 642454
rect 591648 642218 591732 642454
rect 591968 642218 592000 642454
rect 591380 642134 592000 642218
rect 591380 641898 591412 642134
rect 591648 641898 591732 642134
rect 591968 641898 592000 642134
rect 591380 606454 592000 641898
rect 591380 606218 591412 606454
rect 591648 606218 591732 606454
rect 591968 606218 592000 606454
rect 591380 606134 592000 606218
rect 591380 605898 591412 606134
rect 591648 605898 591732 606134
rect 591968 605898 592000 606134
rect 591380 570454 592000 605898
rect 591380 570218 591412 570454
rect 591648 570218 591732 570454
rect 591968 570218 592000 570454
rect 591380 570134 592000 570218
rect 591380 569898 591412 570134
rect 591648 569898 591732 570134
rect 591968 569898 592000 570134
rect 591380 534454 592000 569898
rect 591380 534218 591412 534454
rect 591648 534218 591732 534454
rect 591968 534218 592000 534454
rect 591380 534134 592000 534218
rect 591380 533898 591412 534134
rect 591648 533898 591732 534134
rect 591968 533898 592000 534134
rect 591380 498454 592000 533898
rect 591380 498218 591412 498454
rect 591648 498218 591732 498454
rect 591968 498218 592000 498454
rect 591380 498134 592000 498218
rect 591380 497898 591412 498134
rect 591648 497898 591732 498134
rect 591968 497898 592000 498134
rect 591380 462454 592000 497898
rect 591380 462218 591412 462454
rect 591648 462218 591732 462454
rect 591968 462218 592000 462454
rect 591380 462134 592000 462218
rect 591380 461898 591412 462134
rect 591648 461898 591732 462134
rect 591968 461898 592000 462134
rect 591380 426454 592000 461898
rect 591380 426218 591412 426454
rect 591648 426218 591732 426454
rect 591968 426218 592000 426454
rect 591380 426134 592000 426218
rect 591380 425898 591412 426134
rect 591648 425898 591732 426134
rect 591968 425898 592000 426134
rect 591380 390454 592000 425898
rect 591380 390218 591412 390454
rect 591648 390218 591732 390454
rect 591968 390218 592000 390454
rect 591380 390134 592000 390218
rect 591380 389898 591412 390134
rect 591648 389898 591732 390134
rect 591968 389898 592000 390134
rect 591380 354454 592000 389898
rect 591380 354218 591412 354454
rect 591648 354218 591732 354454
rect 591968 354218 592000 354454
rect 591380 354134 592000 354218
rect 591380 353898 591412 354134
rect 591648 353898 591732 354134
rect 591968 353898 592000 354134
rect 591380 318454 592000 353898
rect 591380 318218 591412 318454
rect 591648 318218 591732 318454
rect 591968 318218 592000 318454
rect 591380 318134 592000 318218
rect 591380 317898 591412 318134
rect 591648 317898 591732 318134
rect 591968 317898 592000 318134
rect 591380 282454 592000 317898
rect 591380 282218 591412 282454
rect 591648 282218 591732 282454
rect 591968 282218 592000 282454
rect 591380 282134 592000 282218
rect 591380 281898 591412 282134
rect 591648 281898 591732 282134
rect 591968 281898 592000 282134
rect 591380 246454 592000 281898
rect 591380 246218 591412 246454
rect 591648 246218 591732 246454
rect 591968 246218 592000 246454
rect 591380 246134 592000 246218
rect 591380 245898 591412 246134
rect 591648 245898 591732 246134
rect 591968 245898 592000 246134
rect 591380 210454 592000 245898
rect 591380 210218 591412 210454
rect 591648 210218 591732 210454
rect 591968 210218 592000 210454
rect 591380 210134 592000 210218
rect 591380 209898 591412 210134
rect 591648 209898 591732 210134
rect 591968 209898 592000 210134
rect 591380 174454 592000 209898
rect 591380 174218 591412 174454
rect 591648 174218 591732 174454
rect 591968 174218 592000 174454
rect 591380 174134 592000 174218
rect 591380 173898 591412 174134
rect 591648 173898 591732 174134
rect 591968 173898 592000 174134
rect 591380 138454 592000 173898
rect 591380 138218 591412 138454
rect 591648 138218 591732 138454
rect 591968 138218 592000 138454
rect 591380 138134 592000 138218
rect 591380 137898 591412 138134
rect 591648 137898 591732 138134
rect 591968 137898 592000 138134
rect 591380 102454 592000 137898
rect 591380 102218 591412 102454
rect 591648 102218 591732 102454
rect 591968 102218 592000 102454
rect 591380 102134 592000 102218
rect 591380 101898 591412 102134
rect 591648 101898 591732 102134
rect 591968 101898 592000 102134
rect 591380 66454 592000 101898
rect 591380 66218 591412 66454
rect 591648 66218 591732 66454
rect 591968 66218 592000 66454
rect 591380 66134 592000 66218
rect 591380 65898 591412 66134
rect 591648 65898 591732 66134
rect 591968 65898 592000 66134
rect 591380 30454 592000 65898
rect 591380 30218 591412 30454
rect 591648 30218 591732 30454
rect 591968 30218 592000 30454
rect 591380 30134 592000 30218
rect 591380 29898 591412 30134
rect 591648 29898 591732 30134
rect 591968 29898 592000 30134
rect 591380 -6416 592000 29898
rect 591380 -6652 591412 -6416
rect 591648 -6652 591732 -6416
rect 591968 -6652 592000 -6416
rect 591380 -6736 592000 -6652
rect 591380 -6972 591412 -6736
rect 591648 -6972 591732 -6736
rect 591968 -6972 592000 -6736
rect 591380 -7004 592000 -6972
rect 592340 682954 592960 711312
rect 592340 682718 592372 682954
rect 592608 682718 592692 682954
rect 592928 682718 592960 682954
rect 592340 682634 592960 682718
rect 592340 682398 592372 682634
rect 592608 682398 592692 682634
rect 592928 682398 592960 682634
rect 592340 646954 592960 682398
rect 592340 646718 592372 646954
rect 592608 646718 592692 646954
rect 592928 646718 592960 646954
rect 592340 646634 592960 646718
rect 592340 646398 592372 646634
rect 592608 646398 592692 646634
rect 592928 646398 592960 646634
rect 592340 610954 592960 646398
rect 592340 610718 592372 610954
rect 592608 610718 592692 610954
rect 592928 610718 592960 610954
rect 592340 610634 592960 610718
rect 592340 610398 592372 610634
rect 592608 610398 592692 610634
rect 592928 610398 592960 610634
rect 592340 574954 592960 610398
rect 592340 574718 592372 574954
rect 592608 574718 592692 574954
rect 592928 574718 592960 574954
rect 592340 574634 592960 574718
rect 592340 574398 592372 574634
rect 592608 574398 592692 574634
rect 592928 574398 592960 574634
rect 592340 538954 592960 574398
rect 592340 538718 592372 538954
rect 592608 538718 592692 538954
rect 592928 538718 592960 538954
rect 592340 538634 592960 538718
rect 592340 538398 592372 538634
rect 592608 538398 592692 538634
rect 592928 538398 592960 538634
rect 592340 502954 592960 538398
rect 592340 502718 592372 502954
rect 592608 502718 592692 502954
rect 592928 502718 592960 502954
rect 592340 502634 592960 502718
rect 592340 502398 592372 502634
rect 592608 502398 592692 502634
rect 592928 502398 592960 502634
rect 592340 466954 592960 502398
rect 592340 466718 592372 466954
rect 592608 466718 592692 466954
rect 592928 466718 592960 466954
rect 592340 466634 592960 466718
rect 592340 466398 592372 466634
rect 592608 466398 592692 466634
rect 592928 466398 592960 466634
rect 592340 430954 592960 466398
rect 592340 430718 592372 430954
rect 592608 430718 592692 430954
rect 592928 430718 592960 430954
rect 592340 430634 592960 430718
rect 592340 430398 592372 430634
rect 592608 430398 592692 430634
rect 592928 430398 592960 430634
rect 592340 394954 592960 430398
rect 592340 394718 592372 394954
rect 592608 394718 592692 394954
rect 592928 394718 592960 394954
rect 592340 394634 592960 394718
rect 592340 394398 592372 394634
rect 592608 394398 592692 394634
rect 592928 394398 592960 394634
rect 592340 358954 592960 394398
rect 592340 358718 592372 358954
rect 592608 358718 592692 358954
rect 592928 358718 592960 358954
rect 592340 358634 592960 358718
rect 592340 358398 592372 358634
rect 592608 358398 592692 358634
rect 592928 358398 592960 358634
rect 592340 322954 592960 358398
rect 592340 322718 592372 322954
rect 592608 322718 592692 322954
rect 592928 322718 592960 322954
rect 592340 322634 592960 322718
rect 592340 322398 592372 322634
rect 592608 322398 592692 322634
rect 592928 322398 592960 322634
rect 592340 286954 592960 322398
rect 592340 286718 592372 286954
rect 592608 286718 592692 286954
rect 592928 286718 592960 286954
rect 592340 286634 592960 286718
rect 592340 286398 592372 286634
rect 592608 286398 592692 286634
rect 592928 286398 592960 286634
rect 592340 250954 592960 286398
rect 592340 250718 592372 250954
rect 592608 250718 592692 250954
rect 592928 250718 592960 250954
rect 592340 250634 592960 250718
rect 592340 250398 592372 250634
rect 592608 250398 592692 250634
rect 592928 250398 592960 250634
rect 592340 214954 592960 250398
rect 592340 214718 592372 214954
rect 592608 214718 592692 214954
rect 592928 214718 592960 214954
rect 592340 214634 592960 214718
rect 592340 214398 592372 214634
rect 592608 214398 592692 214634
rect 592928 214398 592960 214634
rect 592340 178954 592960 214398
rect 592340 178718 592372 178954
rect 592608 178718 592692 178954
rect 592928 178718 592960 178954
rect 592340 178634 592960 178718
rect 592340 178398 592372 178634
rect 592608 178398 592692 178634
rect 592928 178398 592960 178634
rect 592340 142954 592960 178398
rect 592340 142718 592372 142954
rect 592608 142718 592692 142954
rect 592928 142718 592960 142954
rect 592340 142634 592960 142718
rect 592340 142398 592372 142634
rect 592608 142398 592692 142634
rect 592928 142398 592960 142634
rect 592340 106954 592960 142398
rect 592340 106718 592372 106954
rect 592608 106718 592692 106954
rect 592928 106718 592960 106954
rect 592340 106634 592960 106718
rect 592340 106398 592372 106634
rect 592608 106398 592692 106634
rect 592928 106398 592960 106634
rect 592340 70954 592960 106398
rect 592340 70718 592372 70954
rect 592608 70718 592692 70954
rect 592928 70718 592960 70954
rect 592340 70634 592960 70718
rect 592340 70398 592372 70634
rect 592608 70398 592692 70634
rect 592928 70398 592960 70634
rect 592340 34954 592960 70398
rect 592340 34718 592372 34954
rect 592608 34718 592692 34954
rect 592928 34718 592960 34954
rect 592340 34634 592960 34718
rect 592340 34398 592372 34634
rect 592608 34398 592692 34634
rect 592928 34398 592960 34634
rect 592340 -7376 592960 34398
rect 592340 -7612 592372 -7376
rect 592608 -7612 592692 -7376
rect 592928 -7612 592960 -7376
rect 592340 -7696 592960 -7612
rect 592340 -7932 592372 -7696
rect 592608 -7932 592692 -7696
rect 592928 -7932 592960 -7696
rect 592340 -7964 592960 -7932
<< via4 >>
rect -9004 711632 -8768 711868
rect -8684 711632 -8448 711868
rect -9004 711312 -8768 711548
rect -8684 711312 -8448 711548
rect -9004 682718 -8768 682954
rect -8684 682718 -8448 682954
rect -9004 682398 -8768 682634
rect -8684 682398 -8448 682634
rect -9004 646718 -8768 646954
rect -8684 646718 -8448 646954
rect -9004 646398 -8768 646634
rect -8684 646398 -8448 646634
rect -9004 610718 -8768 610954
rect -8684 610718 -8448 610954
rect -9004 610398 -8768 610634
rect -8684 610398 -8448 610634
rect -9004 574718 -8768 574954
rect -8684 574718 -8448 574954
rect -9004 574398 -8768 574634
rect -8684 574398 -8448 574634
rect -9004 538718 -8768 538954
rect -8684 538718 -8448 538954
rect -9004 538398 -8768 538634
rect -8684 538398 -8448 538634
rect -9004 502718 -8768 502954
rect -8684 502718 -8448 502954
rect -9004 502398 -8768 502634
rect -8684 502398 -8448 502634
rect -9004 466718 -8768 466954
rect -8684 466718 -8448 466954
rect -9004 466398 -8768 466634
rect -8684 466398 -8448 466634
rect -9004 430718 -8768 430954
rect -8684 430718 -8448 430954
rect -9004 430398 -8768 430634
rect -8684 430398 -8448 430634
rect -9004 394718 -8768 394954
rect -8684 394718 -8448 394954
rect -9004 394398 -8768 394634
rect -8684 394398 -8448 394634
rect -9004 358718 -8768 358954
rect -8684 358718 -8448 358954
rect -9004 358398 -8768 358634
rect -8684 358398 -8448 358634
rect -9004 322718 -8768 322954
rect -8684 322718 -8448 322954
rect -9004 322398 -8768 322634
rect -8684 322398 -8448 322634
rect -9004 286718 -8768 286954
rect -8684 286718 -8448 286954
rect -9004 286398 -8768 286634
rect -8684 286398 -8448 286634
rect -9004 250718 -8768 250954
rect -8684 250718 -8448 250954
rect -9004 250398 -8768 250634
rect -8684 250398 -8448 250634
rect -9004 214718 -8768 214954
rect -8684 214718 -8448 214954
rect -9004 214398 -8768 214634
rect -8684 214398 -8448 214634
rect -9004 178718 -8768 178954
rect -8684 178718 -8448 178954
rect -9004 178398 -8768 178634
rect -8684 178398 -8448 178634
rect -9004 142718 -8768 142954
rect -8684 142718 -8448 142954
rect -9004 142398 -8768 142634
rect -8684 142398 -8448 142634
rect -9004 106718 -8768 106954
rect -8684 106718 -8448 106954
rect -9004 106398 -8768 106634
rect -8684 106398 -8448 106634
rect -9004 70718 -8768 70954
rect -8684 70718 -8448 70954
rect -9004 70398 -8768 70634
rect -8684 70398 -8448 70634
rect -9004 34718 -8768 34954
rect -8684 34718 -8448 34954
rect -9004 34398 -8768 34634
rect -8684 34398 -8448 34634
rect -8044 710672 -7808 710908
rect -7724 710672 -7488 710908
rect -8044 710352 -7808 710588
rect -7724 710352 -7488 710588
rect -8044 678218 -7808 678454
rect -7724 678218 -7488 678454
rect -8044 677898 -7808 678134
rect -7724 677898 -7488 678134
rect -8044 642218 -7808 642454
rect -7724 642218 -7488 642454
rect -8044 641898 -7808 642134
rect -7724 641898 -7488 642134
rect -8044 606218 -7808 606454
rect -7724 606218 -7488 606454
rect -8044 605898 -7808 606134
rect -7724 605898 -7488 606134
rect -8044 570218 -7808 570454
rect -7724 570218 -7488 570454
rect -8044 569898 -7808 570134
rect -7724 569898 -7488 570134
rect -8044 534218 -7808 534454
rect -7724 534218 -7488 534454
rect -8044 533898 -7808 534134
rect -7724 533898 -7488 534134
rect -8044 498218 -7808 498454
rect -7724 498218 -7488 498454
rect -8044 497898 -7808 498134
rect -7724 497898 -7488 498134
rect -8044 462218 -7808 462454
rect -7724 462218 -7488 462454
rect -8044 461898 -7808 462134
rect -7724 461898 -7488 462134
rect -8044 426218 -7808 426454
rect -7724 426218 -7488 426454
rect -8044 425898 -7808 426134
rect -7724 425898 -7488 426134
rect -8044 390218 -7808 390454
rect -7724 390218 -7488 390454
rect -8044 389898 -7808 390134
rect -7724 389898 -7488 390134
rect -8044 354218 -7808 354454
rect -7724 354218 -7488 354454
rect -8044 353898 -7808 354134
rect -7724 353898 -7488 354134
rect -8044 318218 -7808 318454
rect -7724 318218 -7488 318454
rect -8044 317898 -7808 318134
rect -7724 317898 -7488 318134
rect -8044 282218 -7808 282454
rect -7724 282218 -7488 282454
rect -8044 281898 -7808 282134
rect -7724 281898 -7488 282134
rect -8044 246218 -7808 246454
rect -7724 246218 -7488 246454
rect -8044 245898 -7808 246134
rect -7724 245898 -7488 246134
rect -8044 210218 -7808 210454
rect -7724 210218 -7488 210454
rect -8044 209898 -7808 210134
rect -7724 209898 -7488 210134
rect -8044 174218 -7808 174454
rect -7724 174218 -7488 174454
rect -8044 173898 -7808 174134
rect -7724 173898 -7488 174134
rect -8044 138218 -7808 138454
rect -7724 138218 -7488 138454
rect -8044 137898 -7808 138134
rect -7724 137898 -7488 138134
rect -8044 102218 -7808 102454
rect -7724 102218 -7488 102454
rect -8044 101898 -7808 102134
rect -7724 101898 -7488 102134
rect -8044 66218 -7808 66454
rect -7724 66218 -7488 66454
rect -8044 65898 -7808 66134
rect -7724 65898 -7488 66134
rect -8044 30218 -7808 30454
rect -7724 30218 -7488 30454
rect -8044 29898 -7808 30134
rect -7724 29898 -7488 30134
rect -7084 709712 -6848 709948
rect -6764 709712 -6528 709948
rect -7084 709392 -6848 709628
rect -6764 709392 -6528 709628
rect -7084 673718 -6848 673954
rect -6764 673718 -6528 673954
rect -7084 673398 -6848 673634
rect -6764 673398 -6528 673634
rect -7084 637718 -6848 637954
rect -6764 637718 -6528 637954
rect -7084 637398 -6848 637634
rect -6764 637398 -6528 637634
rect -7084 601718 -6848 601954
rect -6764 601718 -6528 601954
rect -7084 601398 -6848 601634
rect -6764 601398 -6528 601634
rect -7084 565718 -6848 565954
rect -6764 565718 -6528 565954
rect -7084 565398 -6848 565634
rect -6764 565398 -6528 565634
rect -7084 529718 -6848 529954
rect -6764 529718 -6528 529954
rect -7084 529398 -6848 529634
rect -6764 529398 -6528 529634
rect -7084 493718 -6848 493954
rect -6764 493718 -6528 493954
rect -7084 493398 -6848 493634
rect -6764 493398 -6528 493634
rect -7084 457718 -6848 457954
rect -6764 457718 -6528 457954
rect -7084 457398 -6848 457634
rect -6764 457398 -6528 457634
rect -7084 421718 -6848 421954
rect -6764 421718 -6528 421954
rect -7084 421398 -6848 421634
rect -6764 421398 -6528 421634
rect -7084 385718 -6848 385954
rect -6764 385718 -6528 385954
rect -7084 385398 -6848 385634
rect -6764 385398 -6528 385634
rect -7084 349718 -6848 349954
rect -6764 349718 -6528 349954
rect -7084 349398 -6848 349634
rect -6764 349398 -6528 349634
rect -7084 313718 -6848 313954
rect -6764 313718 -6528 313954
rect -7084 313398 -6848 313634
rect -6764 313398 -6528 313634
rect -7084 277718 -6848 277954
rect -6764 277718 -6528 277954
rect -7084 277398 -6848 277634
rect -6764 277398 -6528 277634
rect -7084 241718 -6848 241954
rect -6764 241718 -6528 241954
rect -7084 241398 -6848 241634
rect -6764 241398 -6528 241634
rect -7084 205718 -6848 205954
rect -6764 205718 -6528 205954
rect -7084 205398 -6848 205634
rect -6764 205398 -6528 205634
rect -7084 169718 -6848 169954
rect -6764 169718 -6528 169954
rect -7084 169398 -6848 169634
rect -6764 169398 -6528 169634
rect -7084 133718 -6848 133954
rect -6764 133718 -6528 133954
rect -7084 133398 -6848 133634
rect -6764 133398 -6528 133634
rect -7084 97718 -6848 97954
rect -6764 97718 -6528 97954
rect -7084 97398 -6848 97634
rect -6764 97398 -6528 97634
rect -7084 61718 -6848 61954
rect -6764 61718 -6528 61954
rect -7084 61398 -6848 61634
rect -6764 61398 -6528 61634
rect -7084 25718 -6848 25954
rect -6764 25718 -6528 25954
rect -7084 25398 -6848 25634
rect -6764 25398 -6528 25634
rect -6124 708752 -5888 708988
rect -5804 708752 -5568 708988
rect -6124 708432 -5888 708668
rect -5804 708432 -5568 708668
rect -6124 669218 -5888 669454
rect -5804 669218 -5568 669454
rect -6124 668898 -5888 669134
rect -5804 668898 -5568 669134
rect -6124 633218 -5888 633454
rect -5804 633218 -5568 633454
rect -6124 632898 -5888 633134
rect -5804 632898 -5568 633134
rect -6124 597218 -5888 597454
rect -5804 597218 -5568 597454
rect -6124 596898 -5888 597134
rect -5804 596898 -5568 597134
rect -6124 561218 -5888 561454
rect -5804 561218 -5568 561454
rect -6124 560898 -5888 561134
rect -5804 560898 -5568 561134
rect -6124 525218 -5888 525454
rect -5804 525218 -5568 525454
rect -6124 524898 -5888 525134
rect -5804 524898 -5568 525134
rect -6124 489218 -5888 489454
rect -5804 489218 -5568 489454
rect -6124 488898 -5888 489134
rect -5804 488898 -5568 489134
rect -6124 453218 -5888 453454
rect -5804 453218 -5568 453454
rect -6124 452898 -5888 453134
rect -5804 452898 -5568 453134
rect -6124 417218 -5888 417454
rect -5804 417218 -5568 417454
rect -6124 416898 -5888 417134
rect -5804 416898 -5568 417134
rect -6124 381218 -5888 381454
rect -5804 381218 -5568 381454
rect -6124 380898 -5888 381134
rect -5804 380898 -5568 381134
rect -6124 345218 -5888 345454
rect -5804 345218 -5568 345454
rect -6124 344898 -5888 345134
rect -5804 344898 -5568 345134
rect -6124 309218 -5888 309454
rect -5804 309218 -5568 309454
rect -6124 308898 -5888 309134
rect -5804 308898 -5568 309134
rect -6124 273218 -5888 273454
rect -5804 273218 -5568 273454
rect -6124 272898 -5888 273134
rect -5804 272898 -5568 273134
rect -6124 237218 -5888 237454
rect -5804 237218 -5568 237454
rect -6124 236898 -5888 237134
rect -5804 236898 -5568 237134
rect -6124 201218 -5888 201454
rect -5804 201218 -5568 201454
rect -6124 200898 -5888 201134
rect -5804 200898 -5568 201134
rect -6124 165218 -5888 165454
rect -5804 165218 -5568 165454
rect -6124 164898 -5888 165134
rect -5804 164898 -5568 165134
rect -6124 129218 -5888 129454
rect -5804 129218 -5568 129454
rect -6124 128898 -5888 129134
rect -5804 128898 -5568 129134
rect -6124 93218 -5888 93454
rect -5804 93218 -5568 93454
rect -6124 92898 -5888 93134
rect -5804 92898 -5568 93134
rect -6124 57218 -5888 57454
rect -5804 57218 -5568 57454
rect -6124 56898 -5888 57134
rect -5804 56898 -5568 57134
rect -6124 21218 -5888 21454
rect -5804 21218 -5568 21454
rect -6124 20898 -5888 21134
rect -5804 20898 -5568 21134
rect -5164 707792 -4928 708028
rect -4844 707792 -4608 708028
rect -5164 707472 -4928 707708
rect -4844 707472 -4608 707708
rect -5164 700718 -4928 700954
rect -4844 700718 -4608 700954
rect -5164 700398 -4928 700634
rect -4844 700398 -4608 700634
rect -5164 664718 -4928 664954
rect -4844 664718 -4608 664954
rect -5164 664398 -4928 664634
rect -4844 664398 -4608 664634
rect -5164 628718 -4928 628954
rect -4844 628718 -4608 628954
rect -5164 628398 -4928 628634
rect -4844 628398 -4608 628634
rect -5164 592718 -4928 592954
rect -4844 592718 -4608 592954
rect -5164 592398 -4928 592634
rect -4844 592398 -4608 592634
rect -5164 556718 -4928 556954
rect -4844 556718 -4608 556954
rect -5164 556398 -4928 556634
rect -4844 556398 -4608 556634
rect -5164 520718 -4928 520954
rect -4844 520718 -4608 520954
rect -5164 520398 -4928 520634
rect -4844 520398 -4608 520634
rect -5164 484718 -4928 484954
rect -4844 484718 -4608 484954
rect -5164 484398 -4928 484634
rect -4844 484398 -4608 484634
rect -5164 448718 -4928 448954
rect -4844 448718 -4608 448954
rect -5164 448398 -4928 448634
rect -4844 448398 -4608 448634
rect -5164 412718 -4928 412954
rect -4844 412718 -4608 412954
rect -5164 412398 -4928 412634
rect -4844 412398 -4608 412634
rect -5164 376718 -4928 376954
rect -4844 376718 -4608 376954
rect -5164 376398 -4928 376634
rect -4844 376398 -4608 376634
rect -5164 340718 -4928 340954
rect -4844 340718 -4608 340954
rect -5164 340398 -4928 340634
rect -4844 340398 -4608 340634
rect -5164 304718 -4928 304954
rect -4844 304718 -4608 304954
rect -5164 304398 -4928 304634
rect -4844 304398 -4608 304634
rect -5164 268718 -4928 268954
rect -4844 268718 -4608 268954
rect -5164 268398 -4928 268634
rect -4844 268398 -4608 268634
rect -5164 232718 -4928 232954
rect -4844 232718 -4608 232954
rect -5164 232398 -4928 232634
rect -4844 232398 -4608 232634
rect -5164 196718 -4928 196954
rect -4844 196718 -4608 196954
rect -5164 196398 -4928 196634
rect -4844 196398 -4608 196634
rect -5164 160718 -4928 160954
rect -4844 160718 -4608 160954
rect -5164 160398 -4928 160634
rect -4844 160398 -4608 160634
rect -5164 124718 -4928 124954
rect -4844 124718 -4608 124954
rect -5164 124398 -4928 124634
rect -4844 124398 -4608 124634
rect -5164 88718 -4928 88954
rect -4844 88718 -4608 88954
rect -5164 88398 -4928 88634
rect -4844 88398 -4608 88634
rect -5164 52718 -4928 52954
rect -4844 52718 -4608 52954
rect -5164 52398 -4928 52634
rect -4844 52398 -4608 52634
rect -5164 16718 -4928 16954
rect -4844 16718 -4608 16954
rect -5164 16398 -4928 16634
rect -4844 16398 -4608 16634
rect -4204 706832 -3968 707068
rect -3884 706832 -3648 707068
rect -4204 706512 -3968 706748
rect -3884 706512 -3648 706748
rect -4204 696218 -3968 696454
rect -3884 696218 -3648 696454
rect -4204 695898 -3968 696134
rect -3884 695898 -3648 696134
rect -4204 660218 -3968 660454
rect -3884 660218 -3648 660454
rect -4204 659898 -3968 660134
rect -3884 659898 -3648 660134
rect -4204 624218 -3968 624454
rect -3884 624218 -3648 624454
rect -4204 623898 -3968 624134
rect -3884 623898 -3648 624134
rect -4204 588218 -3968 588454
rect -3884 588218 -3648 588454
rect -4204 587898 -3968 588134
rect -3884 587898 -3648 588134
rect -4204 552218 -3968 552454
rect -3884 552218 -3648 552454
rect -4204 551898 -3968 552134
rect -3884 551898 -3648 552134
rect -4204 516218 -3968 516454
rect -3884 516218 -3648 516454
rect -4204 515898 -3968 516134
rect -3884 515898 -3648 516134
rect -4204 480218 -3968 480454
rect -3884 480218 -3648 480454
rect -4204 479898 -3968 480134
rect -3884 479898 -3648 480134
rect -4204 444218 -3968 444454
rect -3884 444218 -3648 444454
rect -4204 443898 -3968 444134
rect -3884 443898 -3648 444134
rect -4204 408218 -3968 408454
rect -3884 408218 -3648 408454
rect -4204 407898 -3968 408134
rect -3884 407898 -3648 408134
rect -4204 372218 -3968 372454
rect -3884 372218 -3648 372454
rect -4204 371898 -3968 372134
rect -3884 371898 -3648 372134
rect -4204 336218 -3968 336454
rect -3884 336218 -3648 336454
rect -4204 335898 -3968 336134
rect -3884 335898 -3648 336134
rect -4204 300218 -3968 300454
rect -3884 300218 -3648 300454
rect -4204 299898 -3968 300134
rect -3884 299898 -3648 300134
rect -4204 264218 -3968 264454
rect -3884 264218 -3648 264454
rect -4204 263898 -3968 264134
rect -3884 263898 -3648 264134
rect -4204 228218 -3968 228454
rect -3884 228218 -3648 228454
rect -4204 227898 -3968 228134
rect -3884 227898 -3648 228134
rect -4204 192218 -3968 192454
rect -3884 192218 -3648 192454
rect -4204 191898 -3968 192134
rect -3884 191898 -3648 192134
rect -4204 156218 -3968 156454
rect -3884 156218 -3648 156454
rect -4204 155898 -3968 156134
rect -3884 155898 -3648 156134
rect -4204 120218 -3968 120454
rect -3884 120218 -3648 120454
rect -4204 119898 -3968 120134
rect -3884 119898 -3648 120134
rect -4204 84218 -3968 84454
rect -3884 84218 -3648 84454
rect -4204 83898 -3968 84134
rect -3884 83898 -3648 84134
rect -4204 48218 -3968 48454
rect -3884 48218 -3648 48454
rect -4204 47898 -3968 48134
rect -3884 47898 -3648 48134
rect -4204 12218 -3968 12454
rect -3884 12218 -3648 12454
rect -4204 11898 -3968 12134
rect -3884 11898 -3648 12134
rect -3244 705872 -3008 706108
rect -2924 705872 -2688 706108
rect -3244 705552 -3008 705788
rect -2924 705552 -2688 705788
rect -3244 691718 -3008 691954
rect -2924 691718 -2688 691954
rect -3244 691398 -3008 691634
rect -2924 691398 -2688 691634
rect -3244 655718 -3008 655954
rect -2924 655718 -2688 655954
rect -3244 655398 -3008 655634
rect -2924 655398 -2688 655634
rect -3244 619718 -3008 619954
rect -2924 619718 -2688 619954
rect -3244 619398 -3008 619634
rect -2924 619398 -2688 619634
rect -3244 583718 -3008 583954
rect -2924 583718 -2688 583954
rect -3244 583398 -3008 583634
rect -2924 583398 -2688 583634
rect -3244 547718 -3008 547954
rect -2924 547718 -2688 547954
rect -3244 547398 -3008 547634
rect -2924 547398 -2688 547634
rect -3244 511718 -3008 511954
rect -2924 511718 -2688 511954
rect -3244 511398 -3008 511634
rect -2924 511398 -2688 511634
rect -3244 475718 -3008 475954
rect -2924 475718 -2688 475954
rect -3244 475398 -3008 475634
rect -2924 475398 -2688 475634
rect -3244 439718 -3008 439954
rect -2924 439718 -2688 439954
rect -3244 439398 -3008 439634
rect -2924 439398 -2688 439634
rect -3244 403718 -3008 403954
rect -2924 403718 -2688 403954
rect -3244 403398 -3008 403634
rect -2924 403398 -2688 403634
rect -3244 367718 -3008 367954
rect -2924 367718 -2688 367954
rect -3244 367398 -3008 367634
rect -2924 367398 -2688 367634
rect -3244 331718 -3008 331954
rect -2924 331718 -2688 331954
rect -3244 331398 -3008 331634
rect -2924 331398 -2688 331634
rect -3244 295718 -3008 295954
rect -2924 295718 -2688 295954
rect -3244 295398 -3008 295634
rect -2924 295398 -2688 295634
rect -3244 259718 -3008 259954
rect -2924 259718 -2688 259954
rect -3244 259398 -3008 259634
rect -2924 259398 -2688 259634
rect -3244 223718 -3008 223954
rect -2924 223718 -2688 223954
rect -3244 223398 -3008 223634
rect -2924 223398 -2688 223634
rect -3244 187718 -3008 187954
rect -2924 187718 -2688 187954
rect -3244 187398 -3008 187634
rect -2924 187398 -2688 187634
rect -3244 151718 -3008 151954
rect -2924 151718 -2688 151954
rect -3244 151398 -3008 151634
rect -2924 151398 -2688 151634
rect -3244 115718 -3008 115954
rect -2924 115718 -2688 115954
rect -3244 115398 -3008 115634
rect -2924 115398 -2688 115634
rect -3244 79718 -3008 79954
rect -2924 79718 -2688 79954
rect -3244 79398 -3008 79634
rect -2924 79398 -2688 79634
rect -3244 43718 -3008 43954
rect -2924 43718 -2688 43954
rect -3244 43398 -3008 43634
rect -2924 43398 -2688 43634
rect -3244 7718 -3008 7954
rect -2924 7718 -2688 7954
rect -3244 7398 -3008 7634
rect -2924 7398 -2688 7634
rect -2284 704912 -2048 705148
rect -1964 704912 -1728 705148
rect -2284 704592 -2048 704828
rect -1964 704592 -1728 704828
rect -2284 687218 -2048 687454
rect -1964 687218 -1728 687454
rect -2284 686898 -2048 687134
rect -1964 686898 -1728 687134
rect -2284 651218 -2048 651454
rect -1964 651218 -1728 651454
rect -2284 650898 -2048 651134
rect -1964 650898 -1728 651134
rect -2284 615218 -2048 615454
rect -1964 615218 -1728 615454
rect -2284 614898 -2048 615134
rect -1964 614898 -1728 615134
rect -2284 579218 -2048 579454
rect -1964 579218 -1728 579454
rect -2284 578898 -2048 579134
rect -1964 578898 -1728 579134
rect -2284 543218 -2048 543454
rect -1964 543218 -1728 543454
rect -2284 542898 -2048 543134
rect -1964 542898 -1728 543134
rect -2284 507218 -2048 507454
rect -1964 507218 -1728 507454
rect -2284 506898 -2048 507134
rect -1964 506898 -1728 507134
rect -2284 471218 -2048 471454
rect -1964 471218 -1728 471454
rect -2284 470898 -2048 471134
rect -1964 470898 -1728 471134
rect -2284 435218 -2048 435454
rect -1964 435218 -1728 435454
rect -2284 434898 -2048 435134
rect -1964 434898 -1728 435134
rect -2284 399218 -2048 399454
rect -1964 399218 -1728 399454
rect -2284 398898 -2048 399134
rect -1964 398898 -1728 399134
rect -2284 363218 -2048 363454
rect -1964 363218 -1728 363454
rect -2284 362898 -2048 363134
rect -1964 362898 -1728 363134
rect -2284 327218 -2048 327454
rect -1964 327218 -1728 327454
rect -2284 326898 -2048 327134
rect -1964 326898 -1728 327134
rect -2284 291218 -2048 291454
rect -1964 291218 -1728 291454
rect -2284 290898 -2048 291134
rect -1964 290898 -1728 291134
rect -2284 255218 -2048 255454
rect -1964 255218 -1728 255454
rect -2284 254898 -2048 255134
rect -1964 254898 -1728 255134
rect -2284 219218 -2048 219454
rect -1964 219218 -1728 219454
rect -2284 218898 -2048 219134
rect -1964 218898 -1728 219134
rect -2284 183218 -2048 183454
rect -1964 183218 -1728 183454
rect -2284 182898 -2048 183134
rect -1964 182898 -1728 183134
rect -2284 147218 -2048 147454
rect -1964 147218 -1728 147454
rect -2284 146898 -2048 147134
rect -1964 146898 -1728 147134
rect -2284 111218 -2048 111454
rect -1964 111218 -1728 111454
rect -2284 110898 -2048 111134
rect -1964 110898 -1728 111134
rect -2284 75218 -2048 75454
rect -1964 75218 -1728 75454
rect -2284 74898 -2048 75134
rect -1964 74898 -1728 75134
rect -2284 39218 -2048 39454
rect -1964 39218 -1728 39454
rect -2284 38898 -2048 39134
rect -1964 38898 -1728 39134
rect -2284 3218 -2048 3454
rect -1964 3218 -1728 3454
rect -2284 2898 -2048 3134
rect -1964 2898 -1728 3134
rect -2284 -892 -2048 -656
rect -1964 -892 -1728 -656
rect -2284 -1212 -2048 -976
rect -1964 -1212 -1728 -976
rect 1826 704912 2062 705148
rect 2146 704912 2382 705148
rect 1826 704592 2062 704828
rect 2146 704592 2382 704828
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -892 2062 -656
rect 2146 -892 2382 -656
rect 1826 -1212 2062 -976
rect 2146 -1212 2382 -976
rect -3244 -1852 -3008 -1616
rect -2924 -1852 -2688 -1616
rect -3244 -2172 -3008 -1936
rect -2924 -2172 -2688 -1936
rect -4204 -2812 -3968 -2576
rect -3884 -2812 -3648 -2576
rect -4204 -3132 -3968 -2896
rect -3884 -3132 -3648 -2896
rect -5164 -3772 -4928 -3536
rect -4844 -3772 -4608 -3536
rect -5164 -4092 -4928 -3856
rect -4844 -4092 -4608 -3856
rect -6124 -4732 -5888 -4496
rect -5804 -4732 -5568 -4496
rect -6124 -5052 -5888 -4816
rect -5804 -5052 -5568 -4816
rect -7084 -5692 -6848 -5456
rect -6764 -5692 -6528 -5456
rect -7084 -6012 -6848 -5776
rect -6764 -6012 -6528 -5776
rect -8044 -6652 -7808 -6416
rect -7724 -6652 -7488 -6416
rect -8044 -6972 -7808 -6736
rect -7724 -6972 -7488 -6736
rect -9004 -7612 -8768 -7376
rect -8684 -7612 -8448 -7376
rect -9004 -7932 -8768 -7696
rect -8684 -7932 -8448 -7696
rect 6326 705872 6562 706108
rect 6646 705872 6882 706108
rect 6326 705552 6562 705788
rect 6646 705552 6882 705788
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1852 6562 -1616
rect 6646 -1852 6882 -1616
rect 6326 -2172 6562 -1936
rect 6646 -2172 6882 -1936
rect 10826 706832 11062 707068
rect 11146 706832 11382 707068
rect 10826 706512 11062 706748
rect 11146 706512 11382 706748
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2812 11062 -2576
rect 11146 -2812 11382 -2576
rect 10826 -3132 11062 -2896
rect 11146 -3132 11382 -2896
rect 15326 707792 15562 708028
rect 15646 707792 15882 708028
rect 15326 707472 15562 707708
rect 15646 707472 15882 707708
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3772 15562 -3536
rect 15646 -3772 15882 -3536
rect 15326 -4092 15562 -3856
rect 15646 -4092 15882 -3856
rect 19826 708752 20062 708988
rect 20146 708752 20382 708988
rect 19826 708432 20062 708668
rect 20146 708432 20382 708668
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4732 20062 -4496
rect 20146 -4732 20382 -4496
rect 19826 -5052 20062 -4816
rect 20146 -5052 20382 -4816
rect 24326 709712 24562 709948
rect 24646 709712 24882 709948
rect 24326 709392 24562 709628
rect 24646 709392 24882 709628
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5692 24562 -5456
rect 24646 -5692 24882 -5456
rect 24326 -6012 24562 -5776
rect 24646 -6012 24882 -5776
rect 28826 710672 29062 710908
rect 29146 710672 29382 710908
rect 28826 710352 29062 710588
rect 29146 710352 29382 710588
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6652 29062 -6416
rect 29146 -6652 29382 -6416
rect 28826 -6972 29062 -6736
rect 29146 -6972 29382 -6736
rect 33326 711632 33562 711868
rect 33646 711632 33882 711868
rect 33326 711312 33562 711548
rect 33646 711312 33882 711548
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7612 33562 -7376
rect 33646 -7612 33882 -7376
rect 33326 -7932 33562 -7696
rect 33646 -7932 33882 -7696
rect 37826 704912 38062 705148
rect 38146 704912 38382 705148
rect 37826 704592 38062 704828
rect 38146 704592 38382 704828
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -892 38062 -656
rect 38146 -892 38382 -656
rect 37826 -1212 38062 -976
rect 38146 -1212 38382 -976
rect 42326 705872 42562 706108
rect 42646 705872 42882 706108
rect 42326 705552 42562 705788
rect 42646 705552 42882 705788
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1852 42562 -1616
rect 42646 -1852 42882 -1616
rect 42326 -2172 42562 -1936
rect 42646 -2172 42882 -1936
rect 46826 706832 47062 707068
rect 47146 706832 47382 707068
rect 46826 706512 47062 706748
rect 47146 706512 47382 706748
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2812 47062 -2576
rect 47146 -2812 47382 -2576
rect 46826 -3132 47062 -2896
rect 47146 -3132 47382 -2896
rect 51326 707792 51562 708028
rect 51646 707792 51882 708028
rect 51326 707472 51562 707708
rect 51646 707472 51882 707708
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3772 51562 -3536
rect 51646 -3772 51882 -3536
rect 51326 -4092 51562 -3856
rect 51646 -4092 51882 -3856
rect 55826 708752 56062 708988
rect 56146 708752 56382 708988
rect 55826 708432 56062 708668
rect 56146 708432 56382 708668
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4732 56062 -4496
rect 56146 -4732 56382 -4496
rect 55826 -5052 56062 -4816
rect 56146 -5052 56382 -4816
rect 60326 709712 60562 709948
rect 60646 709712 60882 709948
rect 60326 709392 60562 709628
rect 60646 709392 60882 709628
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5692 60562 -5456
rect 60646 -5692 60882 -5456
rect 60326 -6012 60562 -5776
rect 60646 -6012 60882 -5776
rect 64826 710672 65062 710908
rect 65146 710672 65382 710908
rect 64826 710352 65062 710588
rect 65146 710352 65382 710588
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6652 65062 -6416
rect 65146 -6652 65382 -6416
rect 64826 -6972 65062 -6736
rect 65146 -6972 65382 -6736
rect 69326 711632 69562 711868
rect 69646 711632 69882 711868
rect 69326 711312 69562 711548
rect 69646 711312 69882 711548
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7612 69562 -7376
rect 69646 -7612 69882 -7376
rect 69326 -7932 69562 -7696
rect 69646 -7932 69882 -7696
rect 73826 704912 74062 705148
rect 74146 704912 74382 705148
rect 73826 704592 74062 704828
rect 74146 704592 74382 704828
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -892 74062 -656
rect 74146 -892 74382 -656
rect 73826 -1212 74062 -976
rect 74146 -1212 74382 -976
rect 78326 705872 78562 706108
rect 78646 705872 78882 706108
rect 78326 705552 78562 705788
rect 78646 705552 78882 705788
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1852 78562 -1616
rect 78646 -1852 78882 -1616
rect 78326 -2172 78562 -1936
rect 78646 -2172 78882 -1936
rect 82826 706832 83062 707068
rect 83146 706832 83382 707068
rect 82826 706512 83062 706748
rect 83146 706512 83382 706748
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2812 83062 -2576
rect 83146 -2812 83382 -2576
rect 82826 -3132 83062 -2896
rect 83146 -3132 83382 -2896
rect 87326 707792 87562 708028
rect 87646 707792 87882 708028
rect 87326 707472 87562 707708
rect 87646 707472 87882 707708
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3772 87562 -3536
rect 87646 -3772 87882 -3536
rect 87326 -4092 87562 -3856
rect 87646 -4092 87882 -3856
rect 91826 708752 92062 708988
rect 92146 708752 92382 708988
rect 91826 708432 92062 708668
rect 92146 708432 92382 708668
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4732 92062 -4496
rect 92146 -4732 92382 -4496
rect 91826 -5052 92062 -4816
rect 92146 -5052 92382 -4816
rect 96326 709712 96562 709948
rect 96646 709712 96882 709948
rect 96326 709392 96562 709628
rect 96646 709392 96882 709628
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 100826 710672 101062 710908
rect 101146 710672 101382 710908
rect 100826 710352 101062 710588
rect 101146 710352 101382 710588
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 105326 711632 105562 711868
rect 105646 711632 105882 711868
rect 105326 711312 105562 711548
rect 105646 711312 105882 711548
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 109826 704912 110062 705148
rect 110146 704912 110382 705148
rect 109826 704592 110062 704828
rect 110146 704592 110382 704828
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 114326 705872 114562 706108
rect 114646 705872 114882 706108
rect 114326 705552 114562 705788
rect 114646 705552 114882 705788
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 118826 706832 119062 707068
rect 119146 706832 119382 707068
rect 118826 706512 119062 706748
rect 119146 706512 119382 706748
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 123326 707792 123562 708028
rect 123646 707792 123882 708028
rect 123326 707472 123562 707708
rect 123646 707472 123882 707708
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 127826 708752 128062 708988
rect 128146 708752 128382 708988
rect 127826 708432 128062 708668
rect 128146 708432 128382 708668
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 132326 709712 132562 709948
rect 132646 709712 132882 709948
rect 132326 709392 132562 709628
rect 132646 709392 132882 709628
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 136826 710672 137062 710908
rect 137146 710672 137382 710908
rect 136826 710352 137062 710588
rect 137146 710352 137382 710588
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 141326 711632 141562 711868
rect 141646 711632 141882 711868
rect 141326 711312 141562 711548
rect 141646 711312 141882 711548
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 145826 704912 146062 705148
rect 146146 704912 146382 705148
rect 145826 704592 146062 704828
rect 146146 704592 146382 704828
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 150326 705872 150562 706108
rect 150646 705872 150882 706108
rect 150326 705552 150562 705788
rect 150646 705552 150882 705788
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 154826 706832 155062 707068
rect 155146 706832 155382 707068
rect 154826 706512 155062 706748
rect 155146 706512 155382 706748
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 159326 707792 159562 708028
rect 159646 707792 159882 708028
rect 159326 707472 159562 707708
rect 159646 707472 159882 707708
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 163826 708752 164062 708988
rect 164146 708752 164382 708988
rect 163826 708432 164062 708668
rect 164146 708432 164382 708668
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 168326 709712 168562 709948
rect 168646 709712 168882 709948
rect 168326 709392 168562 709628
rect 168646 709392 168882 709628
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 172826 710672 173062 710908
rect 173146 710672 173382 710908
rect 172826 710352 173062 710588
rect 173146 710352 173382 710588
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 119610 367718 119846 367954
rect 119610 367398 119846 367634
rect 150330 367718 150566 367954
rect 150330 367398 150566 367634
rect 104250 363218 104486 363454
rect 104250 362898 104486 363134
rect 134970 363218 135206 363454
rect 134970 362898 135206 363134
rect 165690 363218 165926 363454
rect 165690 362898 165926 363134
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 119610 331718 119846 331954
rect 119610 331398 119846 331634
rect 150330 331718 150566 331954
rect 150330 331398 150566 331634
rect 104250 327218 104486 327454
rect 104250 326898 104486 327134
rect 134970 327218 135206 327454
rect 134970 326898 135206 327134
rect 165690 327218 165926 327454
rect 165690 326898 165926 327134
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 96326 241718 96562 241954
rect 96646 241718 96882 241954
rect 96326 241398 96562 241634
rect 96646 241398 96882 241634
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5692 96562 -5456
rect 96646 -5692 96882 -5456
rect 96326 -6012 96562 -5776
rect 96646 -6012 96882 -5776
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 100826 246218 101062 246454
rect 101146 246218 101382 246454
rect 100826 245898 101062 246134
rect 101146 245898 101382 246134
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6652 101062 -6416
rect 101146 -6652 101382 -6416
rect 100826 -6972 101062 -6736
rect 101146 -6972 101382 -6736
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7612 105562 -7376
rect 105646 -7612 105882 -7376
rect 105326 -7932 105562 -7696
rect 105646 -7932 105882 -7696
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -892 110062 -656
rect 110146 -892 110382 -656
rect 109826 -1212 110062 -976
rect 110146 -1212 110382 -976
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1852 114562 -1616
rect 114646 -1852 114882 -1616
rect 114326 -2172 114562 -1936
rect 114646 -2172 114882 -1936
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 118826 228218 119062 228454
rect 119146 228218 119382 228454
rect 118826 227898 119062 228134
rect 119146 227898 119382 228134
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 118826 120218 119062 120454
rect 119146 120218 119382 120454
rect 118826 119898 119062 120134
rect 119146 119898 119382 120134
rect 118826 84218 119062 84454
rect 119146 84218 119382 84454
rect 118826 83898 119062 84134
rect 119146 83898 119382 84134
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2812 119062 -2576
rect 119146 -2812 119382 -2576
rect 118826 -3132 119062 -2896
rect 119146 -3132 119382 -2896
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 123326 232718 123562 232954
rect 123646 232718 123882 232954
rect 123326 232398 123562 232634
rect 123646 232398 123882 232634
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 123326 124718 123562 124954
rect 123646 124718 123882 124954
rect 123326 124398 123562 124634
rect 123646 124398 123882 124634
rect 123326 88718 123562 88954
rect 123646 88718 123882 88954
rect 123326 88398 123562 88634
rect 123646 88398 123882 88634
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3772 123562 -3536
rect 123646 -3772 123882 -3536
rect 123326 -4092 123562 -3856
rect 123646 -4092 123882 -3856
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4732 128062 -4496
rect 128146 -4732 128382 -4496
rect 127826 -5052 128062 -4816
rect 128146 -5052 128382 -4816
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 132326 241718 132562 241954
rect 132646 241718 132882 241954
rect 132326 241398 132562 241634
rect 132646 241398 132882 241634
rect 132326 205718 132562 205954
rect 132646 205718 132882 205954
rect 132326 205398 132562 205634
rect 132646 205398 132882 205634
rect 132326 169718 132562 169954
rect 132646 169718 132882 169954
rect 132326 169398 132562 169634
rect 132646 169398 132882 169634
rect 132326 133718 132562 133954
rect 132646 133718 132882 133954
rect 132326 133398 132562 133634
rect 132646 133398 132882 133634
rect 132326 97718 132562 97954
rect 132646 97718 132882 97954
rect 132326 97398 132562 97634
rect 132646 97398 132882 97634
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5692 132562 -5456
rect 132646 -5692 132882 -5456
rect 132326 -6012 132562 -5776
rect 132646 -6012 132882 -5776
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 136826 246218 137062 246454
rect 137146 246218 137382 246454
rect 136826 245898 137062 246134
rect 137146 245898 137382 246134
rect 136826 210218 137062 210454
rect 137146 210218 137382 210454
rect 136826 209898 137062 210134
rect 137146 209898 137382 210134
rect 136826 174218 137062 174454
rect 137146 174218 137382 174454
rect 136826 173898 137062 174134
rect 137146 173898 137382 174134
rect 136826 138218 137062 138454
rect 137146 138218 137382 138454
rect 136826 137898 137062 138134
rect 137146 137898 137382 138134
rect 136826 102218 137062 102454
rect 137146 102218 137382 102454
rect 136826 101898 137062 102134
rect 137146 101898 137382 102134
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6652 137062 -6416
rect 137146 -6652 137382 -6416
rect 136826 -6972 137062 -6736
rect 137146 -6972 137382 -6736
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 141326 214718 141562 214954
rect 141646 214718 141882 214954
rect 141326 214398 141562 214634
rect 141646 214398 141882 214634
rect 141326 178718 141562 178954
rect 141646 178718 141882 178954
rect 141326 178398 141562 178634
rect 141646 178398 141882 178634
rect 141326 142718 141562 142954
rect 141646 142718 141882 142954
rect 141326 142398 141562 142634
rect 141646 142398 141882 142634
rect 141326 106718 141562 106954
rect 141646 106718 141882 106954
rect 141326 106398 141562 106634
rect 141646 106398 141882 106634
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 141326 -7612 141562 -7376
rect 141646 -7612 141882 -7376
rect 141326 -7932 141562 -7696
rect 141646 -7932 141882 -7696
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -892 146062 -656
rect 146146 -892 146382 -656
rect 145826 -1212 146062 -976
rect 146146 -1212 146382 -976
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 150326 223718 150562 223954
rect 150646 223718 150882 223954
rect 150326 223398 150562 223634
rect 150646 223398 150882 223634
rect 150326 187718 150562 187954
rect 150646 187718 150882 187954
rect 150326 187398 150562 187634
rect 150646 187398 150882 187634
rect 150326 151718 150562 151954
rect 150646 151718 150882 151954
rect 150326 151398 150562 151634
rect 150646 151398 150882 151634
rect 150326 115718 150562 115954
rect 150646 115718 150882 115954
rect 150326 115398 150562 115634
rect 150646 115398 150882 115634
rect 150326 79718 150562 79954
rect 150646 79718 150882 79954
rect 150326 79398 150562 79634
rect 150646 79398 150882 79634
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1852 150562 -1616
rect 150646 -1852 150882 -1616
rect 150326 -2172 150562 -1936
rect 150646 -2172 150882 -1936
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 154826 228218 155062 228454
rect 155146 228218 155382 228454
rect 154826 227898 155062 228134
rect 155146 227898 155382 228134
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 154826 156218 155062 156454
rect 155146 156218 155382 156454
rect 154826 155898 155062 156134
rect 155146 155898 155382 156134
rect 154826 120218 155062 120454
rect 155146 120218 155382 120454
rect 154826 119898 155062 120134
rect 155146 119898 155382 120134
rect 154826 84218 155062 84454
rect 155146 84218 155382 84454
rect 154826 83898 155062 84134
rect 155146 83898 155382 84134
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2812 155062 -2576
rect 155146 -2812 155382 -2576
rect 154826 -3132 155062 -2896
rect 155146 -3132 155382 -2896
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 159326 232718 159562 232954
rect 159646 232718 159882 232954
rect 159326 232398 159562 232634
rect 159646 232398 159882 232634
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 159326 160718 159562 160954
rect 159646 160718 159882 160954
rect 159326 160398 159562 160634
rect 159646 160398 159882 160634
rect 159326 124718 159562 124954
rect 159646 124718 159882 124954
rect 159326 124398 159562 124634
rect 159646 124398 159882 124634
rect 159326 88718 159562 88954
rect 159646 88718 159882 88954
rect 159326 88398 159562 88634
rect 159646 88398 159882 88634
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3772 159562 -3536
rect 159646 -3772 159882 -3536
rect 159326 -4092 159562 -3856
rect 159646 -4092 159882 -3856
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4732 164062 -4496
rect 164146 -4732 164382 -4496
rect 163826 -5052 164062 -4816
rect 164146 -5052 164382 -4816
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 168326 241718 168562 241954
rect 168646 241718 168882 241954
rect 168326 241398 168562 241634
rect 168646 241398 168882 241634
rect 168326 205718 168562 205954
rect 168646 205718 168882 205954
rect 168326 205398 168562 205634
rect 168646 205398 168882 205634
rect 168326 169718 168562 169954
rect 168646 169718 168882 169954
rect 168326 169398 168562 169634
rect 168646 169398 168882 169634
rect 168326 133718 168562 133954
rect 168646 133718 168882 133954
rect 168326 133398 168562 133634
rect 168646 133398 168882 133634
rect 168326 97718 168562 97954
rect 168646 97718 168882 97954
rect 168326 97398 168562 97634
rect 168646 97398 168882 97634
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5692 168562 -5456
rect 168646 -5692 168882 -5456
rect 168326 -6012 168562 -5776
rect 168646 -6012 168882 -5776
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 172826 246218 173062 246454
rect 173146 246218 173382 246454
rect 172826 245898 173062 246134
rect 173146 245898 173382 246134
rect 172826 210218 173062 210454
rect 173146 210218 173382 210454
rect 172826 209898 173062 210134
rect 173146 209898 173382 210134
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 172826 138218 173062 138454
rect 173146 138218 173382 138454
rect 172826 137898 173062 138134
rect 173146 137898 173382 138134
rect 172826 102218 173062 102454
rect 173146 102218 173382 102454
rect 172826 101898 173062 102134
rect 173146 101898 173382 102134
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6652 173062 -6416
rect 173146 -6652 173382 -6416
rect 172826 -6972 173062 -6736
rect 173146 -6972 173382 -6736
rect 177326 711632 177562 711868
rect 177646 711632 177882 711868
rect 177326 711312 177562 711548
rect 177646 711312 177882 711548
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 177326 214718 177562 214954
rect 177646 214718 177882 214954
rect 177326 214398 177562 214634
rect 177646 214398 177882 214634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 177326 106718 177562 106954
rect 177646 106718 177882 106954
rect 177326 106398 177562 106634
rect 177646 106398 177882 106634
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7612 177562 -7376
rect 177646 -7612 177882 -7376
rect 177326 -7932 177562 -7696
rect 177646 -7932 177882 -7696
rect 181826 704912 182062 705148
rect 182146 704912 182382 705148
rect 181826 704592 182062 704828
rect 182146 704592 182382 704828
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -892 182062 -656
rect 182146 -892 182382 -656
rect 181826 -1212 182062 -976
rect 182146 -1212 182382 -976
rect 186326 705872 186562 706108
rect 186646 705872 186882 706108
rect 186326 705552 186562 705788
rect 186646 705552 186882 705788
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1852 186562 -1616
rect 186646 -1852 186882 -1616
rect 186326 -2172 186562 -1936
rect 186646 -2172 186882 -1936
rect 190826 706832 191062 707068
rect 191146 706832 191382 707068
rect 190826 706512 191062 706748
rect 191146 706512 191382 706748
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 190826 228218 191062 228454
rect 191146 228218 191382 228454
rect 190826 227898 191062 228134
rect 191146 227898 191382 228134
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2812 191062 -2576
rect 191146 -2812 191382 -2576
rect 190826 -3132 191062 -2896
rect 191146 -3132 191382 -2896
rect 195326 707792 195562 708028
rect 195646 707792 195882 708028
rect 195326 707472 195562 707708
rect 195646 707472 195882 707708
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3772 195562 -3536
rect 195646 -3772 195882 -3536
rect 195326 -4092 195562 -3856
rect 195646 -4092 195882 -3856
rect 199826 708752 200062 708988
rect 200146 708752 200382 708988
rect 199826 708432 200062 708668
rect 200146 708432 200382 708668
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4732 200062 -4496
rect 200146 -4732 200382 -4496
rect 199826 -5052 200062 -4816
rect 200146 -5052 200382 -4816
rect 204326 709712 204562 709948
rect 204646 709712 204882 709948
rect 204326 709392 204562 709628
rect 204646 709392 204882 709628
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 204326 241718 204562 241954
rect 204646 241718 204882 241954
rect 204326 241398 204562 241634
rect 204646 241398 204882 241634
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5692 204562 -5456
rect 204646 -5692 204882 -5456
rect 204326 -6012 204562 -5776
rect 204646 -6012 204882 -5776
rect 208826 710672 209062 710908
rect 209146 710672 209382 710908
rect 208826 710352 209062 710588
rect 209146 710352 209382 710588
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 213326 711632 213562 711868
rect 213646 711632 213882 711868
rect 213326 711312 213562 711548
rect 213646 711312 213882 711548
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 217826 704912 218062 705148
rect 218146 704912 218382 705148
rect 217826 704592 218062 704828
rect 218146 704592 218382 704828
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 222326 705872 222562 706108
rect 222646 705872 222882 706108
rect 222326 705552 222562 705788
rect 222646 705552 222882 705788
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 226826 706832 227062 707068
rect 227146 706832 227382 707068
rect 226826 706512 227062 706748
rect 227146 706512 227382 706748
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 231326 707792 231562 708028
rect 231646 707792 231882 708028
rect 231326 707472 231562 707708
rect 231646 707472 231882 707708
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 235826 708752 236062 708988
rect 236146 708752 236382 708988
rect 235826 708432 236062 708668
rect 236146 708432 236382 708668
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 240326 709712 240562 709948
rect 240646 709712 240882 709948
rect 240326 709392 240562 709628
rect 240646 709392 240882 709628
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 244826 710672 245062 710908
rect 245146 710672 245382 710908
rect 244826 710352 245062 710588
rect 245146 710352 245382 710588
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 249326 711632 249562 711868
rect 249646 711632 249882 711868
rect 249326 711312 249562 711548
rect 249646 711312 249882 711548
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 253826 704912 254062 705148
rect 254146 704912 254382 705148
rect 253826 704592 254062 704828
rect 254146 704592 254382 704828
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 258326 705872 258562 706108
rect 258646 705872 258882 706108
rect 258326 705552 258562 705788
rect 258646 705552 258882 705788
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 262826 706832 263062 707068
rect 263146 706832 263382 707068
rect 262826 706512 263062 706748
rect 263146 706512 263382 706748
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 267326 707792 267562 708028
rect 267646 707792 267882 708028
rect 267326 707472 267562 707708
rect 267646 707472 267882 707708
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 271826 708752 272062 708988
rect 272146 708752 272382 708988
rect 271826 708432 272062 708668
rect 272146 708432 272382 708668
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 276326 709712 276562 709948
rect 276646 709712 276882 709948
rect 276326 709392 276562 709628
rect 276646 709392 276882 709628
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 280826 710672 281062 710908
rect 281146 710672 281382 710908
rect 280826 710352 281062 710588
rect 281146 710352 281382 710588
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 285326 711632 285562 711868
rect 285646 711632 285882 711868
rect 285326 711312 285562 711548
rect 285646 711312 285882 711548
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 289826 704912 290062 705148
rect 290146 704912 290382 705148
rect 289826 704592 290062 704828
rect 290146 704592 290382 704828
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 294326 705872 294562 706108
rect 294646 705872 294882 706108
rect 294326 705552 294562 705788
rect 294646 705552 294882 705788
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 298826 706832 299062 707068
rect 299146 706832 299382 707068
rect 298826 706512 299062 706748
rect 299146 706512 299382 706748
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 303326 707792 303562 708028
rect 303646 707792 303882 708028
rect 303326 707472 303562 707708
rect 303646 707472 303882 707708
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 307826 708752 308062 708988
rect 308146 708752 308382 708988
rect 307826 708432 308062 708668
rect 308146 708432 308382 708668
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 312326 709712 312562 709948
rect 312646 709712 312882 709948
rect 312326 709392 312562 709628
rect 312646 709392 312882 709628
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 316826 710672 317062 710908
rect 317146 710672 317382 710908
rect 316826 710352 317062 710588
rect 317146 710352 317382 710588
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 321326 711632 321562 711868
rect 321646 711632 321882 711868
rect 321326 711312 321562 711548
rect 321646 711312 321882 711548
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 325826 704912 326062 705148
rect 326146 704912 326382 705148
rect 325826 704592 326062 704828
rect 326146 704592 326382 704828
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 330326 705872 330562 706108
rect 330646 705872 330882 706108
rect 330326 705552 330562 705788
rect 330646 705552 330882 705788
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 334826 706832 335062 707068
rect 335146 706832 335382 707068
rect 334826 706512 335062 706748
rect 335146 706512 335382 706748
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 339326 707792 339562 708028
rect 339646 707792 339882 708028
rect 339326 707472 339562 707708
rect 339646 707472 339882 707708
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 343826 708752 344062 708988
rect 344146 708752 344382 708988
rect 343826 708432 344062 708668
rect 344146 708432 344382 708668
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 348326 709712 348562 709948
rect 348646 709712 348882 709948
rect 348326 709392 348562 709628
rect 348646 709392 348882 709628
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 352826 710672 353062 710908
rect 353146 710672 353382 710908
rect 352826 710352 353062 710588
rect 353146 710352 353382 710588
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 357326 711632 357562 711868
rect 357646 711632 357882 711868
rect 357326 711312 357562 711548
rect 357646 711312 357882 711548
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 361826 704912 362062 705148
rect 362146 704912 362382 705148
rect 361826 704592 362062 704828
rect 362146 704592 362382 704828
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 220328 547718 220564 547954
rect 220328 547398 220564 547634
rect 356056 547718 356292 547954
rect 356056 547398 356292 547634
rect 221008 543218 221244 543454
rect 221008 542898 221244 543134
rect 355376 543218 355612 543454
rect 355376 542898 355612 543134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 220328 511718 220564 511954
rect 220328 511398 220564 511634
rect 356056 511718 356292 511954
rect 356056 511398 356292 511634
rect 221008 507218 221244 507454
rect 221008 506898 221244 507134
rect 355376 507218 355612 507454
rect 355376 506898 355612 507134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 208826 246218 209062 246454
rect 209146 246218 209382 246454
rect 208826 245898 209062 246134
rect 209146 245898 209382 246134
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 208826 -6652 209062 -6416
rect 209146 -6652 209382 -6416
rect 208826 -6972 209062 -6736
rect 209146 -6972 209382 -6736
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 252010 403718 252246 403954
rect 252010 403398 252246 403634
rect 282730 403718 282966 403954
rect 282730 403398 282966 403634
rect 313450 403718 313686 403954
rect 313450 403398 313686 403634
rect 344170 403718 344406 403954
rect 344170 403398 344406 403634
rect 236650 399218 236886 399454
rect 236650 398898 236886 399134
rect 267370 399218 267606 399454
rect 267370 398898 267606 399134
rect 298090 399218 298326 399454
rect 298090 398898 298326 399134
rect 328810 399218 329046 399454
rect 328810 398898 329046 399134
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 252010 367718 252246 367954
rect 252010 367398 252246 367634
rect 282730 367718 282966 367954
rect 282730 367398 282966 367634
rect 313450 367718 313686 367954
rect 313450 367398 313686 367634
rect 344170 367718 344406 367954
rect 344170 367398 344406 367634
rect 236650 363218 236886 363454
rect 236650 362898 236886 363134
rect 267370 363218 267606 363454
rect 267370 362898 267606 363134
rect 298090 363218 298326 363454
rect 298090 362898 298326 363134
rect 328810 363218 329046 363454
rect 328810 362898 329046 363134
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 252010 331718 252246 331954
rect 252010 331398 252246 331634
rect 282730 331718 282966 331954
rect 282730 331398 282966 331634
rect 313450 331718 313686 331954
rect 313450 331398 313686 331634
rect 344170 331718 344406 331954
rect 344170 331398 344406 331634
rect 236650 327218 236886 327454
rect 236650 326898 236886 327134
rect 267370 327218 267606 327454
rect 267370 326898 267606 327134
rect 298090 327218 298326 327454
rect 298090 326898 298326 327134
rect 328810 327218 329046 327454
rect 328810 326898 329046 327134
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 244826 246218 245062 246454
rect 245146 246218 245382 246454
rect 244826 245898 245062 246134
rect 245146 245898 245382 246134
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 280826 246218 281062 246454
rect 281146 246218 281382 246454
rect 280826 245898 281062 246134
rect 281146 245898 281382 246134
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 316826 246218 317062 246454
rect 317146 246218 317382 246454
rect 316826 245898 317062 246134
rect 317146 245898 317382 246134
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 220328 223718 220564 223954
rect 220328 223398 220564 223634
rect 356056 223718 356292 223954
rect 356056 223398 356292 223634
rect 221008 219218 221244 219454
rect 221008 218898 221244 219134
rect 355376 219218 355612 219454
rect 355376 218898 355612 219134
rect 220328 187718 220564 187954
rect 220328 187398 220564 187634
rect 356056 187718 356292 187954
rect 356056 187398 356292 187634
rect 221008 183218 221244 183454
rect 221008 182898 221244 183134
rect 355376 183218 355612 183454
rect 355376 182898 355612 183134
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 213326 -7612 213562 -7376
rect 213646 -7612 213882 -7376
rect 213326 -7932 213562 -7696
rect 213646 -7932 213882 -7696
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -892 218062 -656
rect 218146 -892 218382 -656
rect 217826 -1212 218062 -976
rect 218146 -1212 218382 -976
rect 222326 -1852 222562 -1616
rect 222646 -1852 222882 -1616
rect 222326 -2172 222562 -1936
rect 222646 -2172 222882 -1936
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2812 227062 -2576
rect 227146 -2812 227382 -2576
rect 226826 -3132 227062 -2896
rect 227146 -3132 227382 -2896
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3772 231562 -3536
rect 231646 -3772 231882 -3536
rect 231326 -4092 231562 -3856
rect 231646 -4092 231882 -3856
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4732 236062 -4496
rect 236146 -4732 236382 -4496
rect 235826 -5052 236062 -4816
rect 236146 -5052 236382 -4816
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5692 240562 -5456
rect 240646 -5692 240882 -5456
rect 240326 -6012 240562 -5776
rect 240646 -6012 240882 -5776
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6652 245062 -6416
rect 245146 -6652 245382 -6416
rect 244826 -6972 245062 -6736
rect 245146 -6972 245382 -6736
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7612 249562 -7376
rect 249646 -7612 249882 -7376
rect 249326 -7932 249562 -7696
rect 249646 -7932 249882 -7696
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -892 254062 -656
rect 254146 -892 254382 -656
rect 253826 -1212 254062 -976
rect 254146 -1212 254382 -976
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1852 258562 -1616
rect 258646 -1852 258882 -1616
rect 258326 -2172 258562 -1936
rect 258646 -2172 258882 -1936
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2812 263062 -2576
rect 263146 -2812 263382 -2576
rect 262826 -3132 263062 -2896
rect 263146 -3132 263382 -2896
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3772 267562 -3536
rect 267646 -3772 267882 -3536
rect 267326 -4092 267562 -3856
rect 267646 -4092 267882 -3856
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4732 272062 -4496
rect 272146 -4732 272382 -4496
rect 271826 -5052 272062 -4816
rect 272146 -5052 272382 -4816
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5692 276562 -5456
rect 276646 -5692 276882 -5456
rect 276326 -6012 276562 -5776
rect 276646 -6012 276882 -5776
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6652 281062 -6416
rect 281146 -6652 281382 -6416
rect 280826 -6972 281062 -6736
rect 281146 -6972 281382 -6736
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7612 285562 -7376
rect 285646 -7612 285882 -7376
rect 285326 -7932 285562 -7696
rect 285646 -7932 285882 -7696
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -892 290062 -656
rect 290146 -892 290382 -656
rect 289826 -1212 290062 -976
rect 290146 -1212 290382 -976
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1852 294562 -1616
rect 294646 -1852 294882 -1616
rect 294326 -2172 294562 -1936
rect 294646 -2172 294882 -1936
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2812 299062 -2576
rect 299146 -2812 299382 -2576
rect 298826 -3132 299062 -2896
rect 299146 -3132 299382 -2896
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3772 303562 -3536
rect 303646 -3772 303882 -3536
rect 303326 -4092 303562 -3856
rect 303646 -4092 303882 -3856
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4732 308062 -4496
rect 308146 -4732 308382 -4496
rect 307826 -5052 308062 -4816
rect 308146 -5052 308382 -4816
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5692 312562 -5456
rect 312646 -5692 312882 -5456
rect 312326 -6012 312562 -5776
rect 312646 -6012 312882 -5776
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6652 317062 -6416
rect 317146 -6652 317382 -6416
rect 316826 -6972 317062 -6736
rect 317146 -6972 317382 -6736
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7612 321562 -7376
rect 321646 -7612 321882 -7376
rect 321326 -7932 321562 -7696
rect 321646 -7932 321882 -7696
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -892 326062 -656
rect 326146 -892 326382 -656
rect 325826 -1212 326062 -976
rect 326146 -1212 326382 -976
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1852 330562 -1616
rect 330646 -1852 330882 -1616
rect 330326 -2172 330562 -1936
rect 330646 -2172 330882 -1936
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2812 335062 -2576
rect 335146 -2812 335382 -2576
rect 334826 -3132 335062 -2896
rect 335146 -3132 335382 -2896
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3772 339562 -3536
rect 339646 -3772 339882 -3536
rect 339326 -4092 339562 -3856
rect 339646 -4092 339882 -3856
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4732 344062 -4496
rect 344146 -4732 344382 -4496
rect 343826 -5052 344062 -4816
rect 344146 -5052 344382 -4816
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5692 348562 -5456
rect 348646 -5692 348882 -5456
rect 348326 -6012 348562 -5776
rect 348646 -6012 348882 -5776
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6652 353062 -6416
rect 353146 -6652 353382 -6416
rect 352826 -6972 353062 -6736
rect 353146 -6972 353382 -6736
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 366326 705872 366562 706108
rect 366646 705872 366882 706108
rect 366326 705552 366562 705788
rect 366646 705552 366882 705788
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 370826 706832 371062 707068
rect 371146 706832 371382 707068
rect 370826 706512 371062 706748
rect 371146 706512 371382 706748
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 357326 -7612 357562 -7376
rect 357646 -7612 357882 -7376
rect 357326 -7932 357562 -7696
rect 357646 -7932 357882 -7696
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -892 362062 -656
rect 362146 -892 362382 -656
rect 361826 -1212 362062 -976
rect 362146 -1212 362382 -976
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 366326 -1852 366562 -1616
rect 366646 -1852 366882 -1616
rect 366326 -2172 366562 -1936
rect 366646 -2172 366882 -1936
rect 370826 -2812 371062 -2576
rect 371146 -2812 371382 -2576
rect 370826 -3132 371062 -2896
rect 371146 -3132 371382 -2896
rect 375326 707792 375562 708028
rect 375646 707792 375882 708028
rect 375326 707472 375562 707708
rect 375646 707472 375882 707708
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3772 375562 -3536
rect 375646 -3772 375882 -3536
rect 375326 -4092 375562 -3856
rect 375646 -4092 375882 -3856
rect 379826 708752 380062 708988
rect 380146 708752 380382 708988
rect 379826 708432 380062 708668
rect 380146 708432 380382 708668
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4732 380062 -4496
rect 380146 -4732 380382 -4496
rect 379826 -5052 380062 -4816
rect 380146 -5052 380382 -4816
rect 384326 709712 384562 709948
rect 384646 709712 384882 709948
rect 384326 709392 384562 709628
rect 384646 709392 384882 709628
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5692 384562 -5456
rect 384646 -5692 384882 -5456
rect 384326 -6012 384562 -5776
rect 384646 -6012 384882 -5776
rect 388826 710672 389062 710908
rect 389146 710672 389382 710908
rect 388826 710352 389062 710588
rect 389146 710352 389382 710588
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6652 389062 -6416
rect 389146 -6652 389382 -6416
rect 388826 -6972 389062 -6736
rect 389146 -6972 389382 -6736
rect 393326 711632 393562 711868
rect 393646 711632 393882 711868
rect 393326 711312 393562 711548
rect 393646 711312 393882 711548
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7612 393562 -7376
rect 393646 -7612 393882 -7376
rect 393326 -7932 393562 -7696
rect 393646 -7932 393882 -7696
rect 397826 704912 398062 705148
rect 398146 704912 398382 705148
rect 397826 704592 398062 704828
rect 398146 704592 398382 704828
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -892 398062 -656
rect 398146 -892 398382 -656
rect 397826 -1212 398062 -976
rect 398146 -1212 398382 -976
rect 402326 705872 402562 706108
rect 402646 705872 402882 706108
rect 402326 705552 402562 705788
rect 402646 705552 402882 705788
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1852 402562 -1616
rect 402646 -1852 402882 -1616
rect 402326 -2172 402562 -1936
rect 402646 -2172 402882 -1936
rect 406826 706832 407062 707068
rect 407146 706832 407382 707068
rect 406826 706512 407062 706748
rect 407146 706512 407382 706748
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2812 407062 -2576
rect 407146 -2812 407382 -2576
rect 406826 -3132 407062 -2896
rect 407146 -3132 407382 -2896
rect 411326 707792 411562 708028
rect 411646 707792 411882 708028
rect 411326 707472 411562 707708
rect 411646 707472 411882 707708
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3772 411562 -3536
rect 411646 -3772 411882 -3536
rect 411326 -4092 411562 -3856
rect 411646 -4092 411882 -3856
rect 415826 708752 416062 708988
rect 416146 708752 416382 708988
rect 415826 708432 416062 708668
rect 416146 708432 416382 708668
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4732 416062 -4496
rect 416146 -4732 416382 -4496
rect 415826 -5052 416062 -4816
rect 416146 -5052 416382 -4816
rect 420326 709712 420562 709948
rect 420646 709712 420882 709948
rect 420326 709392 420562 709628
rect 420646 709392 420882 709628
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5692 420562 -5456
rect 420646 -5692 420882 -5456
rect 420326 -6012 420562 -5776
rect 420646 -6012 420882 -5776
rect 424826 710672 425062 710908
rect 425146 710672 425382 710908
rect 424826 710352 425062 710588
rect 425146 710352 425382 710588
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6652 425062 -6416
rect 425146 -6652 425382 -6416
rect 424826 -6972 425062 -6736
rect 425146 -6972 425382 -6736
rect 429326 711632 429562 711868
rect 429646 711632 429882 711868
rect 429326 711312 429562 711548
rect 429646 711312 429882 711548
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7612 429562 -7376
rect 429646 -7612 429882 -7376
rect 429326 -7932 429562 -7696
rect 429646 -7932 429882 -7696
rect 433826 704912 434062 705148
rect 434146 704912 434382 705148
rect 433826 704592 434062 704828
rect 434146 704592 434382 704828
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -892 434062 -656
rect 434146 -892 434382 -656
rect 433826 -1212 434062 -976
rect 434146 -1212 434382 -976
rect 438326 705872 438562 706108
rect 438646 705872 438882 706108
rect 438326 705552 438562 705788
rect 438646 705552 438882 705788
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1852 438562 -1616
rect 438646 -1852 438882 -1616
rect 438326 -2172 438562 -1936
rect 438646 -2172 438882 -1936
rect 442826 706832 443062 707068
rect 443146 706832 443382 707068
rect 442826 706512 443062 706748
rect 443146 706512 443382 706748
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2812 443062 -2576
rect 443146 -2812 443382 -2576
rect 442826 -3132 443062 -2896
rect 443146 -3132 443382 -2896
rect 447326 707792 447562 708028
rect 447646 707792 447882 708028
rect 447326 707472 447562 707708
rect 447646 707472 447882 707708
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3772 447562 -3536
rect 447646 -3772 447882 -3536
rect 447326 -4092 447562 -3856
rect 447646 -4092 447882 -3856
rect 451826 708752 452062 708988
rect 452146 708752 452382 708988
rect 451826 708432 452062 708668
rect 452146 708432 452382 708668
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4732 452062 -4496
rect 452146 -4732 452382 -4496
rect 451826 -5052 452062 -4816
rect 452146 -5052 452382 -4816
rect 456326 709712 456562 709948
rect 456646 709712 456882 709948
rect 456326 709392 456562 709628
rect 456646 709392 456882 709628
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5692 456562 -5456
rect 456646 -5692 456882 -5456
rect 456326 -6012 456562 -5776
rect 456646 -6012 456882 -5776
rect 460826 710672 461062 710908
rect 461146 710672 461382 710908
rect 460826 710352 461062 710588
rect 461146 710352 461382 710588
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6652 461062 -6416
rect 461146 -6652 461382 -6416
rect 460826 -6972 461062 -6736
rect 461146 -6972 461382 -6736
rect 465326 711632 465562 711868
rect 465646 711632 465882 711868
rect 465326 711312 465562 711548
rect 465646 711312 465882 711548
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7612 465562 -7376
rect 465646 -7612 465882 -7376
rect 465326 -7932 465562 -7696
rect 465646 -7932 465882 -7696
rect 469826 704912 470062 705148
rect 470146 704912 470382 705148
rect 469826 704592 470062 704828
rect 470146 704592 470382 704828
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -892 470062 -656
rect 470146 -892 470382 -656
rect 469826 -1212 470062 -976
rect 470146 -1212 470382 -976
rect 474326 705872 474562 706108
rect 474646 705872 474882 706108
rect 474326 705552 474562 705788
rect 474646 705552 474882 705788
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1852 474562 -1616
rect 474646 -1852 474882 -1616
rect 474326 -2172 474562 -1936
rect 474646 -2172 474882 -1936
rect 478826 706832 479062 707068
rect 479146 706832 479382 707068
rect 478826 706512 479062 706748
rect 479146 706512 479382 706748
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2812 479062 -2576
rect 479146 -2812 479382 -2576
rect 478826 -3132 479062 -2896
rect 479146 -3132 479382 -2896
rect 483326 707792 483562 708028
rect 483646 707792 483882 708028
rect 483326 707472 483562 707708
rect 483646 707472 483882 707708
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3772 483562 -3536
rect 483646 -3772 483882 -3536
rect 483326 -4092 483562 -3856
rect 483646 -4092 483882 -3856
rect 487826 708752 488062 708988
rect 488146 708752 488382 708988
rect 487826 708432 488062 708668
rect 488146 708432 488382 708668
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4732 488062 -4496
rect 488146 -4732 488382 -4496
rect 487826 -5052 488062 -4816
rect 488146 -5052 488382 -4816
rect 492326 709712 492562 709948
rect 492646 709712 492882 709948
rect 492326 709392 492562 709628
rect 492646 709392 492882 709628
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5692 492562 -5456
rect 492646 -5692 492882 -5456
rect 492326 -6012 492562 -5776
rect 492646 -6012 492882 -5776
rect 496826 710672 497062 710908
rect 497146 710672 497382 710908
rect 496826 710352 497062 710588
rect 497146 710352 497382 710588
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6652 497062 -6416
rect 497146 -6652 497382 -6416
rect 496826 -6972 497062 -6736
rect 497146 -6972 497382 -6736
rect 501326 711632 501562 711868
rect 501646 711632 501882 711868
rect 501326 711312 501562 711548
rect 501646 711312 501882 711548
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7612 501562 -7376
rect 501646 -7612 501882 -7376
rect 501326 -7932 501562 -7696
rect 501646 -7932 501882 -7696
rect 505826 704912 506062 705148
rect 506146 704912 506382 705148
rect 505826 704592 506062 704828
rect 506146 704592 506382 704828
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -892 506062 -656
rect 506146 -892 506382 -656
rect 505826 -1212 506062 -976
rect 506146 -1212 506382 -976
rect 510326 705872 510562 706108
rect 510646 705872 510882 706108
rect 510326 705552 510562 705788
rect 510646 705552 510882 705788
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1852 510562 -1616
rect 510646 -1852 510882 -1616
rect 510326 -2172 510562 -1936
rect 510646 -2172 510882 -1936
rect 514826 706832 515062 707068
rect 515146 706832 515382 707068
rect 514826 706512 515062 706748
rect 515146 706512 515382 706748
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2812 515062 -2576
rect 515146 -2812 515382 -2576
rect 514826 -3132 515062 -2896
rect 515146 -3132 515382 -2896
rect 519326 707792 519562 708028
rect 519646 707792 519882 708028
rect 519326 707472 519562 707708
rect 519646 707472 519882 707708
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3772 519562 -3536
rect 519646 -3772 519882 -3536
rect 519326 -4092 519562 -3856
rect 519646 -4092 519882 -3856
rect 523826 708752 524062 708988
rect 524146 708752 524382 708988
rect 523826 708432 524062 708668
rect 524146 708432 524382 708668
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4732 524062 -4496
rect 524146 -4732 524382 -4496
rect 523826 -5052 524062 -4816
rect 524146 -5052 524382 -4816
rect 528326 709712 528562 709948
rect 528646 709712 528882 709948
rect 528326 709392 528562 709628
rect 528646 709392 528882 709628
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5692 528562 -5456
rect 528646 -5692 528882 -5456
rect 528326 -6012 528562 -5776
rect 528646 -6012 528882 -5776
rect 532826 710672 533062 710908
rect 533146 710672 533382 710908
rect 532826 710352 533062 710588
rect 533146 710352 533382 710588
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6652 533062 -6416
rect 533146 -6652 533382 -6416
rect 532826 -6972 533062 -6736
rect 533146 -6972 533382 -6736
rect 537326 711632 537562 711868
rect 537646 711632 537882 711868
rect 537326 711312 537562 711548
rect 537646 711312 537882 711548
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7612 537562 -7376
rect 537646 -7612 537882 -7376
rect 537326 -7932 537562 -7696
rect 537646 -7932 537882 -7696
rect 541826 704912 542062 705148
rect 542146 704912 542382 705148
rect 541826 704592 542062 704828
rect 542146 704592 542382 704828
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -892 542062 -656
rect 542146 -892 542382 -656
rect 541826 -1212 542062 -976
rect 542146 -1212 542382 -976
rect 546326 705872 546562 706108
rect 546646 705872 546882 706108
rect 546326 705552 546562 705788
rect 546646 705552 546882 705788
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1852 546562 -1616
rect 546646 -1852 546882 -1616
rect 546326 -2172 546562 -1936
rect 546646 -2172 546882 -1936
rect 550826 706832 551062 707068
rect 551146 706832 551382 707068
rect 550826 706512 551062 706748
rect 551146 706512 551382 706748
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2812 551062 -2576
rect 551146 -2812 551382 -2576
rect 550826 -3132 551062 -2896
rect 551146 -3132 551382 -2896
rect 555326 707792 555562 708028
rect 555646 707792 555882 708028
rect 555326 707472 555562 707708
rect 555646 707472 555882 707708
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3772 555562 -3536
rect 555646 -3772 555882 -3536
rect 555326 -4092 555562 -3856
rect 555646 -4092 555882 -3856
rect 559826 708752 560062 708988
rect 560146 708752 560382 708988
rect 559826 708432 560062 708668
rect 560146 708432 560382 708668
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4732 560062 -4496
rect 560146 -4732 560382 -4496
rect 559826 -5052 560062 -4816
rect 560146 -5052 560382 -4816
rect 564326 709712 564562 709948
rect 564646 709712 564882 709948
rect 564326 709392 564562 709628
rect 564646 709392 564882 709628
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5692 564562 -5456
rect 564646 -5692 564882 -5456
rect 564326 -6012 564562 -5776
rect 564646 -6012 564882 -5776
rect 568826 710672 569062 710908
rect 569146 710672 569382 710908
rect 568826 710352 569062 710588
rect 569146 710352 569382 710588
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6652 569062 -6416
rect 569146 -6652 569382 -6416
rect 568826 -6972 569062 -6736
rect 569146 -6972 569382 -6736
rect 573326 711632 573562 711868
rect 573646 711632 573882 711868
rect 573326 711312 573562 711548
rect 573646 711312 573882 711548
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7612 573562 -7376
rect 573646 -7612 573882 -7376
rect 573326 -7932 573562 -7696
rect 573646 -7932 573882 -7696
rect 577826 704912 578062 705148
rect 578146 704912 578382 705148
rect 577826 704592 578062 704828
rect 578146 704592 578382 704828
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -892 578062 -656
rect 578146 -892 578382 -656
rect 577826 -1212 578062 -976
rect 578146 -1212 578382 -976
rect 592372 711632 592608 711868
rect 592692 711632 592928 711868
rect 592372 711312 592608 711548
rect 592692 711312 592928 711548
rect 591412 710672 591648 710908
rect 591732 710672 591968 710908
rect 591412 710352 591648 710588
rect 591732 710352 591968 710588
rect 590452 709712 590688 709948
rect 590772 709712 591008 709948
rect 590452 709392 590688 709628
rect 590772 709392 591008 709628
rect 589492 708752 589728 708988
rect 589812 708752 590048 708988
rect 589492 708432 589728 708668
rect 589812 708432 590048 708668
rect 588532 707792 588768 708028
rect 588852 707792 589088 708028
rect 588532 707472 588768 707708
rect 588852 707472 589088 707708
rect 587572 706832 587808 707068
rect 587892 706832 588128 707068
rect 587572 706512 587808 706748
rect 587892 706512 588128 706748
rect 582326 705872 582562 706108
rect 582646 705872 582882 706108
rect 582326 705552 582562 705788
rect 582646 705552 582882 705788
rect 586612 705872 586848 706108
rect 586932 705872 587168 706108
rect 586612 705552 586848 705788
rect 586932 705552 587168 705788
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585652 704912 585888 705148
rect 585972 704912 586208 705148
rect 585652 704592 585888 704828
rect 585972 704592 586208 704828
rect 585652 687218 585888 687454
rect 585972 687218 586208 687454
rect 585652 686898 585888 687134
rect 585972 686898 586208 687134
rect 585652 651218 585888 651454
rect 585972 651218 586208 651454
rect 585652 650898 585888 651134
rect 585972 650898 586208 651134
rect 585652 615218 585888 615454
rect 585972 615218 586208 615454
rect 585652 614898 585888 615134
rect 585972 614898 586208 615134
rect 585652 579218 585888 579454
rect 585972 579218 586208 579454
rect 585652 578898 585888 579134
rect 585972 578898 586208 579134
rect 585652 543218 585888 543454
rect 585972 543218 586208 543454
rect 585652 542898 585888 543134
rect 585972 542898 586208 543134
rect 585652 507218 585888 507454
rect 585972 507218 586208 507454
rect 585652 506898 585888 507134
rect 585972 506898 586208 507134
rect 585652 471218 585888 471454
rect 585972 471218 586208 471454
rect 585652 470898 585888 471134
rect 585972 470898 586208 471134
rect 585652 435218 585888 435454
rect 585972 435218 586208 435454
rect 585652 434898 585888 435134
rect 585972 434898 586208 435134
rect 585652 399218 585888 399454
rect 585972 399218 586208 399454
rect 585652 398898 585888 399134
rect 585972 398898 586208 399134
rect 585652 363218 585888 363454
rect 585972 363218 586208 363454
rect 585652 362898 585888 363134
rect 585972 362898 586208 363134
rect 585652 327218 585888 327454
rect 585972 327218 586208 327454
rect 585652 326898 585888 327134
rect 585972 326898 586208 327134
rect 585652 291218 585888 291454
rect 585972 291218 586208 291454
rect 585652 290898 585888 291134
rect 585972 290898 586208 291134
rect 585652 255218 585888 255454
rect 585972 255218 586208 255454
rect 585652 254898 585888 255134
rect 585972 254898 586208 255134
rect 585652 219218 585888 219454
rect 585972 219218 586208 219454
rect 585652 218898 585888 219134
rect 585972 218898 586208 219134
rect 585652 183218 585888 183454
rect 585972 183218 586208 183454
rect 585652 182898 585888 183134
rect 585972 182898 586208 183134
rect 585652 147218 585888 147454
rect 585972 147218 586208 147454
rect 585652 146898 585888 147134
rect 585972 146898 586208 147134
rect 585652 111218 585888 111454
rect 585972 111218 586208 111454
rect 585652 110898 585888 111134
rect 585972 110898 586208 111134
rect 585652 75218 585888 75454
rect 585972 75218 586208 75454
rect 585652 74898 585888 75134
rect 585972 74898 586208 75134
rect 585652 39218 585888 39454
rect 585972 39218 586208 39454
rect 585652 38898 585888 39134
rect 585972 38898 586208 39134
rect 585652 3218 585888 3454
rect 585972 3218 586208 3454
rect 585652 2898 585888 3134
rect 585972 2898 586208 3134
rect 585652 -892 585888 -656
rect 585972 -892 586208 -656
rect 585652 -1212 585888 -976
rect 585972 -1212 586208 -976
rect 586612 691718 586848 691954
rect 586932 691718 587168 691954
rect 586612 691398 586848 691634
rect 586932 691398 587168 691634
rect 586612 655718 586848 655954
rect 586932 655718 587168 655954
rect 586612 655398 586848 655634
rect 586932 655398 587168 655634
rect 586612 619718 586848 619954
rect 586932 619718 587168 619954
rect 586612 619398 586848 619634
rect 586932 619398 587168 619634
rect 586612 583718 586848 583954
rect 586932 583718 587168 583954
rect 586612 583398 586848 583634
rect 586932 583398 587168 583634
rect 586612 547718 586848 547954
rect 586932 547718 587168 547954
rect 586612 547398 586848 547634
rect 586932 547398 587168 547634
rect 586612 511718 586848 511954
rect 586932 511718 587168 511954
rect 586612 511398 586848 511634
rect 586932 511398 587168 511634
rect 586612 475718 586848 475954
rect 586932 475718 587168 475954
rect 586612 475398 586848 475634
rect 586932 475398 587168 475634
rect 586612 439718 586848 439954
rect 586932 439718 587168 439954
rect 586612 439398 586848 439634
rect 586932 439398 587168 439634
rect 586612 403718 586848 403954
rect 586932 403718 587168 403954
rect 586612 403398 586848 403634
rect 586932 403398 587168 403634
rect 586612 367718 586848 367954
rect 586932 367718 587168 367954
rect 586612 367398 586848 367634
rect 586932 367398 587168 367634
rect 586612 331718 586848 331954
rect 586932 331718 587168 331954
rect 586612 331398 586848 331634
rect 586932 331398 587168 331634
rect 586612 295718 586848 295954
rect 586932 295718 587168 295954
rect 586612 295398 586848 295634
rect 586932 295398 587168 295634
rect 586612 259718 586848 259954
rect 586932 259718 587168 259954
rect 586612 259398 586848 259634
rect 586932 259398 587168 259634
rect 586612 223718 586848 223954
rect 586932 223718 587168 223954
rect 586612 223398 586848 223634
rect 586932 223398 587168 223634
rect 586612 187718 586848 187954
rect 586932 187718 587168 187954
rect 586612 187398 586848 187634
rect 586932 187398 587168 187634
rect 586612 151718 586848 151954
rect 586932 151718 587168 151954
rect 586612 151398 586848 151634
rect 586932 151398 587168 151634
rect 586612 115718 586848 115954
rect 586932 115718 587168 115954
rect 586612 115398 586848 115634
rect 586932 115398 587168 115634
rect 586612 79718 586848 79954
rect 586932 79718 587168 79954
rect 586612 79398 586848 79634
rect 586932 79398 587168 79634
rect 586612 43718 586848 43954
rect 586932 43718 587168 43954
rect 586612 43398 586848 43634
rect 586932 43398 587168 43634
rect 586612 7718 586848 7954
rect 586932 7718 587168 7954
rect 586612 7398 586848 7634
rect 586932 7398 587168 7634
rect 582326 -1852 582562 -1616
rect 582646 -1852 582882 -1616
rect 582326 -2172 582562 -1936
rect 582646 -2172 582882 -1936
rect 586612 -1852 586848 -1616
rect 586932 -1852 587168 -1616
rect 586612 -2172 586848 -1936
rect 586932 -2172 587168 -1936
rect 587572 696218 587808 696454
rect 587892 696218 588128 696454
rect 587572 695898 587808 696134
rect 587892 695898 588128 696134
rect 587572 660218 587808 660454
rect 587892 660218 588128 660454
rect 587572 659898 587808 660134
rect 587892 659898 588128 660134
rect 587572 624218 587808 624454
rect 587892 624218 588128 624454
rect 587572 623898 587808 624134
rect 587892 623898 588128 624134
rect 587572 588218 587808 588454
rect 587892 588218 588128 588454
rect 587572 587898 587808 588134
rect 587892 587898 588128 588134
rect 587572 552218 587808 552454
rect 587892 552218 588128 552454
rect 587572 551898 587808 552134
rect 587892 551898 588128 552134
rect 587572 516218 587808 516454
rect 587892 516218 588128 516454
rect 587572 515898 587808 516134
rect 587892 515898 588128 516134
rect 587572 480218 587808 480454
rect 587892 480218 588128 480454
rect 587572 479898 587808 480134
rect 587892 479898 588128 480134
rect 587572 444218 587808 444454
rect 587892 444218 588128 444454
rect 587572 443898 587808 444134
rect 587892 443898 588128 444134
rect 587572 408218 587808 408454
rect 587892 408218 588128 408454
rect 587572 407898 587808 408134
rect 587892 407898 588128 408134
rect 587572 372218 587808 372454
rect 587892 372218 588128 372454
rect 587572 371898 587808 372134
rect 587892 371898 588128 372134
rect 587572 336218 587808 336454
rect 587892 336218 588128 336454
rect 587572 335898 587808 336134
rect 587892 335898 588128 336134
rect 587572 300218 587808 300454
rect 587892 300218 588128 300454
rect 587572 299898 587808 300134
rect 587892 299898 588128 300134
rect 587572 264218 587808 264454
rect 587892 264218 588128 264454
rect 587572 263898 587808 264134
rect 587892 263898 588128 264134
rect 587572 228218 587808 228454
rect 587892 228218 588128 228454
rect 587572 227898 587808 228134
rect 587892 227898 588128 228134
rect 587572 192218 587808 192454
rect 587892 192218 588128 192454
rect 587572 191898 587808 192134
rect 587892 191898 588128 192134
rect 587572 156218 587808 156454
rect 587892 156218 588128 156454
rect 587572 155898 587808 156134
rect 587892 155898 588128 156134
rect 587572 120218 587808 120454
rect 587892 120218 588128 120454
rect 587572 119898 587808 120134
rect 587892 119898 588128 120134
rect 587572 84218 587808 84454
rect 587892 84218 588128 84454
rect 587572 83898 587808 84134
rect 587892 83898 588128 84134
rect 587572 48218 587808 48454
rect 587892 48218 588128 48454
rect 587572 47898 587808 48134
rect 587892 47898 588128 48134
rect 587572 12218 587808 12454
rect 587892 12218 588128 12454
rect 587572 11898 587808 12134
rect 587892 11898 588128 12134
rect 587572 -2812 587808 -2576
rect 587892 -2812 588128 -2576
rect 587572 -3132 587808 -2896
rect 587892 -3132 588128 -2896
rect 588532 700718 588768 700954
rect 588852 700718 589088 700954
rect 588532 700398 588768 700634
rect 588852 700398 589088 700634
rect 588532 664718 588768 664954
rect 588852 664718 589088 664954
rect 588532 664398 588768 664634
rect 588852 664398 589088 664634
rect 588532 628718 588768 628954
rect 588852 628718 589088 628954
rect 588532 628398 588768 628634
rect 588852 628398 589088 628634
rect 588532 592718 588768 592954
rect 588852 592718 589088 592954
rect 588532 592398 588768 592634
rect 588852 592398 589088 592634
rect 588532 556718 588768 556954
rect 588852 556718 589088 556954
rect 588532 556398 588768 556634
rect 588852 556398 589088 556634
rect 588532 520718 588768 520954
rect 588852 520718 589088 520954
rect 588532 520398 588768 520634
rect 588852 520398 589088 520634
rect 588532 484718 588768 484954
rect 588852 484718 589088 484954
rect 588532 484398 588768 484634
rect 588852 484398 589088 484634
rect 588532 448718 588768 448954
rect 588852 448718 589088 448954
rect 588532 448398 588768 448634
rect 588852 448398 589088 448634
rect 588532 412718 588768 412954
rect 588852 412718 589088 412954
rect 588532 412398 588768 412634
rect 588852 412398 589088 412634
rect 588532 376718 588768 376954
rect 588852 376718 589088 376954
rect 588532 376398 588768 376634
rect 588852 376398 589088 376634
rect 588532 340718 588768 340954
rect 588852 340718 589088 340954
rect 588532 340398 588768 340634
rect 588852 340398 589088 340634
rect 588532 304718 588768 304954
rect 588852 304718 589088 304954
rect 588532 304398 588768 304634
rect 588852 304398 589088 304634
rect 588532 268718 588768 268954
rect 588852 268718 589088 268954
rect 588532 268398 588768 268634
rect 588852 268398 589088 268634
rect 588532 232718 588768 232954
rect 588852 232718 589088 232954
rect 588532 232398 588768 232634
rect 588852 232398 589088 232634
rect 588532 196718 588768 196954
rect 588852 196718 589088 196954
rect 588532 196398 588768 196634
rect 588852 196398 589088 196634
rect 588532 160718 588768 160954
rect 588852 160718 589088 160954
rect 588532 160398 588768 160634
rect 588852 160398 589088 160634
rect 588532 124718 588768 124954
rect 588852 124718 589088 124954
rect 588532 124398 588768 124634
rect 588852 124398 589088 124634
rect 588532 88718 588768 88954
rect 588852 88718 589088 88954
rect 588532 88398 588768 88634
rect 588852 88398 589088 88634
rect 588532 52718 588768 52954
rect 588852 52718 589088 52954
rect 588532 52398 588768 52634
rect 588852 52398 589088 52634
rect 588532 16718 588768 16954
rect 588852 16718 589088 16954
rect 588532 16398 588768 16634
rect 588852 16398 589088 16634
rect 588532 -3772 588768 -3536
rect 588852 -3772 589088 -3536
rect 588532 -4092 588768 -3856
rect 588852 -4092 589088 -3856
rect 589492 669218 589728 669454
rect 589812 669218 590048 669454
rect 589492 668898 589728 669134
rect 589812 668898 590048 669134
rect 589492 633218 589728 633454
rect 589812 633218 590048 633454
rect 589492 632898 589728 633134
rect 589812 632898 590048 633134
rect 589492 597218 589728 597454
rect 589812 597218 590048 597454
rect 589492 596898 589728 597134
rect 589812 596898 590048 597134
rect 589492 561218 589728 561454
rect 589812 561218 590048 561454
rect 589492 560898 589728 561134
rect 589812 560898 590048 561134
rect 589492 525218 589728 525454
rect 589812 525218 590048 525454
rect 589492 524898 589728 525134
rect 589812 524898 590048 525134
rect 589492 489218 589728 489454
rect 589812 489218 590048 489454
rect 589492 488898 589728 489134
rect 589812 488898 590048 489134
rect 589492 453218 589728 453454
rect 589812 453218 590048 453454
rect 589492 452898 589728 453134
rect 589812 452898 590048 453134
rect 589492 417218 589728 417454
rect 589812 417218 590048 417454
rect 589492 416898 589728 417134
rect 589812 416898 590048 417134
rect 589492 381218 589728 381454
rect 589812 381218 590048 381454
rect 589492 380898 589728 381134
rect 589812 380898 590048 381134
rect 589492 345218 589728 345454
rect 589812 345218 590048 345454
rect 589492 344898 589728 345134
rect 589812 344898 590048 345134
rect 589492 309218 589728 309454
rect 589812 309218 590048 309454
rect 589492 308898 589728 309134
rect 589812 308898 590048 309134
rect 589492 273218 589728 273454
rect 589812 273218 590048 273454
rect 589492 272898 589728 273134
rect 589812 272898 590048 273134
rect 589492 237218 589728 237454
rect 589812 237218 590048 237454
rect 589492 236898 589728 237134
rect 589812 236898 590048 237134
rect 589492 201218 589728 201454
rect 589812 201218 590048 201454
rect 589492 200898 589728 201134
rect 589812 200898 590048 201134
rect 589492 165218 589728 165454
rect 589812 165218 590048 165454
rect 589492 164898 589728 165134
rect 589812 164898 590048 165134
rect 589492 129218 589728 129454
rect 589812 129218 590048 129454
rect 589492 128898 589728 129134
rect 589812 128898 590048 129134
rect 589492 93218 589728 93454
rect 589812 93218 590048 93454
rect 589492 92898 589728 93134
rect 589812 92898 590048 93134
rect 589492 57218 589728 57454
rect 589812 57218 590048 57454
rect 589492 56898 589728 57134
rect 589812 56898 590048 57134
rect 589492 21218 589728 21454
rect 589812 21218 590048 21454
rect 589492 20898 589728 21134
rect 589812 20898 590048 21134
rect 589492 -4732 589728 -4496
rect 589812 -4732 590048 -4496
rect 589492 -5052 589728 -4816
rect 589812 -5052 590048 -4816
rect 590452 673718 590688 673954
rect 590772 673718 591008 673954
rect 590452 673398 590688 673634
rect 590772 673398 591008 673634
rect 590452 637718 590688 637954
rect 590772 637718 591008 637954
rect 590452 637398 590688 637634
rect 590772 637398 591008 637634
rect 590452 601718 590688 601954
rect 590772 601718 591008 601954
rect 590452 601398 590688 601634
rect 590772 601398 591008 601634
rect 590452 565718 590688 565954
rect 590772 565718 591008 565954
rect 590452 565398 590688 565634
rect 590772 565398 591008 565634
rect 590452 529718 590688 529954
rect 590772 529718 591008 529954
rect 590452 529398 590688 529634
rect 590772 529398 591008 529634
rect 590452 493718 590688 493954
rect 590772 493718 591008 493954
rect 590452 493398 590688 493634
rect 590772 493398 591008 493634
rect 590452 457718 590688 457954
rect 590772 457718 591008 457954
rect 590452 457398 590688 457634
rect 590772 457398 591008 457634
rect 590452 421718 590688 421954
rect 590772 421718 591008 421954
rect 590452 421398 590688 421634
rect 590772 421398 591008 421634
rect 590452 385718 590688 385954
rect 590772 385718 591008 385954
rect 590452 385398 590688 385634
rect 590772 385398 591008 385634
rect 590452 349718 590688 349954
rect 590772 349718 591008 349954
rect 590452 349398 590688 349634
rect 590772 349398 591008 349634
rect 590452 313718 590688 313954
rect 590772 313718 591008 313954
rect 590452 313398 590688 313634
rect 590772 313398 591008 313634
rect 590452 277718 590688 277954
rect 590772 277718 591008 277954
rect 590452 277398 590688 277634
rect 590772 277398 591008 277634
rect 590452 241718 590688 241954
rect 590772 241718 591008 241954
rect 590452 241398 590688 241634
rect 590772 241398 591008 241634
rect 590452 205718 590688 205954
rect 590772 205718 591008 205954
rect 590452 205398 590688 205634
rect 590772 205398 591008 205634
rect 590452 169718 590688 169954
rect 590772 169718 591008 169954
rect 590452 169398 590688 169634
rect 590772 169398 591008 169634
rect 590452 133718 590688 133954
rect 590772 133718 591008 133954
rect 590452 133398 590688 133634
rect 590772 133398 591008 133634
rect 590452 97718 590688 97954
rect 590772 97718 591008 97954
rect 590452 97398 590688 97634
rect 590772 97398 591008 97634
rect 590452 61718 590688 61954
rect 590772 61718 591008 61954
rect 590452 61398 590688 61634
rect 590772 61398 591008 61634
rect 590452 25718 590688 25954
rect 590772 25718 591008 25954
rect 590452 25398 590688 25634
rect 590772 25398 591008 25634
rect 590452 -5692 590688 -5456
rect 590772 -5692 591008 -5456
rect 590452 -6012 590688 -5776
rect 590772 -6012 591008 -5776
rect 591412 678218 591648 678454
rect 591732 678218 591968 678454
rect 591412 677898 591648 678134
rect 591732 677898 591968 678134
rect 591412 642218 591648 642454
rect 591732 642218 591968 642454
rect 591412 641898 591648 642134
rect 591732 641898 591968 642134
rect 591412 606218 591648 606454
rect 591732 606218 591968 606454
rect 591412 605898 591648 606134
rect 591732 605898 591968 606134
rect 591412 570218 591648 570454
rect 591732 570218 591968 570454
rect 591412 569898 591648 570134
rect 591732 569898 591968 570134
rect 591412 534218 591648 534454
rect 591732 534218 591968 534454
rect 591412 533898 591648 534134
rect 591732 533898 591968 534134
rect 591412 498218 591648 498454
rect 591732 498218 591968 498454
rect 591412 497898 591648 498134
rect 591732 497898 591968 498134
rect 591412 462218 591648 462454
rect 591732 462218 591968 462454
rect 591412 461898 591648 462134
rect 591732 461898 591968 462134
rect 591412 426218 591648 426454
rect 591732 426218 591968 426454
rect 591412 425898 591648 426134
rect 591732 425898 591968 426134
rect 591412 390218 591648 390454
rect 591732 390218 591968 390454
rect 591412 389898 591648 390134
rect 591732 389898 591968 390134
rect 591412 354218 591648 354454
rect 591732 354218 591968 354454
rect 591412 353898 591648 354134
rect 591732 353898 591968 354134
rect 591412 318218 591648 318454
rect 591732 318218 591968 318454
rect 591412 317898 591648 318134
rect 591732 317898 591968 318134
rect 591412 282218 591648 282454
rect 591732 282218 591968 282454
rect 591412 281898 591648 282134
rect 591732 281898 591968 282134
rect 591412 246218 591648 246454
rect 591732 246218 591968 246454
rect 591412 245898 591648 246134
rect 591732 245898 591968 246134
rect 591412 210218 591648 210454
rect 591732 210218 591968 210454
rect 591412 209898 591648 210134
rect 591732 209898 591968 210134
rect 591412 174218 591648 174454
rect 591732 174218 591968 174454
rect 591412 173898 591648 174134
rect 591732 173898 591968 174134
rect 591412 138218 591648 138454
rect 591732 138218 591968 138454
rect 591412 137898 591648 138134
rect 591732 137898 591968 138134
rect 591412 102218 591648 102454
rect 591732 102218 591968 102454
rect 591412 101898 591648 102134
rect 591732 101898 591968 102134
rect 591412 66218 591648 66454
rect 591732 66218 591968 66454
rect 591412 65898 591648 66134
rect 591732 65898 591968 66134
rect 591412 30218 591648 30454
rect 591732 30218 591968 30454
rect 591412 29898 591648 30134
rect 591732 29898 591968 30134
rect 591412 -6652 591648 -6416
rect 591732 -6652 591968 -6416
rect 591412 -6972 591648 -6736
rect 591732 -6972 591968 -6736
rect 592372 682718 592608 682954
rect 592692 682718 592928 682954
rect 592372 682398 592608 682634
rect 592692 682398 592928 682634
rect 592372 646718 592608 646954
rect 592692 646718 592928 646954
rect 592372 646398 592608 646634
rect 592692 646398 592928 646634
rect 592372 610718 592608 610954
rect 592692 610718 592928 610954
rect 592372 610398 592608 610634
rect 592692 610398 592928 610634
rect 592372 574718 592608 574954
rect 592692 574718 592928 574954
rect 592372 574398 592608 574634
rect 592692 574398 592928 574634
rect 592372 538718 592608 538954
rect 592692 538718 592928 538954
rect 592372 538398 592608 538634
rect 592692 538398 592928 538634
rect 592372 502718 592608 502954
rect 592692 502718 592928 502954
rect 592372 502398 592608 502634
rect 592692 502398 592928 502634
rect 592372 466718 592608 466954
rect 592692 466718 592928 466954
rect 592372 466398 592608 466634
rect 592692 466398 592928 466634
rect 592372 430718 592608 430954
rect 592692 430718 592928 430954
rect 592372 430398 592608 430634
rect 592692 430398 592928 430634
rect 592372 394718 592608 394954
rect 592692 394718 592928 394954
rect 592372 394398 592608 394634
rect 592692 394398 592928 394634
rect 592372 358718 592608 358954
rect 592692 358718 592928 358954
rect 592372 358398 592608 358634
rect 592692 358398 592928 358634
rect 592372 322718 592608 322954
rect 592692 322718 592928 322954
rect 592372 322398 592608 322634
rect 592692 322398 592928 322634
rect 592372 286718 592608 286954
rect 592692 286718 592928 286954
rect 592372 286398 592608 286634
rect 592692 286398 592928 286634
rect 592372 250718 592608 250954
rect 592692 250718 592928 250954
rect 592372 250398 592608 250634
rect 592692 250398 592928 250634
rect 592372 214718 592608 214954
rect 592692 214718 592928 214954
rect 592372 214398 592608 214634
rect 592692 214398 592928 214634
rect 592372 178718 592608 178954
rect 592692 178718 592928 178954
rect 592372 178398 592608 178634
rect 592692 178398 592928 178634
rect 592372 142718 592608 142954
rect 592692 142718 592928 142954
rect 592372 142398 592608 142634
rect 592692 142398 592928 142634
rect 592372 106718 592608 106954
rect 592692 106718 592928 106954
rect 592372 106398 592608 106634
rect 592692 106398 592928 106634
rect 592372 70718 592608 70954
rect 592692 70718 592928 70954
rect 592372 70398 592608 70634
rect 592692 70398 592928 70634
rect 592372 34718 592608 34954
rect 592692 34718 592928 34954
rect 592372 34398 592608 34634
rect 592692 34398 592928 34634
rect 592372 -7612 592608 -7376
rect 592692 -7612 592928 -7376
rect 592372 -7932 592608 -7696
rect 592692 -7932 592928 -7696
<< metal5 >>
rect -9036 711868 592960 711900
rect -9036 711632 -9004 711868
rect -8768 711632 -8684 711868
rect -8448 711632 33326 711868
rect 33562 711632 33646 711868
rect 33882 711632 69326 711868
rect 69562 711632 69646 711868
rect 69882 711632 105326 711868
rect 105562 711632 105646 711868
rect 105882 711632 141326 711868
rect 141562 711632 141646 711868
rect 141882 711632 177326 711868
rect 177562 711632 177646 711868
rect 177882 711632 213326 711868
rect 213562 711632 213646 711868
rect 213882 711632 249326 711868
rect 249562 711632 249646 711868
rect 249882 711632 285326 711868
rect 285562 711632 285646 711868
rect 285882 711632 321326 711868
rect 321562 711632 321646 711868
rect 321882 711632 357326 711868
rect 357562 711632 357646 711868
rect 357882 711632 393326 711868
rect 393562 711632 393646 711868
rect 393882 711632 429326 711868
rect 429562 711632 429646 711868
rect 429882 711632 465326 711868
rect 465562 711632 465646 711868
rect 465882 711632 501326 711868
rect 501562 711632 501646 711868
rect 501882 711632 537326 711868
rect 537562 711632 537646 711868
rect 537882 711632 573326 711868
rect 573562 711632 573646 711868
rect 573882 711632 592372 711868
rect 592608 711632 592692 711868
rect 592928 711632 592960 711868
rect -9036 711548 592960 711632
rect -9036 711312 -9004 711548
rect -8768 711312 -8684 711548
rect -8448 711312 33326 711548
rect 33562 711312 33646 711548
rect 33882 711312 69326 711548
rect 69562 711312 69646 711548
rect 69882 711312 105326 711548
rect 105562 711312 105646 711548
rect 105882 711312 141326 711548
rect 141562 711312 141646 711548
rect 141882 711312 177326 711548
rect 177562 711312 177646 711548
rect 177882 711312 213326 711548
rect 213562 711312 213646 711548
rect 213882 711312 249326 711548
rect 249562 711312 249646 711548
rect 249882 711312 285326 711548
rect 285562 711312 285646 711548
rect 285882 711312 321326 711548
rect 321562 711312 321646 711548
rect 321882 711312 357326 711548
rect 357562 711312 357646 711548
rect 357882 711312 393326 711548
rect 393562 711312 393646 711548
rect 393882 711312 429326 711548
rect 429562 711312 429646 711548
rect 429882 711312 465326 711548
rect 465562 711312 465646 711548
rect 465882 711312 501326 711548
rect 501562 711312 501646 711548
rect 501882 711312 537326 711548
rect 537562 711312 537646 711548
rect 537882 711312 573326 711548
rect 573562 711312 573646 711548
rect 573882 711312 592372 711548
rect 592608 711312 592692 711548
rect 592928 711312 592960 711548
rect -9036 711280 592960 711312
rect -8076 710908 592000 710940
rect -8076 710672 -8044 710908
rect -7808 710672 -7724 710908
rect -7488 710672 28826 710908
rect 29062 710672 29146 710908
rect 29382 710672 64826 710908
rect 65062 710672 65146 710908
rect 65382 710672 100826 710908
rect 101062 710672 101146 710908
rect 101382 710672 136826 710908
rect 137062 710672 137146 710908
rect 137382 710672 172826 710908
rect 173062 710672 173146 710908
rect 173382 710672 208826 710908
rect 209062 710672 209146 710908
rect 209382 710672 244826 710908
rect 245062 710672 245146 710908
rect 245382 710672 280826 710908
rect 281062 710672 281146 710908
rect 281382 710672 316826 710908
rect 317062 710672 317146 710908
rect 317382 710672 352826 710908
rect 353062 710672 353146 710908
rect 353382 710672 388826 710908
rect 389062 710672 389146 710908
rect 389382 710672 424826 710908
rect 425062 710672 425146 710908
rect 425382 710672 460826 710908
rect 461062 710672 461146 710908
rect 461382 710672 496826 710908
rect 497062 710672 497146 710908
rect 497382 710672 532826 710908
rect 533062 710672 533146 710908
rect 533382 710672 568826 710908
rect 569062 710672 569146 710908
rect 569382 710672 591412 710908
rect 591648 710672 591732 710908
rect 591968 710672 592000 710908
rect -8076 710588 592000 710672
rect -8076 710352 -8044 710588
rect -7808 710352 -7724 710588
rect -7488 710352 28826 710588
rect 29062 710352 29146 710588
rect 29382 710352 64826 710588
rect 65062 710352 65146 710588
rect 65382 710352 100826 710588
rect 101062 710352 101146 710588
rect 101382 710352 136826 710588
rect 137062 710352 137146 710588
rect 137382 710352 172826 710588
rect 173062 710352 173146 710588
rect 173382 710352 208826 710588
rect 209062 710352 209146 710588
rect 209382 710352 244826 710588
rect 245062 710352 245146 710588
rect 245382 710352 280826 710588
rect 281062 710352 281146 710588
rect 281382 710352 316826 710588
rect 317062 710352 317146 710588
rect 317382 710352 352826 710588
rect 353062 710352 353146 710588
rect 353382 710352 388826 710588
rect 389062 710352 389146 710588
rect 389382 710352 424826 710588
rect 425062 710352 425146 710588
rect 425382 710352 460826 710588
rect 461062 710352 461146 710588
rect 461382 710352 496826 710588
rect 497062 710352 497146 710588
rect 497382 710352 532826 710588
rect 533062 710352 533146 710588
rect 533382 710352 568826 710588
rect 569062 710352 569146 710588
rect 569382 710352 591412 710588
rect 591648 710352 591732 710588
rect 591968 710352 592000 710588
rect -8076 710320 592000 710352
rect -7116 709948 591040 709980
rect -7116 709712 -7084 709948
rect -6848 709712 -6764 709948
rect -6528 709712 24326 709948
rect 24562 709712 24646 709948
rect 24882 709712 60326 709948
rect 60562 709712 60646 709948
rect 60882 709712 96326 709948
rect 96562 709712 96646 709948
rect 96882 709712 132326 709948
rect 132562 709712 132646 709948
rect 132882 709712 168326 709948
rect 168562 709712 168646 709948
rect 168882 709712 204326 709948
rect 204562 709712 204646 709948
rect 204882 709712 240326 709948
rect 240562 709712 240646 709948
rect 240882 709712 276326 709948
rect 276562 709712 276646 709948
rect 276882 709712 312326 709948
rect 312562 709712 312646 709948
rect 312882 709712 348326 709948
rect 348562 709712 348646 709948
rect 348882 709712 384326 709948
rect 384562 709712 384646 709948
rect 384882 709712 420326 709948
rect 420562 709712 420646 709948
rect 420882 709712 456326 709948
rect 456562 709712 456646 709948
rect 456882 709712 492326 709948
rect 492562 709712 492646 709948
rect 492882 709712 528326 709948
rect 528562 709712 528646 709948
rect 528882 709712 564326 709948
rect 564562 709712 564646 709948
rect 564882 709712 590452 709948
rect 590688 709712 590772 709948
rect 591008 709712 591040 709948
rect -7116 709628 591040 709712
rect -7116 709392 -7084 709628
rect -6848 709392 -6764 709628
rect -6528 709392 24326 709628
rect 24562 709392 24646 709628
rect 24882 709392 60326 709628
rect 60562 709392 60646 709628
rect 60882 709392 96326 709628
rect 96562 709392 96646 709628
rect 96882 709392 132326 709628
rect 132562 709392 132646 709628
rect 132882 709392 168326 709628
rect 168562 709392 168646 709628
rect 168882 709392 204326 709628
rect 204562 709392 204646 709628
rect 204882 709392 240326 709628
rect 240562 709392 240646 709628
rect 240882 709392 276326 709628
rect 276562 709392 276646 709628
rect 276882 709392 312326 709628
rect 312562 709392 312646 709628
rect 312882 709392 348326 709628
rect 348562 709392 348646 709628
rect 348882 709392 384326 709628
rect 384562 709392 384646 709628
rect 384882 709392 420326 709628
rect 420562 709392 420646 709628
rect 420882 709392 456326 709628
rect 456562 709392 456646 709628
rect 456882 709392 492326 709628
rect 492562 709392 492646 709628
rect 492882 709392 528326 709628
rect 528562 709392 528646 709628
rect 528882 709392 564326 709628
rect 564562 709392 564646 709628
rect 564882 709392 590452 709628
rect 590688 709392 590772 709628
rect 591008 709392 591040 709628
rect -7116 709360 591040 709392
rect -6156 708988 590080 709020
rect -6156 708752 -6124 708988
rect -5888 708752 -5804 708988
rect -5568 708752 19826 708988
rect 20062 708752 20146 708988
rect 20382 708752 55826 708988
rect 56062 708752 56146 708988
rect 56382 708752 91826 708988
rect 92062 708752 92146 708988
rect 92382 708752 127826 708988
rect 128062 708752 128146 708988
rect 128382 708752 163826 708988
rect 164062 708752 164146 708988
rect 164382 708752 199826 708988
rect 200062 708752 200146 708988
rect 200382 708752 235826 708988
rect 236062 708752 236146 708988
rect 236382 708752 271826 708988
rect 272062 708752 272146 708988
rect 272382 708752 307826 708988
rect 308062 708752 308146 708988
rect 308382 708752 343826 708988
rect 344062 708752 344146 708988
rect 344382 708752 379826 708988
rect 380062 708752 380146 708988
rect 380382 708752 415826 708988
rect 416062 708752 416146 708988
rect 416382 708752 451826 708988
rect 452062 708752 452146 708988
rect 452382 708752 487826 708988
rect 488062 708752 488146 708988
rect 488382 708752 523826 708988
rect 524062 708752 524146 708988
rect 524382 708752 559826 708988
rect 560062 708752 560146 708988
rect 560382 708752 589492 708988
rect 589728 708752 589812 708988
rect 590048 708752 590080 708988
rect -6156 708668 590080 708752
rect -6156 708432 -6124 708668
rect -5888 708432 -5804 708668
rect -5568 708432 19826 708668
rect 20062 708432 20146 708668
rect 20382 708432 55826 708668
rect 56062 708432 56146 708668
rect 56382 708432 91826 708668
rect 92062 708432 92146 708668
rect 92382 708432 127826 708668
rect 128062 708432 128146 708668
rect 128382 708432 163826 708668
rect 164062 708432 164146 708668
rect 164382 708432 199826 708668
rect 200062 708432 200146 708668
rect 200382 708432 235826 708668
rect 236062 708432 236146 708668
rect 236382 708432 271826 708668
rect 272062 708432 272146 708668
rect 272382 708432 307826 708668
rect 308062 708432 308146 708668
rect 308382 708432 343826 708668
rect 344062 708432 344146 708668
rect 344382 708432 379826 708668
rect 380062 708432 380146 708668
rect 380382 708432 415826 708668
rect 416062 708432 416146 708668
rect 416382 708432 451826 708668
rect 452062 708432 452146 708668
rect 452382 708432 487826 708668
rect 488062 708432 488146 708668
rect 488382 708432 523826 708668
rect 524062 708432 524146 708668
rect 524382 708432 559826 708668
rect 560062 708432 560146 708668
rect 560382 708432 589492 708668
rect 589728 708432 589812 708668
rect 590048 708432 590080 708668
rect -6156 708400 590080 708432
rect -5196 708028 589120 708060
rect -5196 707792 -5164 708028
rect -4928 707792 -4844 708028
rect -4608 707792 15326 708028
rect 15562 707792 15646 708028
rect 15882 707792 51326 708028
rect 51562 707792 51646 708028
rect 51882 707792 87326 708028
rect 87562 707792 87646 708028
rect 87882 707792 123326 708028
rect 123562 707792 123646 708028
rect 123882 707792 159326 708028
rect 159562 707792 159646 708028
rect 159882 707792 195326 708028
rect 195562 707792 195646 708028
rect 195882 707792 231326 708028
rect 231562 707792 231646 708028
rect 231882 707792 267326 708028
rect 267562 707792 267646 708028
rect 267882 707792 303326 708028
rect 303562 707792 303646 708028
rect 303882 707792 339326 708028
rect 339562 707792 339646 708028
rect 339882 707792 375326 708028
rect 375562 707792 375646 708028
rect 375882 707792 411326 708028
rect 411562 707792 411646 708028
rect 411882 707792 447326 708028
rect 447562 707792 447646 708028
rect 447882 707792 483326 708028
rect 483562 707792 483646 708028
rect 483882 707792 519326 708028
rect 519562 707792 519646 708028
rect 519882 707792 555326 708028
rect 555562 707792 555646 708028
rect 555882 707792 588532 708028
rect 588768 707792 588852 708028
rect 589088 707792 589120 708028
rect -5196 707708 589120 707792
rect -5196 707472 -5164 707708
rect -4928 707472 -4844 707708
rect -4608 707472 15326 707708
rect 15562 707472 15646 707708
rect 15882 707472 51326 707708
rect 51562 707472 51646 707708
rect 51882 707472 87326 707708
rect 87562 707472 87646 707708
rect 87882 707472 123326 707708
rect 123562 707472 123646 707708
rect 123882 707472 159326 707708
rect 159562 707472 159646 707708
rect 159882 707472 195326 707708
rect 195562 707472 195646 707708
rect 195882 707472 231326 707708
rect 231562 707472 231646 707708
rect 231882 707472 267326 707708
rect 267562 707472 267646 707708
rect 267882 707472 303326 707708
rect 303562 707472 303646 707708
rect 303882 707472 339326 707708
rect 339562 707472 339646 707708
rect 339882 707472 375326 707708
rect 375562 707472 375646 707708
rect 375882 707472 411326 707708
rect 411562 707472 411646 707708
rect 411882 707472 447326 707708
rect 447562 707472 447646 707708
rect 447882 707472 483326 707708
rect 483562 707472 483646 707708
rect 483882 707472 519326 707708
rect 519562 707472 519646 707708
rect 519882 707472 555326 707708
rect 555562 707472 555646 707708
rect 555882 707472 588532 707708
rect 588768 707472 588852 707708
rect 589088 707472 589120 707708
rect -5196 707440 589120 707472
rect -4236 707068 588160 707100
rect -4236 706832 -4204 707068
rect -3968 706832 -3884 707068
rect -3648 706832 10826 707068
rect 11062 706832 11146 707068
rect 11382 706832 46826 707068
rect 47062 706832 47146 707068
rect 47382 706832 82826 707068
rect 83062 706832 83146 707068
rect 83382 706832 118826 707068
rect 119062 706832 119146 707068
rect 119382 706832 154826 707068
rect 155062 706832 155146 707068
rect 155382 706832 190826 707068
rect 191062 706832 191146 707068
rect 191382 706832 226826 707068
rect 227062 706832 227146 707068
rect 227382 706832 262826 707068
rect 263062 706832 263146 707068
rect 263382 706832 298826 707068
rect 299062 706832 299146 707068
rect 299382 706832 334826 707068
rect 335062 706832 335146 707068
rect 335382 706832 370826 707068
rect 371062 706832 371146 707068
rect 371382 706832 406826 707068
rect 407062 706832 407146 707068
rect 407382 706832 442826 707068
rect 443062 706832 443146 707068
rect 443382 706832 478826 707068
rect 479062 706832 479146 707068
rect 479382 706832 514826 707068
rect 515062 706832 515146 707068
rect 515382 706832 550826 707068
rect 551062 706832 551146 707068
rect 551382 706832 587572 707068
rect 587808 706832 587892 707068
rect 588128 706832 588160 707068
rect -4236 706748 588160 706832
rect -4236 706512 -4204 706748
rect -3968 706512 -3884 706748
rect -3648 706512 10826 706748
rect 11062 706512 11146 706748
rect 11382 706512 46826 706748
rect 47062 706512 47146 706748
rect 47382 706512 82826 706748
rect 83062 706512 83146 706748
rect 83382 706512 118826 706748
rect 119062 706512 119146 706748
rect 119382 706512 154826 706748
rect 155062 706512 155146 706748
rect 155382 706512 190826 706748
rect 191062 706512 191146 706748
rect 191382 706512 226826 706748
rect 227062 706512 227146 706748
rect 227382 706512 262826 706748
rect 263062 706512 263146 706748
rect 263382 706512 298826 706748
rect 299062 706512 299146 706748
rect 299382 706512 334826 706748
rect 335062 706512 335146 706748
rect 335382 706512 370826 706748
rect 371062 706512 371146 706748
rect 371382 706512 406826 706748
rect 407062 706512 407146 706748
rect 407382 706512 442826 706748
rect 443062 706512 443146 706748
rect 443382 706512 478826 706748
rect 479062 706512 479146 706748
rect 479382 706512 514826 706748
rect 515062 706512 515146 706748
rect 515382 706512 550826 706748
rect 551062 706512 551146 706748
rect 551382 706512 587572 706748
rect 587808 706512 587892 706748
rect 588128 706512 588160 706748
rect -4236 706480 588160 706512
rect -3276 706108 587200 706140
rect -3276 705872 -3244 706108
rect -3008 705872 -2924 706108
rect -2688 705872 6326 706108
rect 6562 705872 6646 706108
rect 6882 705872 42326 706108
rect 42562 705872 42646 706108
rect 42882 705872 78326 706108
rect 78562 705872 78646 706108
rect 78882 705872 114326 706108
rect 114562 705872 114646 706108
rect 114882 705872 150326 706108
rect 150562 705872 150646 706108
rect 150882 705872 186326 706108
rect 186562 705872 186646 706108
rect 186882 705872 222326 706108
rect 222562 705872 222646 706108
rect 222882 705872 258326 706108
rect 258562 705872 258646 706108
rect 258882 705872 294326 706108
rect 294562 705872 294646 706108
rect 294882 705872 330326 706108
rect 330562 705872 330646 706108
rect 330882 705872 366326 706108
rect 366562 705872 366646 706108
rect 366882 705872 402326 706108
rect 402562 705872 402646 706108
rect 402882 705872 438326 706108
rect 438562 705872 438646 706108
rect 438882 705872 474326 706108
rect 474562 705872 474646 706108
rect 474882 705872 510326 706108
rect 510562 705872 510646 706108
rect 510882 705872 546326 706108
rect 546562 705872 546646 706108
rect 546882 705872 582326 706108
rect 582562 705872 582646 706108
rect 582882 705872 586612 706108
rect 586848 705872 586932 706108
rect 587168 705872 587200 706108
rect -3276 705788 587200 705872
rect -3276 705552 -3244 705788
rect -3008 705552 -2924 705788
rect -2688 705552 6326 705788
rect 6562 705552 6646 705788
rect 6882 705552 42326 705788
rect 42562 705552 42646 705788
rect 42882 705552 78326 705788
rect 78562 705552 78646 705788
rect 78882 705552 114326 705788
rect 114562 705552 114646 705788
rect 114882 705552 150326 705788
rect 150562 705552 150646 705788
rect 150882 705552 186326 705788
rect 186562 705552 186646 705788
rect 186882 705552 222326 705788
rect 222562 705552 222646 705788
rect 222882 705552 258326 705788
rect 258562 705552 258646 705788
rect 258882 705552 294326 705788
rect 294562 705552 294646 705788
rect 294882 705552 330326 705788
rect 330562 705552 330646 705788
rect 330882 705552 366326 705788
rect 366562 705552 366646 705788
rect 366882 705552 402326 705788
rect 402562 705552 402646 705788
rect 402882 705552 438326 705788
rect 438562 705552 438646 705788
rect 438882 705552 474326 705788
rect 474562 705552 474646 705788
rect 474882 705552 510326 705788
rect 510562 705552 510646 705788
rect 510882 705552 546326 705788
rect 546562 705552 546646 705788
rect 546882 705552 582326 705788
rect 582562 705552 582646 705788
rect 582882 705552 586612 705788
rect 586848 705552 586932 705788
rect 587168 705552 587200 705788
rect -3276 705520 587200 705552
rect -2316 705148 586240 705180
rect -2316 704912 -2284 705148
rect -2048 704912 -1964 705148
rect -1728 704912 1826 705148
rect 2062 704912 2146 705148
rect 2382 704912 37826 705148
rect 38062 704912 38146 705148
rect 38382 704912 73826 705148
rect 74062 704912 74146 705148
rect 74382 704912 109826 705148
rect 110062 704912 110146 705148
rect 110382 704912 145826 705148
rect 146062 704912 146146 705148
rect 146382 704912 181826 705148
rect 182062 704912 182146 705148
rect 182382 704912 217826 705148
rect 218062 704912 218146 705148
rect 218382 704912 253826 705148
rect 254062 704912 254146 705148
rect 254382 704912 289826 705148
rect 290062 704912 290146 705148
rect 290382 704912 325826 705148
rect 326062 704912 326146 705148
rect 326382 704912 361826 705148
rect 362062 704912 362146 705148
rect 362382 704912 397826 705148
rect 398062 704912 398146 705148
rect 398382 704912 433826 705148
rect 434062 704912 434146 705148
rect 434382 704912 469826 705148
rect 470062 704912 470146 705148
rect 470382 704912 505826 705148
rect 506062 704912 506146 705148
rect 506382 704912 541826 705148
rect 542062 704912 542146 705148
rect 542382 704912 577826 705148
rect 578062 704912 578146 705148
rect 578382 704912 585652 705148
rect 585888 704912 585972 705148
rect 586208 704912 586240 705148
rect -2316 704828 586240 704912
rect -2316 704592 -2284 704828
rect -2048 704592 -1964 704828
rect -1728 704592 1826 704828
rect 2062 704592 2146 704828
rect 2382 704592 37826 704828
rect 38062 704592 38146 704828
rect 38382 704592 73826 704828
rect 74062 704592 74146 704828
rect 74382 704592 109826 704828
rect 110062 704592 110146 704828
rect 110382 704592 145826 704828
rect 146062 704592 146146 704828
rect 146382 704592 181826 704828
rect 182062 704592 182146 704828
rect 182382 704592 217826 704828
rect 218062 704592 218146 704828
rect 218382 704592 253826 704828
rect 254062 704592 254146 704828
rect 254382 704592 289826 704828
rect 290062 704592 290146 704828
rect 290382 704592 325826 704828
rect 326062 704592 326146 704828
rect 326382 704592 361826 704828
rect 362062 704592 362146 704828
rect 362382 704592 397826 704828
rect 398062 704592 398146 704828
rect 398382 704592 433826 704828
rect 434062 704592 434146 704828
rect 434382 704592 469826 704828
rect 470062 704592 470146 704828
rect 470382 704592 505826 704828
rect 506062 704592 506146 704828
rect 506382 704592 541826 704828
rect 542062 704592 542146 704828
rect 542382 704592 577826 704828
rect 578062 704592 578146 704828
rect 578382 704592 585652 704828
rect 585888 704592 585972 704828
rect 586208 704592 586240 704828
rect -2316 704560 586240 704592
rect -9036 700954 592960 700986
rect -9036 700718 -5164 700954
rect -4928 700718 -4844 700954
rect -4608 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588532 700954
rect 588768 700718 588852 700954
rect 589088 700718 592960 700954
rect -9036 700634 592960 700718
rect -9036 700398 -5164 700634
rect -4928 700398 -4844 700634
rect -4608 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588532 700634
rect 588768 700398 588852 700634
rect 589088 700398 592960 700634
rect -9036 700366 592960 700398
rect -9036 696454 592960 696486
rect -9036 696218 -4204 696454
rect -3968 696218 -3884 696454
rect -3648 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587572 696454
rect 587808 696218 587892 696454
rect 588128 696218 592960 696454
rect -9036 696134 592960 696218
rect -9036 695898 -4204 696134
rect -3968 695898 -3884 696134
rect -3648 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587572 696134
rect 587808 695898 587892 696134
rect 588128 695898 592960 696134
rect -9036 695866 592960 695898
rect -9036 691954 592960 691986
rect -9036 691718 -3244 691954
rect -3008 691718 -2924 691954
rect -2688 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586612 691954
rect 586848 691718 586932 691954
rect 587168 691718 592960 691954
rect -9036 691634 592960 691718
rect -9036 691398 -3244 691634
rect -3008 691398 -2924 691634
rect -2688 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586612 691634
rect 586848 691398 586932 691634
rect 587168 691398 592960 691634
rect -9036 691366 592960 691398
rect -9036 687454 592960 687486
rect -9036 687218 -2284 687454
rect -2048 687218 -1964 687454
rect -1728 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585652 687454
rect 585888 687218 585972 687454
rect 586208 687218 592960 687454
rect -9036 687134 592960 687218
rect -9036 686898 -2284 687134
rect -2048 686898 -1964 687134
rect -1728 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585652 687134
rect 585888 686898 585972 687134
rect 586208 686898 592960 687134
rect -9036 686866 592960 686898
rect -9036 682954 592960 682986
rect -9036 682718 -9004 682954
rect -8768 682718 -8684 682954
rect -8448 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592372 682954
rect 592608 682718 592692 682954
rect 592928 682718 592960 682954
rect -9036 682634 592960 682718
rect -9036 682398 -9004 682634
rect -8768 682398 -8684 682634
rect -8448 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592372 682634
rect 592608 682398 592692 682634
rect 592928 682398 592960 682634
rect -9036 682366 592960 682398
rect -9036 678454 592960 678486
rect -9036 678218 -8044 678454
rect -7808 678218 -7724 678454
rect -7488 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591412 678454
rect 591648 678218 591732 678454
rect 591968 678218 592960 678454
rect -9036 678134 592960 678218
rect -9036 677898 -8044 678134
rect -7808 677898 -7724 678134
rect -7488 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591412 678134
rect 591648 677898 591732 678134
rect 591968 677898 592960 678134
rect -9036 677866 592960 677898
rect -9036 673954 592960 673986
rect -9036 673718 -7084 673954
rect -6848 673718 -6764 673954
rect -6528 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590452 673954
rect 590688 673718 590772 673954
rect 591008 673718 592960 673954
rect -9036 673634 592960 673718
rect -9036 673398 -7084 673634
rect -6848 673398 -6764 673634
rect -6528 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590452 673634
rect 590688 673398 590772 673634
rect 591008 673398 592960 673634
rect -9036 673366 592960 673398
rect -9036 669454 592960 669486
rect -9036 669218 -6124 669454
rect -5888 669218 -5804 669454
rect -5568 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589492 669454
rect 589728 669218 589812 669454
rect 590048 669218 592960 669454
rect -9036 669134 592960 669218
rect -9036 668898 -6124 669134
rect -5888 668898 -5804 669134
rect -5568 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589492 669134
rect 589728 668898 589812 669134
rect 590048 668898 592960 669134
rect -9036 668866 592960 668898
rect -9036 664954 592960 664986
rect -9036 664718 -5164 664954
rect -4928 664718 -4844 664954
rect -4608 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588532 664954
rect 588768 664718 588852 664954
rect 589088 664718 592960 664954
rect -9036 664634 592960 664718
rect -9036 664398 -5164 664634
rect -4928 664398 -4844 664634
rect -4608 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588532 664634
rect 588768 664398 588852 664634
rect 589088 664398 592960 664634
rect -9036 664366 592960 664398
rect -9036 660454 592960 660486
rect -9036 660218 -4204 660454
rect -3968 660218 -3884 660454
rect -3648 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587572 660454
rect 587808 660218 587892 660454
rect 588128 660218 592960 660454
rect -9036 660134 592960 660218
rect -9036 659898 -4204 660134
rect -3968 659898 -3884 660134
rect -3648 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587572 660134
rect 587808 659898 587892 660134
rect 588128 659898 592960 660134
rect -9036 659866 592960 659898
rect -9036 655954 592960 655986
rect -9036 655718 -3244 655954
rect -3008 655718 -2924 655954
rect -2688 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586612 655954
rect 586848 655718 586932 655954
rect 587168 655718 592960 655954
rect -9036 655634 592960 655718
rect -9036 655398 -3244 655634
rect -3008 655398 -2924 655634
rect -2688 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586612 655634
rect 586848 655398 586932 655634
rect 587168 655398 592960 655634
rect -9036 655366 592960 655398
rect -9036 651454 592960 651486
rect -9036 651218 -2284 651454
rect -2048 651218 -1964 651454
rect -1728 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585652 651454
rect 585888 651218 585972 651454
rect 586208 651218 592960 651454
rect -9036 651134 592960 651218
rect -9036 650898 -2284 651134
rect -2048 650898 -1964 651134
rect -1728 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585652 651134
rect 585888 650898 585972 651134
rect 586208 650898 592960 651134
rect -9036 650866 592960 650898
rect -9036 646954 592960 646986
rect -9036 646718 -9004 646954
rect -8768 646718 -8684 646954
rect -8448 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592372 646954
rect 592608 646718 592692 646954
rect 592928 646718 592960 646954
rect -9036 646634 592960 646718
rect -9036 646398 -9004 646634
rect -8768 646398 -8684 646634
rect -8448 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592372 646634
rect 592608 646398 592692 646634
rect 592928 646398 592960 646634
rect -9036 646366 592960 646398
rect -9036 642454 592960 642486
rect -9036 642218 -8044 642454
rect -7808 642218 -7724 642454
rect -7488 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591412 642454
rect 591648 642218 591732 642454
rect 591968 642218 592960 642454
rect -9036 642134 592960 642218
rect -9036 641898 -8044 642134
rect -7808 641898 -7724 642134
rect -7488 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591412 642134
rect 591648 641898 591732 642134
rect 591968 641898 592960 642134
rect -9036 641866 592960 641898
rect -9036 637954 592960 637986
rect -9036 637718 -7084 637954
rect -6848 637718 -6764 637954
rect -6528 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590452 637954
rect 590688 637718 590772 637954
rect 591008 637718 592960 637954
rect -9036 637634 592960 637718
rect -9036 637398 -7084 637634
rect -6848 637398 -6764 637634
rect -6528 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590452 637634
rect 590688 637398 590772 637634
rect 591008 637398 592960 637634
rect -9036 637366 592960 637398
rect -9036 633454 592960 633486
rect -9036 633218 -6124 633454
rect -5888 633218 -5804 633454
rect -5568 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589492 633454
rect 589728 633218 589812 633454
rect 590048 633218 592960 633454
rect -9036 633134 592960 633218
rect -9036 632898 -6124 633134
rect -5888 632898 -5804 633134
rect -5568 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589492 633134
rect 589728 632898 589812 633134
rect 590048 632898 592960 633134
rect -9036 632866 592960 632898
rect -9036 628954 592960 628986
rect -9036 628718 -5164 628954
rect -4928 628718 -4844 628954
rect -4608 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588532 628954
rect 588768 628718 588852 628954
rect 589088 628718 592960 628954
rect -9036 628634 592960 628718
rect -9036 628398 -5164 628634
rect -4928 628398 -4844 628634
rect -4608 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588532 628634
rect 588768 628398 588852 628634
rect 589088 628398 592960 628634
rect -9036 628366 592960 628398
rect -9036 624454 592960 624486
rect -9036 624218 -4204 624454
rect -3968 624218 -3884 624454
rect -3648 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587572 624454
rect 587808 624218 587892 624454
rect 588128 624218 592960 624454
rect -9036 624134 592960 624218
rect -9036 623898 -4204 624134
rect -3968 623898 -3884 624134
rect -3648 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587572 624134
rect 587808 623898 587892 624134
rect 588128 623898 592960 624134
rect -9036 623866 592960 623898
rect -9036 619954 592960 619986
rect -9036 619718 -3244 619954
rect -3008 619718 -2924 619954
rect -2688 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586612 619954
rect 586848 619718 586932 619954
rect 587168 619718 592960 619954
rect -9036 619634 592960 619718
rect -9036 619398 -3244 619634
rect -3008 619398 -2924 619634
rect -2688 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586612 619634
rect 586848 619398 586932 619634
rect 587168 619398 592960 619634
rect -9036 619366 592960 619398
rect -9036 615454 592960 615486
rect -9036 615218 -2284 615454
rect -2048 615218 -1964 615454
rect -1728 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585652 615454
rect 585888 615218 585972 615454
rect 586208 615218 592960 615454
rect -9036 615134 592960 615218
rect -9036 614898 -2284 615134
rect -2048 614898 -1964 615134
rect -1728 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585652 615134
rect 585888 614898 585972 615134
rect 586208 614898 592960 615134
rect -9036 614866 592960 614898
rect -9036 610954 592960 610986
rect -9036 610718 -9004 610954
rect -8768 610718 -8684 610954
rect -8448 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592372 610954
rect 592608 610718 592692 610954
rect 592928 610718 592960 610954
rect -9036 610634 592960 610718
rect -9036 610398 -9004 610634
rect -8768 610398 -8684 610634
rect -8448 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592372 610634
rect 592608 610398 592692 610634
rect 592928 610398 592960 610634
rect -9036 610366 592960 610398
rect -9036 606454 592960 606486
rect -9036 606218 -8044 606454
rect -7808 606218 -7724 606454
rect -7488 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591412 606454
rect 591648 606218 591732 606454
rect 591968 606218 592960 606454
rect -9036 606134 592960 606218
rect -9036 605898 -8044 606134
rect -7808 605898 -7724 606134
rect -7488 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591412 606134
rect 591648 605898 591732 606134
rect 591968 605898 592960 606134
rect -9036 605866 592960 605898
rect -9036 601954 592960 601986
rect -9036 601718 -7084 601954
rect -6848 601718 -6764 601954
rect -6528 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590452 601954
rect 590688 601718 590772 601954
rect 591008 601718 592960 601954
rect -9036 601634 592960 601718
rect -9036 601398 -7084 601634
rect -6848 601398 -6764 601634
rect -6528 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590452 601634
rect 590688 601398 590772 601634
rect 591008 601398 592960 601634
rect -9036 601366 592960 601398
rect -9036 597454 592960 597486
rect -9036 597218 -6124 597454
rect -5888 597218 -5804 597454
rect -5568 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589492 597454
rect 589728 597218 589812 597454
rect 590048 597218 592960 597454
rect -9036 597134 592960 597218
rect -9036 596898 -6124 597134
rect -5888 596898 -5804 597134
rect -5568 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589492 597134
rect 589728 596898 589812 597134
rect 590048 596898 592960 597134
rect -9036 596866 592960 596898
rect -9036 592954 592960 592986
rect -9036 592718 -5164 592954
rect -4928 592718 -4844 592954
rect -4608 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588532 592954
rect 588768 592718 588852 592954
rect 589088 592718 592960 592954
rect -9036 592634 592960 592718
rect -9036 592398 -5164 592634
rect -4928 592398 -4844 592634
rect -4608 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588532 592634
rect 588768 592398 588852 592634
rect 589088 592398 592960 592634
rect -9036 592366 592960 592398
rect -9036 588454 592960 588486
rect -9036 588218 -4204 588454
rect -3968 588218 -3884 588454
rect -3648 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587572 588454
rect 587808 588218 587892 588454
rect 588128 588218 592960 588454
rect -9036 588134 592960 588218
rect -9036 587898 -4204 588134
rect -3968 587898 -3884 588134
rect -3648 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587572 588134
rect 587808 587898 587892 588134
rect 588128 587898 592960 588134
rect -9036 587866 592960 587898
rect -9036 583954 592960 583986
rect -9036 583718 -3244 583954
rect -3008 583718 -2924 583954
rect -2688 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586612 583954
rect 586848 583718 586932 583954
rect 587168 583718 592960 583954
rect -9036 583634 592960 583718
rect -9036 583398 -3244 583634
rect -3008 583398 -2924 583634
rect -2688 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586612 583634
rect 586848 583398 586932 583634
rect 587168 583398 592960 583634
rect -9036 583366 592960 583398
rect -9036 579454 592960 579486
rect -9036 579218 -2284 579454
rect -2048 579218 -1964 579454
rect -1728 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585652 579454
rect 585888 579218 585972 579454
rect 586208 579218 592960 579454
rect -9036 579134 592960 579218
rect -9036 578898 -2284 579134
rect -2048 578898 -1964 579134
rect -1728 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585652 579134
rect 585888 578898 585972 579134
rect 586208 578898 592960 579134
rect -9036 578866 592960 578898
rect -9036 574954 592960 574986
rect -9036 574718 -9004 574954
rect -8768 574718 -8684 574954
rect -8448 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592372 574954
rect 592608 574718 592692 574954
rect 592928 574718 592960 574954
rect -9036 574634 592960 574718
rect -9036 574398 -9004 574634
rect -8768 574398 -8684 574634
rect -8448 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592372 574634
rect 592608 574398 592692 574634
rect 592928 574398 592960 574634
rect -9036 574366 592960 574398
rect -9036 570454 592960 570486
rect -9036 570218 -8044 570454
rect -7808 570218 -7724 570454
rect -7488 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591412 570454
rect 591648 570218 591732 570454
rect 591968 570218 592960 570454
rect -9036 570134 592960 570218
rect -9036 569898 -8044 570134
rect -7808 569898 -7724 570134
rect -7488 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591412 570134
rect 591648 569898 591732 570134
rect 591968 569898 592960 570134
rect -9036 569866 592960 569898
rect -9036 565954 592960 565986
rect -9036 565718 -7084 565954
rect -6848 565718 -6764 565954
rect -6528 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590452 565954
rect 590688 565718 590772 565954
rect 591008 565718 592960 565954
rect -9036 565634 592960 565718
rect -9036 565398 -7084 565634
rect -6848 565398 -6764 565634
rect -6528 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590452 565634
rect 590688 565398 590772 565634
rect 591008 565398 592960 565634
rect -9036 565366 592960 565398
rect -9036 561454 592960 561486
rect -9036 561218 -6124 561454
rect -5888 561218 -5804 561454
rect -5568 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589492 561454
rect 589728 561218 589812 561454
rect 590048 561218 592960 561454
rect -9036 561134 592960 561218
rect -9036 560898 -6124 561134
rect -5888 560898 -5804 561134
rect -5568 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589492 561134
rect 589728 560898 589812 561134
rect 590048 560898 592960 561134
rect -9036 560866 592960 560898
rect -9036 556954 592960 556986
rect -9036 556718 -5164 556954
rect -4928 556718 -4844 556954
rect -4608 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588532 556954
rect 588768 556718 588852 556954
rect 589088 556718 592960 556954
rect -9036 556634 592960 556718
rect -9036 556398 -5164 556634
rect -4928 556398 -4844 556634
rect -4608 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588532 556634
rect 588768 556398 588852 556634
rect 589088 556398 592960 556634
rect -9036 556366 592960 556398
rect -9036 552454 592960 552486
rect -9036 552218 -4204 552454
rect -3968 552218 -3884 552454
rect -3648 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587572 552454
rect 587808 552218 587892 552454
rect 588128 552218 592960 552454
rect -9036 552134 592960 552218
rect -9036 551898 -4204 552134
rect -3968 551898 -3884 552134
rect -3648 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587572 552134
rect 587808 551898 587892 552134
rect 588128 551898 592960 552134
rect -9036 551866 592960 551898
rect -9036 547954 592960 547986
rect -9036 547718 -3244 547954
rect -3008 547718 -2924 547954
rect -2688 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 220328 547954
rect 220564 547718 356056 547954
rect 356292 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586612 547954
rect 586848 547718 586932 547954
rect 587168 547718 592960 547954
rect -9036 547634 592960 547718
rect -9036 547398 -3244 547634
rect -3008 547398 -2924 547634
rect -2688 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 220328 547634
rect 220564 547398 356056 547634
rect 356292 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586612 547634
rect 586848 547398 586932 547634
rect 587168 547398 592960 547634
rect -9036 547366 592960 547398
rect -9036 543454 592960 543486
rect -9036 543218 -2284 543454
rect -2048 543218 -1964 543454
rect -1728 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 221008 543454
rect 221244 543218 355376 543454
rect 355612 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585652 543454
rect 585888 543218 585972 543454
rect 586208 543218 592960 543454
rect -9036 543134 592960 543218
rect -9036 542898 -2284 543134
rect -2048 542898 -1964 543134
rect -1728 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 221008 543134
rect 221244 542898 355376 543134
rect 355612 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585652 543134
rect 585888 542898 585972 543134
rect 586208 542898 592960 543134
rect -9036 542866 592960 542898
rect -9036 538954 592960 538986
rect -9036 538718 -9004 538954
rect -8768 538718 -8684 538954
rect -8448 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592372 538954
rect 592608 538718 592692 538954
rect 592928 538718 592960 538954
rect -9036 538634 592960 538718
rect -9036 538398 -9004 538634
rect -8768 538398 -8684 538634
rect -8448 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592372 538634
rect 592608 538398 592692 538634
rect 592928 538398 592960 538634
rect -9036 538366 592960 538398
rect -9036 534454 592960 534486
rect -9036 534218 -8044 534454
rect -7808 534218 -7724 534454
rect -7488 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591412 534454
rect 591648 534218 591732 534454
rect 591968 534218 592960 534454
rect -9036 534134 592960 534218
rect -9036 533898 -8044 534134
rect -7808 533898 -7724 534134
rect -7488 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591412 534134
rect 591648 533898 591732 534134
rect 591968 533898 592960 534134
rect -9036 533866 592960 533898
rect -9036 529954 592960 529986
rect -9036 529718 -7084 529954
rect -6848 529718 -6764 529954
rect -6528 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590452 529954
rect 590688 529718 590772 529954
rect 591008 529718 592960 529954
rect -9036 529634 592960 529718
rect -9036 529398 -7084 529634
rect -6848 529398 -6764 529634
rect -6528 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590452 529634
rect 590688 529398 590772 529634
rect 591008 529398 592960 529634
rect -9036 529366 592960 529398
rect -9036 525454 592960 525486
rect -9036 525218 -6124 525454
rect -5888 525218 -5804 525454
rect -5568 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589492 525454
rect 589728 525218 589812 525454
rect 590048 525218 592960 525454
rect -9036 525134 592960 525218
rect -9036 524898 -6124 525134
rect -5888 524898 -5804 525134
rect -5568 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589492 525134
rect 589728 524898 589812 525134
rect 590048 524898 592960 525134
rect -9036 524866 592960 524898
rect -9036 520954 592960 520986
rect -9036 520718 -5164 520954
rect -4928 520718 -4844 520954
rect -4608 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588532 520954
rect 588768 520718 588852 520954
rect 589088 520718 592960 520954
rect -9036 520634 592960 520718
rect -9036 520398 -5164 520634
rect -4928 520398 -4844 520634
rect -4608 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588532 520634
rect 588768 520398 588852 520634
rect 589088 520398 592960 520634
rect -9036 520366 592960 520398
rect -9036 516454 592960 516486
rect -9036 516218 -4204 516454
rect -3968 516218 -3884 516454
rect -3648 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587572 516454
rect 587808 516218 587892 516454
rect 588128 516218 592960 516454
rect -9036 516134 592960 516218
rect -9036 515898 -4204 516134
rect -3968 515898 -3884 516134
rect -3648 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587572 516134
rect 587808 515898 587892 516134
rect 588128 515898 592960 516134
rect -9036 515866 592960 515898
rect -9036 511954 592960 511986
rect -9036 511718 -3244 511954
rect -3008 511718 -2924 511954
rect -2688 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 220328 511954
rect 220564 511718 356056 511954
rect 356292 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586612 511954
rect 586848 511718 586932 511954
rect 587168 511718 592960 511954
rect -9036 511634 592960 511718
rect -9036 511398 -3244 511634
rect -3008 511398 -2924 511634
rect -2688 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 220328 511634
rect 220564 511398 356056 511634
rect 356292 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586612 511634
rect 586848 511398 586932 511634
rect 587168 511398 592960 511634
rect -9036 511366 592960 511398
rect -9036 507454 592960 507486
rect -9036 507218 -2284 507454
rect -2048 507218 -1964 507454
rect -1728 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 221008 507454
rect 221244 507218 355376 507454
rect 355612 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585652 507454
rect 585888 507218 585972 507454
rect 586208 507218 592960 507454
rect -9036 507134 592960 507218
rect -9036 506898 -2284 507134
rect -2048 506898 -1964 507134
rect -1728 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 221008 507134
rect 221244 506898 355376 507134
rect 355612 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585652 507134
rect 585888 506898 585972 507134
rect 586208 506898 592960 507134
rect -9036 506866 592960 506898
rect -9036 502954 592960 502986
rect -9036 502718 -9004 502954
rect -8768 502718 -8684 502954
rect -8448 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592372 502954
rect 592608 502718 592692 502954
rect 592928 502718 592960 502954
rect -9036 502634 592960 502718
rect -9036 502398 -9004 502634
rect -8768 502398 -8684 502634
rect -8448 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592372 502634
rect 592608 502398 592692 502634
rect 592928 502398 592960 502634
rect -9036 502366 592960 502398
rect -9036 498454 592960 498486
rect -9036 498218 -8044 498454
rect -7808 498218 -7724 498454
rect -7488 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591412 498454
rect 591648 498218 591732 498454
rect 591968 498218 592960 498454
rect -9036 498134 592960 498218
rect -9036 497898 -8044 498134
rect -7808 497898 -7724 498134
rect -7488 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591412 498134
rect 591648 497898 591732 498134
rect 591968 497898 592960 498134
rect -9036 497866 592960 497898
rect -9036 493954 592960 493986
rect -9036 493718 -7084 493954
rect -6848 493718 -6764 493954
rect -6528 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590452 493954
rect 590688 493718 590772 493954
rect 591008 493718 592960 493954
rect -9036 493634 592960 493718
rect -9036 493398 -7084 493634
rect -6848 493398 -6764 493634
rect -6528 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590452 493634
rect 590688 493398 590772 493634
rect 591008 493398 592960 493634
rect -9036 493366 592960 493398
rect -9036 489454 592960 489486
rect -9036 489218 -6124 489454
rect -5888 489218 -5804 489454
rect -5568 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589492 489454
rect 589728 489218 589812 489454
rect 590048 489218 592960 489454
rect -9036 489134 592960 489218
rect -9036 488898 -6124 489134
rect -5888 488898 -5804 489134
rect -5568 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589492 489134
rect 589728 488898 589812 489134
rect 590048 488898 592960 489134
rect -9036 488866 592960 488898
rect -9036 484954 592960 484986
rect -9036 484718 -5164 484954
rect -4928 484718 -4844 484954
rect -4608 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588532 484954
rect 588768 484718 588852 484954
rect 589088 484718 592960 484954
rect -9036 484634 592960 484718
rect -9036 484398 -5164 484634
rect -4928 484398 -4844 484634
rect -4608 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588532 484634
rect 588768 484398 588852 484634
rect 589088 484398 592960 484634
rect -9036 484366 592960 484398
rect -9036 480454 592960 480486
rect -9036 480218 -4204 480454
rect -3968 480218 -3884 480454
rect -3648 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587572 480454
rect 587808 480218 587892 480454
rect 588128 480218 592960 480454
rect -9036 480134 592960 480218
rect -9036 479898 -4204 480134
rect -3968 479898 -3884 480134
rect -3648 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587572 480134
rect 587808 479898 587892 480134
rect 588128 479898 592960 480134
rect -9036 479866 592960 479898
rect -9036 475954 592960 475986
rect -9036 475718 -3244 475954
rect -3008 475718 -2924 475954
rect -2688 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586612 475954
rect 586848 475718 586932 475954
rect 587168 475718 592960 475954
rect -9036 475634 592960 475718
rect -9036 475398 -3244 475634
rect -3008 475398 -2924 475634
rect -2688 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586612 475634
rect 586848 475398 586932 475634
rect 587168 475398 592960 475634
rect -9036 475366 592960 475398
rect -9036 471454 592960 471486
rect -9036 471218 -2284 471454
rect -2048 471218 -1964 471454
rect -1728 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585652 471454
rect 585888 471218 585972 471454
rect 586208 471218 592960 471454
rect -9036 471134 592960 471218
rect -9036 470898 -2284 471134
rect -2048 470898 -1964 471134
rect -1728 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585652 471134
rect 585888 470898 585972 471134
rect 586208 470898 592960 471134
rect -9036 470866 592960 470898
rect -9036 466954 592960 466986
rect -9036 466718 -9004 466954
rect -8768 466718 -8684 466954
rect -8448 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592372 466954
rect 592608 466718 592692 466954
rect 592928 466718 592960 466954
rect -9036 466634 592960 466718
rect -9036 466398 -9004 466634
rect -8768 466398 -8684 466634
rect -8448 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592372 466634
rect 592608 466398 592692 466634
rect 592928 466398 592960 466634
rect -9036 466366 592960 466398
rect -9036 462454 592960 462486
rect -9036 462218 -8044 462454
rect -7808 462218 -7724 462454
rect -7488 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591412 462454
rect 591648 462218 591732 462454
rect 591968 462218 592960 462454
rect -9036 462134 592960 462218
rect -9036 461898 -8044 462134
rect -7808 461898 -7724 462134
rect -7488 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591412 462134
rect 591648 461898 591732 462134
rect 591968 461898 592960 462134
rect -9036 461866 592960 461898
rect -9036 457954 592960 457986
rect -9036 457718 -7084 457954
rect -6848 457718 -6764 457954
rect -6528 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590452 457954
rect 590688 457718 590772 457954
rect 591008 457718 592960 457954
rect -9036 457634 592960 457718
rect -9036 457398 -7084 457634
rect -6848 457398 -6764 457634
rect -6528 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590452 457634
rect 590688 457398 590772 457634
rect 591008 457398 592960 457634
rect -9036 457366 592960 457398
rect -9036 453454 592960 453486
rect -9036 453218 -6124 453454
rect -5888 453218 -5804 453454
rect -5568 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589492 453454
rect 589728 453218 589812 453454
rect 590048 453218 592960 453454
rect -9036 453134 592960 453218
rect -9036 452898 -6124 453134
rect -5888 452898 -5804 453134
rect -5568 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589492 453134
rect 589728 452898 589812 453134
rect 590048 452898 592960 453134
rect -9036 452866 592960 452898
rect -9036 448954 592960 448986
rect -9036 448718 -5164 448954
rect -4928 448718 -4844 448954
rect -4608 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588532 448954
rect 588768 448718 588852 448954
rect 589088 448718 592960 448954
rect -9036 448634 592960 448718
rect -9036 448398 -5164 448634
rect -4928 448398 -4844 448634
rect -4608 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588532 448634
rect 588768 448398 588852 448634
rect 589088 448398 592960 448634
rect -9036 448366 592960 448398
rect -9036 444454 592960 444486
rect -9036 444218 -4204 444454
rect -3968 444218 -3884 444454
rect -3648 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587572 444454
rect 587808 444218 587892 444454
rect 588128 444218 592960 444454
rect -9036 444134 592960 444218
rect -9036 443898 -4204 444134
rect -3968 443898 -3884 444134
rect -3648 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587572 444134
rect 587808 443898 587892 444134
rect 588128 443898 592960 444134
rect -9036 443866 592960 443898
rect -9036 439954 592960 439986
rect -9036 439718 -3244 439954
rect -3008 439718 -2924 439954
rect -2688 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586612 439954
rect 586848 439718 586932 439954
rect 587168 439718 592960 439954
rect -9036 439634 592960 439718
rect -9036 439398 -3244 439634
rect -3008 439398 -2924 439634
rect -2688 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586612 439634
rect 586848 439398 586932 439634
rect 587168 439398 592960 439634
rect -9036 439366 592960 439398
rect -9036 435454 592960 435486
rect -9036 435218 -2284 435454
rect -2048 435218 -1964 435454
rect -1728 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585652 435454
rect 585888 435218 585972 435454
rect 586208 435218 592960 435454
rect -9036 435134 592960 435218
rect -9036 434898 -2284 435134
rect -2048 434898 -1964 435134
rect -1728 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585652 435134
rect 585888 434898 585972 435134
rect 586208 434898 592960 435134
rect -9036 434866 592960 434898
rect -9036 430954 592960 430986
rect -9036 430718 -9004 430954
rect -8768 430718 -8684 430954
rect -8448 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592372 430954
rect 592608 430718 592692 430954
rect 592928 430718 592960 430954
rect -9036 430634 592960 430718
rect -9036 430398 -9004 430634
rect -8768 430398 -8684 430634
rect -8448 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592372 430634
rect 592608 430398 592692 430634
rect 592928 430398 592960 430634
rect -9036 430366 592960 430398
rect -9036 426454 592960 426486
rect -9036 426218 -8044 426454
rect -7808 426218 -7724 426454
rect -7488 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591412 426454
rect 591648 426218 591732 426454
rect 591968 426218 592960 426454
rect -9036 426134 592960 426218
rect -9036 425898 -8044 426134
rect -7808 425898 -7724 426134
rect -7488 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591412 426134
rect 591648 425898 591732 426134
rect 591968 425898 592960 426134
rect -9036 425866 592960 425898
rect -9036 421954 592960 421986
rect -9036 421718 -7084 421954
rect -6848 421718 -6764 421954
rect -6528 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590452 421954
rect 590688 421718 590772 421954
rect 591008 421718 592960 421954
rect -9036 421634 592960 421718
rect -9036 421398 -7084 421634
rect -6848 421398 -6764 421634
rect -6528 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590452 421634
rect 590688 421398 590772 421634
rect 591008 421398 592960 421634
rect -9036 421366 592960 421398
rect -9036 417454 592960 417486
rect -9036 417218 -6124 417454
rect -5888 417218 -5804 417454
rect -5568 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589492 417454
rect 589728 417218 589812 417454
rect 590048 417218 592960 417454
rect -9036 417134 592960 417218
rect -9036 416898 -6124 417134
rect -5888 416898 -5804 417134
rect -5568 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589492 417134
rect 589728 416898 589812 417134
rect 590048 416898 592960 417134
rect -9036 416866 592960 416898
rect -9036 412954 592960 412986
rect -9036 412718 -5164 412954
rect -4928 412718 -4844 412954
rect -4608 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588532 412954
rect 588768 412718 588852 412954
rect 589088 412718 592960 412954
rect -9036 412634 592960 412718
rect -9036 412398 -5164 412634
rect -4928 412398 -4844 412634
rect -4608 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588532 412634
rect 588768 412398 588852 412634
rect 589088 412398 592960 412634
rect -9036 412366 592960 412398
rect -9036 408454 592960 408486
rect -9036 408218 -4204 408454
rect -3968 408218 -3884 408454
rect -3648 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587572 408454
rect 587808 408218 587892 408454
rect 588128 408218 592960 408454
rect -9036 408134 592960 408218
rect -9036 407898 -4204 408134
rect -3968 407898 -3884 408134
rect -3648 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587572 408134
rect 587808 407898 587892 408134
rect 588128 407898 592960 408134
rect -9036 407866 592960 407898
rect -9036 403954 592960 403986
rect -9036 403718 -3244 403954
rect -3008 403718 -2924 403954
rect -2688 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 252010 403954
rect 252246 403718 282730 403954
rect 282966 403718 313450 403954
rect 313686 403718 344170 403954
rect 344406 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586612 403954
rect 586848 403718 586932 403954
rect 587168 403718 592960 403954
rect -9036 403634 592960 403718
rect -9036 403398 -3244 403634
rect -3008 403398 -2924 403634
rect -2688 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 252010 403634
rect 252246 403398 282730 403634
rect 282966 403398 313450 403634
rect 313686 403398 344170 403634
rect 344406 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586612 403634
rect 586848 403398 586932 403634
rect 587168 403398 592960 403634
rect -9036 403366 592960 403398
rect -9036 399454 592960 399486
rect -9036 399218 -2284 399454
rect -2048 399218 -1964 399454
rect -1728 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 236650 399454
rect 236886 399218 267370 399454
rect 267606 399218 298090 399454
rect 298326 399218 328810 399454
rect 329046 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585652 399454
rect 585888 399218 585972 399454
rect 586208 399218 592960 399454
rect -9036 399134 592960 399218
rect -9036 398898 -2284 399134
rect -2048 398898 -1964 399134
rect -1728 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 236650 399134
rect 236886 398898 267370 399134
rect 267606 398898 298090 399134
rect 298326 398898 328810 399134
rect 329046 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585652 399134
rect 585888 398898 585972 399134
rect 586208 398898 592960 399134
rect -9036 398866 592960 398898
rect -9036 394954 592960 394986
rect -9036 394718 -9004 394954
rect -8768 394718 -8684 394954
rect -8448 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592372 394954
rect 592608 394718 592692 394954
rect 592928 394718 592960 394954
rect -9036 394634 592960 394718
rect -9036 394398 -9004 394634
rect -8768 394398 -8684 394634
rect -8448 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592372 394634
rect 592608 394398 592692 394634
rect 592928 394398 592960 394634
rect -9036 394366 592960 394398
rect -9036 390454 592960 390486
rect -9036 390218 -8044 390454
rect -7808 390218 -7724 390454
rect -7488 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591412 390454
rect 591648 390218 591732 390454
rect 591968 390218 592960 390454
rect -9036 390134 592960 390218
rect -9036 389898 -8044 390134
rect -7808 389898 -7724 390134
rect -7488 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591412 390134
rect 591648 389898 591732 390134
rect 591968 389898 592960 390134
rect -9036 389866 592960 389898
rect -9036 385954 592960 385986
rect -9036 385718 -7084 385954
rect -6848 385718 -6764 385954
rect -6528 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590452 385954
rect 590688 385718 590772 385954
rect 591008 385718 592960 385954
rect -9036 385634 592960 385718
rect -9036 385398 -7084 385634
rect -6848 385398 -6764 385634
rect -6528 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590452 385634
rect 590688 385398 590772 385634
rect 591008 385398 592960 385634
rect -9036 385366 592960 385398
rect -9036 381454 592960 381486
rect -9036 381218 -6124 381454
rect -5888 381218 -5804 381454
rect -5568 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589492 381454
rect 589728 381218 589812 381454
rect 590048 381218 592960 381454
rect -9036 381134 592960 381218
rect -9036 380898 -6124 381134
rect -5888 380898 -5804 381134
rect -5568 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589492 381134
rect 589728 380898 589812 381134
rect 590048 380898 592960 381134
rect -9036 380866 592960 380898
rect -9036 376954 592960 376986
rect -9036 376718 -5164 376954
rect -4928 376718 -4844 376954
rect -4608 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588532 376954
rect 588768 376718 588852 376954
rect 589088 376718 592960 376954
rect -9036 376634 592960 376718
rect -9036 376398 -5164 376634
rect -4928 376398 -4844 376634
rect -4608 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588532 376634
rect 588768 376398 588852 376634
rect 589088 376398 592960 376634
rect -9036 376366 592960 376398
rect -9036 372454 592960 372486
rect -9036 372218 -4204 372454
rect -3968 372218 -3884 372454
rect -3648 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587572 372454
rect 587808 372218 587892 372454
rect 588128 372218 592960 372454
rect -9036 372134 592960 372218
rect -9036 371898 -4204 372134
rect -3968 371898 -3884 372134
rect -3648 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587572 372134
rect 587808 371898 587892 372134
rect 588128 371898 592960 372134
rect -9036 371866 592960 371898
rect -9036 367954 592960 367986
rect -9036 367718 -3244 367954
rect -3008 367718 -2924 367954
rect -2688 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 119610 367954
rect 119846 367718 150330 367954
rect 150566 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 252010 367954
rect 252246 367718 282730 367954
rect 282966 367718 313450 367954
rect 313686 367718 344170 367954
rect 344406 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586612 367954
rect 586848 367718 586932 367954
rect 587168 367718 592960 367954
rect -9036 367634 592960 367718
rect -9036 367398 -3244 367634
rect -3008 367398 -2924 367634
rect -2688 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 119610 367634
rect 119846 367398 150330 367634
rect 150566 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 252010 367634
rect 252246 367398 282730 367634
rect 282966 367398 313450 367634
rect 313686 367398 344170 367634
rect 344406 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586612 367634
rect 586848 367398 586932 367634
rect 587168 367398 592960 367634
rect -9036 367366 592960 367398
rect -9036 363454 592960 363486
rect -9036 363218 -2284 363454
rect -2048 363218 -1964 363454
rect -1728 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 104250 363454
rect 104486 363218 134970 363454
rect 135206 363218 165690 363454
rect 165926 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 236650 363454
rect 236886 363218 267370 363454
rect 267606 363218 298090 363454
rect 298326 363218 328810 363454
rect 329046 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585652 363454
rect 585888 363218 585972 363454
rect 586208 363218 592960 363454
rect -9036 363134 592960 363218
rect -9036 362898 -2284 363134
rect -2048 362898 -1964 363134
rect -1728 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 104250 363134
rect 104486 362898 134970 363134
rect 135206 362898 165690 363134
rect 165926 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 236650 363134
rect 236886 362898 267370 363134
rect 267606 362898 298090 363134
rect 298326 362898 328810 363134
rect 329046 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585652 363134
rect 585888 362898 585972 363134
rect 586208 362898 592960 363134
rect -9036 362866 592960 362898
rect -9036 358954 592960 358986
rect -9036 358718 -9004 358954
rect -8768 358718 -8684 358954
rect -8448 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592372 358954
rect 592608 358718 592692 358954
rect 592928 358718 592960 358954
rect -9036 358634 592960 358718
rect -9036 358398 -9004 358634
rect -8768 358398 -8684 358634
rect -8448 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592372 358634
rect 592608 358398 592692 358634
rect 592928 358398 592960 358634
rect -9036 358366 592960 358398
rect -9036 354454 592960 354486
rect -9036 354218 -8044 354454
rect -7808 354218 -7724 354454
rect -7488 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591412 354454
rect 591648 354218 591732 354454
rect 591968 354218 592960 354454
rect -9036 354134 592960 354218
rect -9036 353898 -8044 354134
rect -7808 353898 -7724 354134
rect -7488 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591412 354134
rect 591648 353898 591732 354134
rect 591968 353898 592960 354134
rect -9036 353866 592960 353898
rect -9036 349954 592960 349986
rect -9036 349718 -7084 349954
rect -6848 349718 -6764 349954
rect -6528 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590452 349954
rect 590688 349718 590772 349954
rect 591008 349718 592960 349954
rect -9036 349634 592960 349718
rect -9036 349398 -7084 349634
rect -6848 349398 -6764 349634
rect -6528 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590452 349634
rect 590688 349398 590772 349634
rect 591008 349398 592960 349634
rect -9036 349366 592960 349398
rect -9036 345454 592960 345486
rect -9036 345218 -6124 345454
rect -5888 345218 -5804 345454
rect -5568 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589492 345454
rect 589728 345218 589812 345454
rect 590048 345218 592960 345454
rect -9036 345134 592960 345218
rect -9036 344898 -6124 345134
rect -5888 344898 -5804 345134
rect -5568 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589492 345134
rect 589728 344898 589812 345134
rect 590048 344898 592960 345134
rect -9036 344866 592960 344898
rect -9036 340954 592960 340986
rect -9036 340718 -5164 340954
rect -4928 340718 -4844 340954
rect -4608 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588532 340954
rect 588768 340718 588852 340954
rect 589088 340718 592960 340954
rect -9036 340634 592960 340718
rect -9036 340398 -5164 340634
rect -4928 340398 -4844 340634
rect -4608 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588532 340634
rect 588768 340398 588852 340634
rect 589088 340398 592960 340634
rect -9036 340366 592960 340398
rect -9036 336454 592960 336486
rect -9036 336218 -4204 336454
rect -3968 336218 -3884 336454
rect -3648 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587572 336454
rect 587808 336218 587892 336454
rect 588128 336218 592960 336454
rect -9036 336134 592960 336218
rect -9036 335898 -4204 336134
rect -3968 335898 -3884 336134
rect -3648 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587572 336134
rect 587808 335898 587892 336134
rect 588128 335898 592960 336134
rect -9036 335866 592960 335898
rect -9036 331954 592960 331986
rect -9036 331718 -3244 331954
rect -3008 331718 -2924 331954
rect -2688 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 119610 331954
rect 119846 331718 150330 331954
rect 150566 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 252010 331954
rect 252246 331718 282730 331954
rect 282966 331718 313450 331954
rect 313686 331718 344170 331954
rect 344406 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586612 331954
rect 586848 331718 586932 331954
rect 587168 331718 592960 331954
rect -9036 331634 592960 331718
rect -9036 331398 -3244 331634
rect -3008 331398 -2924 331634
rect -2688 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 119610 331634
rect 119846 331398 150330 331634
rect 150566 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 252010 331634
rect 252246 331398 282730 331634
rect 282966 331398 313450 331634
rect 313686 331398 344170 331634
rect 344406 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586612 331634
rect 586848 331398 586932 331634
rect 587168 331398 592960 331634
rect -9036 331366 592960 331398
rect -9036 327454 592960 327486
rect -9036 327218 -2284 327454
rect -2048 327218 -1964 327454
rect -1728 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 104250 327454
rect 104486 327218 134970 327454
rect 135206 327218 165690 327454
rect 165926 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 236650 327454
rect 236886 327218 267370 327454
rect 267606 327218 298090 327454
rect 298326 327218 328810 327454
rect 329046 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585652 327454
rect 585888 327218 585972 327454
rect 586208 327218 592960 327454
rect -9036 327134 592960 327218
rect -9036 326898 -2284 327134
rect -2048 326898 -1964 327134
rect -1728 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 104250 327134
rect 104486 326898 134970 327134
rect 135206 326898 165690 327134
rect 165926 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 236650 327134
rect 236886 326898 267370 327134
rect 267606 326898 298090 327134
rect 298326 326898 328810 327134
rect 329046 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585652 327134
rect 585888 326898 585972 327134
rect 586208 326898 592960 327134
rect -9036 326866 592960 326898
rect -9036 322954 592960 322986
rect -9036 322718 -9004 322954
rect -8768 322718 -8684 322954
rect -8448 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592372 322954
rect 592608 322718 592692 322954
rect 592928 322718 592960 322954
rect -9036 322634 592960 322718
rect -9036 322398 -9004 322634
rect -8768 322398 -8684 322634
rect -8448 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592372 322634
rect 592608 322398 592692 322634
rect 592928 322398 592960 322634
rect -9036 322366 592960 322398
rect -9036 318454 592960 318486
rect -9036 318218 -8044 318454
rect -7808 318218 -7724 318454
rect -7488 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591412 318454
rect 591648 318218 591732 318454
rect 591968 318218 592960 318454
rect -9036 318134 592960 318218
rect -9036 317898 -8044 318134
rect -7808 317898 -7724 318134
rect -7488 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591412 318134
rect 591648 317898 591732 318134
rect 591968 317898 592960 318134
rect -9036 317866 592960 317898
rect -9036 313954 592960 313986
rect -9036 313718 -7084 313954
rect -6848 313718 -6764 313954
rect -6528 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590452 313954
rect 590688 313718 590772 313954
rect 591008 313718 592960 313954
rect -9036 313634 592960 313718
rect -9036 313398 -7084 313634
rect -6848 313398 -6764 313634
rect -6528 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590452 313634
rect 590688 313398 590772 313634
rect 591008 313398 592960 313634
rect -9036 313366 592960 313398
rect -9036 309454 592960 309486
rect -9036 309218 -6124 309454
rect -5888 309218 -5804 309454
rect -5568 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589492 309454
rect 589728 309218 589812 309454
rect 590048 309218 592960 309454
rect -9036 309134 592960 309218
rect -9036 308898 -6124 309134
rect -5888 308898 -5804 309134
rect -5568 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589492 309134
rect 589728 308898 589812 309134
rect 590048 308898 592960 309134
rect -9036 308866 592960 308898
rect -9036 304954 592960 304986
rect -9036 304718 -5164 304954
rect -4928 304718 -4844 304954
rect -4608 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588532 304954
rect 588768 304718 588852 304954
rect 589088 304718 592960 304954
rect -9036 304634 592960 304718
rect -9036 304398 -5164 304634
rect -4928 304398 -4844 304634
rect -4608 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588532 304634
rect 588768 304398 588852 304634
rect 589088 304398 592960 304634
rect -9036 304366 592960 304398
rect -9036 300454 592960 300486
rect -9036 300218 -4204 300454
rect -3968 300218 -3884 300454
rect -3648 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587572 300454
rect 587808 300218 587892 300454
rect 588128 300218 592960 300454
rect -9036 300134 592960 300218
rect -9036 299898 -4204 300134
rect -3968 299898 -3884 300134
rect -3648 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587572 300134
rect 587808 299898 587892 300134
rect 588128 299898 592960 300134
rect -9036 299866 592960 299898
rect -9036 295954 592960 295986
rect -9036 295718 -3244 295954
rect -3008 295718 -2924 295954
rect -2688 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586612 295954
rect 586848 295718 586932 295954
rect 587168 295718 592960 295954
rect -9036 295634 592960 295718
rect -9036 295398 -3244 295634
rect -3008 295398 -2924 295634
rect -2688 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586612 295634
rect 586848 295398 586932 295634
rect 587168 295398 592960 295634
rect -9036 295366 592960 295398
rect -9036 291454 592960 291486
rect -9036 291218 -2284 291454
rect -2048 291218 -1964 291454
rect -1728 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585652 291454
rect 585888 291218 585972 291454
rect 586208 291218 592960 291454
rect -9036 291134 592960 291218
rect -9036 290898 -2284 291134
rect -2048 290898 -1964 291134
rect -1728 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585652 291134
rect 585888 290898 585972 291134
rect 586208 290898 592960 291134
rect -9036 290866 592960 290898
rect -9036 286954 592960 286986
rect -9036 286718 -9004 286954
rect -8768 286718 -8684 286954
rect -8448 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592372 286954
rect 592608 286718 592692 286954
rect 592928 286718 592960 286954
rect -9036 286634 592960 286718
rect -9036 286398 -9004 286634
rect -8768 286398 -8684 286634
rect -8448 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592372 286634
rect 592608 286398 592692 286634
rect 592928 286398 592960 286634
rect -9036 286366 592960 286398
rect -9036 282454 592960 282486
rect -9036 282218 -8044 282454
rect -7808 282218 -7724 282454
rect -7488 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591412 282454
rect 591648 282218 591732 282454
rect 591968 282218 592960 282454
rect -9036 282134 592960 282218
rect -9036 281898 -8044 282134
rect -7808 281898 -7724 282134
rect -7488 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591412 282134
rect 591648 281898 591732 282134
rect 591968 281898 592960 282134
rect -9036 281866 592960 281898
rect -9036 277954 592960 277986
rect -9036 277718 -7084 277954
rect -6848 277718 -6764 277954
rect -6528 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590452 277954
rect 590688 277718 590772 277954
rect 591008 277718 592960 277954
rect -9036 277634 592960 277718
rect -9036 277398 -7084 277634
rect -6848 277398 -6764 277634
rect -6528 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590452 277634
rect 590688 277398 590772 277634
rect 591008 277398 592960 277634
rect -9036 277366 592960 277398
rect -9036 273454 592960 273486
rect -9036 273218 -6124 273454
rect -5888 273218 -5804 273454
rect -5568 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589492 273454
rect 589728 273218 589812 273454
rect 590048 273218 592960 273454
rect -9036 273134 592960 273218
rect -9036 272898 -6124 273134
rect -5888 272898 -5804 273134
rect -5568 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589492 273134
rect 589728 272898 589812 273134
rect 590048 272898 592960 273134
rect -9036 272866 592960 272898
rect -9036 268954 592960 268986
rect -9036 268718 -5164 268954
rect -4928 268718 -4844 268954
rect -4608 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588532 268954
rect 588768 268718 588852 268954
rect 589088 268718 592960 268954
rect -9036 268634 592960 268718
rect -9036 268398 -5164 268634
rect -4928 268398 -4844 268634
rect -4608 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588532 268634
rect 588768 268398 588852 268634
rect 589088 268398 592960 268634
rect -9036 268366 592960 268398
rect -9036 264454 592960 264486
rect -9036 264218 -4204 264454
rect -3968 264218 -3884 264454
rect -3648 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587572 264454
rect 587808 264218 587892 264454
rect 588128 264218 592960 264454
rect -9036 264134 592960 264218
rect -9036 263898 -4204 264134
rect -3968 263898 -3884 264134
rect -3648 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587572 264134
rect 587808 263898 587892 264134
rect 588128 263898 592960 264134
rect -9036 263866 592960 263898
rect -9036 259954 592960 259986
rect -9036 259718 -3244 259954
rect -3008 259718 -2924 259954
rect -2688 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586612 259954
rect 586848 259718 586932 259954
rect 587168 259718 592960 259954
rect -9036 259634 592960 259718
rect -9036 259398 -3244 259634
rect -3008 259398 -2924 259634
rect -2688 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586612 259634
rect 586848 259398 586932 259634
rect 587168 259398 592960 259634
rect -9036 259366 592960 259398
rect -9036 255454 592960 255486
rect -9036 255218 -2284 255454
rect -2048 255218 -1964 255454
rect -1728 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585652 255454
rect 585888 255218 585972 255454
rect 586208 255218 592960 255454
rect -9036 255134 592960 255218
rect -9036 254898 -2284 255134
rect -2048 254898 -1964 255134
rect -1728 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585652 255134
rect 585888 254898 585972 255134
rect 586208 254898 592960 255134
rect -9036 254866 592960 254898
rect -9036 250954 592960 250986
rect -9036 250718 -9004 250954
rect -8768 250718 -8684 250954
rect -8448 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592372 250954
rect 592608 250718 592692 250954
rect 592928 250718 592960 250954
rect -9036 250634 592960 250718
rect -9036 250398 -9004 250634
rect -8768 250398 -8684 250634
rect -8448 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592372 250634
rect 592608 250398 592692 250634
rect 592928 250398 592960 250634
rect -9036 250366 592960 250398
rect -9036 246454 592960 246486
rect -9036 246218 -8044 246454
rect -7808 246218 -7724 246454
rect -7488 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591412 246454
rect 591648 246218 591732 246454
rect 591968 246218 592960 246454
rect -9036 246134 592960 246218
rect -9036 245898 -8044 246134
rect -7808 245898 -7724 246134
rect -7488 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591412 246134
rect 591648 245898 591732 246134
rect 591968 245898 592960 246134
rect -9036 245866 592960 245898
rect -9036 241954 592960 241986
rect -9036 241718 -7084 241954
rect -6848 241718 -6764 241954
rect -6528 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590452 241954
rect 590688 241718 590772 241954
rect 591008 241718 592960 241954
rect -9036 241634 592960 241718
rect -9036 241398 -7084 241634
rect -6848 241398 -6764 241634
rect -6528 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590452 241634
rect 590688 241398 590772 241634
rect 591008 241398 592960 241634
rect -9036 241366 592960 241398
rect -9036 237454 592960 237486
rect -9036 237218 -6124 237454
rect -5888 237218 -5804 237454
rect -5568 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589492 237454
rect 589728 237218 589812 237454
rect 590048 237218 592960 237454
rect -9036 237134 592960 237218
rect -9036 236898 -6124 237134
rect -5888 236898 -5804 237134
rect -5568 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589492 237134
rect 589728 236898 589812 237134
rect 590048 236898 592960 237134
rect -9036 236866 592960 236898
rect -9036 232954 592960 232986
rect -9036 232718 -5164 232954
rect -4928 232718 -4844 232954
rect -4608 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588532 232954
rect 588768 232718 588852 232954
rect 589088 232718 592960 232954
rect -9036 232634 592960 232718
rect -9036 232398 -5164 232634
rect -4928 232398 -4844 232634
rect -4608 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588532 232634
rect 588768 232398 588852 232634
rect 589088 232398 592960 232634
rect -9036 232366 592960 232398
rect -9036 228454 592960 228486
rect -9036 228218 -4204 228454
rect -3968 228218 -3884 228454
rect -3648 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587572 228454
rect 587808 228218 587892 228454
rect 588128 228218 592960 228454
rect -9036 228134 592960 228218
rect -9036 227898 -4204 228134
rect -3968 227898 -3884 228134
rect -3648 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587572 228134
rect 587808 227898 587892 228134
rect 588128 227898 592960 228134
rect -9036 227866 592960 227898
rect -9036 223954 592960 223986
rect -9036 223718 -3244 223954
rect -3008 223718 -2924 223954
rect -2688 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 220328 223954
rect 220564 223718 356056 223954
rect 356292 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586612 223954
rect 586848 223718 586932 223954
rect 587168 223718 592960 223954
rect -9036 223634 592960 223718
rect -9036 223398 -3244 223634
rect -3008 223398 -2924 223634
rect -2688 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 220328 223634
rect 220564 223398 356056 223634
rect 356292 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586612 223634
rect 586848 223398 586932 223634
rect 587168 223398 592960 223634
rect -9036 223366 592960 223398
rect -9036 219454 592960 219486
rect -9036 219218 -2284 219454
rect -2048 219218 -1964 219454
rect -1728 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 221008 219454
rect 221244 219218 355376 219454
rect 355612 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585652 219454
rect 585888 219218 585972 219454
rect 586208 219218 592960 219454
rect -9036 219134 592960 219218
rect -9036 218898 -2284 219134
rect -2048 218898 -1964 219134
rect -1728 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 221008 219134
rect 221244 218898 355376 219134
rect 355612 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585652 219134
rect 585888 218898 585972 219134
rect 586208 218898 592960 219134
rect -9036 218866 592960 218898
rect -9036 214954 592960 214986
rect -9036 214718 -9004 214954
rect -8768 214718 -8684 214954
rect -8448 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592372 214954
rect 592608 214718 592692 214954
rect 592928 214718 592960 214954
rect -9036 214634 592960 214718
rect -9036 214398 -9004 214634
rect -8768 214398 -8684 214634
rect -8448 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592372 214634
rect 592608 214398 592692 214634
rect 592928 214398 592960 214634
rect -9036 214366 592960 214398
rect -9036 210454 592960 210486
rect -9036 210218 -8044 210454
rect -7808 210218 -7724 210454
rect -7488 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591412 210454
rect 591648 210218 591732 210454
rect 591968 210218 592960 210454
rect -9036 210134 592960 210218
rect -9036 209898 -8044 210134
rect -7808 209898 -7724 210134
rect -7488 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591412 210134
rect 591648 209898 591732 210134
rect 591968 209898 592960 210134
rect -9036 209866 592960 209898
rect -9036 205954 592960 205986
rect -9036 205718 -7084 205954
rect -6848 205718 -6764 205954
rect -6528 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590452 205954
rect 590688 205718 590772 205954
rect 591008 205718 592960 205954
rect -9036 205634 592960 205718
rect -9036 205398 -7084 205634
rect -6848 205398 -6764 205634
rect -6528 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590452 205634
rect 590688 205398 590772 205634
rect 591008 205398 592960 205634
rect -9036 205366 592960 205398
rect -9036 201454 592960 201486
rect -9036 201218 -6124 201454
rect -5888 201218 -5804 201454
rect -5568 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589492 201454
rect 589728 201218 589812 201454
rect 590048 201218 592960 201454
rect -9036 201134 592960 201218
rect -9036 200898 -6124 201134
rect -5888 200898 -5804 201134
rect -5568 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589492 201134
rect 589728 200898 589812 201134
rect 590048 200898 592960 201134
rect -9036 200866 592960 200898
rect -9036 196954 592960 196986
rect -9036 196718 -5164 196954
rect -4928 196718 -4844 196954
rect -4608 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588532 196954
rect 588768 196718 588852 196954
rect 589088 196718 592960 196954
rect -9036 196634 592960 196718
rect -9036 196398 -5164 196634
rect -4928 196398 -4844 196634
rect -4608 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588532 196634
rect 588768 196398 588852 196634
rect 589088 196398 592960 196634
rect -9036 196366 592960 196398
rect -9036 192454 592960 192486
rect -9036 192218 -4204 192454
rect -3968 192218 -3884 192454
rect -3648 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587572 192454
rect 587808 192218 587892 192454
rect 588128 192218 592960 192454
rect -9036 192134 592960 192218
rect -9036 191898 -4204 192134
rect -3968 191898 -3884 192134
rect -3648 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587572 192134
rect 587808 191898 587892 192134
rect 588128 191898 592960 192134
rect -9036 191866 592960 191898
rect -9036 187954 592960 187986
rect -9036 187718 -3244 187954
rect -3008 187718 -2924 187954
rect -2688 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 220328 187954
rect 220564 187718 356056 187954
rect 356292 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586612 187954
rect 586848 187718 586932 187954
rect 587168 187718 592960 187954
rect -9036 187634 592960 187718
rect -9036 187398 -3244 187634
rect -3008 187398 -2924 187634
rect -2688 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 220328 187634
rect 220564 187398 356056 187634
rect 356292 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586612 187634
rect 586848 187398 586932 187634
rect 587168 187398 592960 187634
rect -9036 187366 592960 187398
rect -9036 183454 592960 183486
rect -9036 183218 -2284 183454
rect -2048 183218 -1964 183454
rect -1728 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 221008 183454
rect 221244 183218 355376 183454
rect 355612 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585652 183454
rect 585888 183218 585972 183454
rect 586208 183218 592960 183454
rect -9036 183134 592960 183218
rect -9036 182898 -2284 183134
rect -2048 182898 -1964 183134
rect -1728 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 221008 183134
rect 221244 182898 355376 183134
rect 355612 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585652 183134
rect 585888 182898 585972 183134
rect 586208 182898 592960 183134
rect -9036 182866 592960 182898
rect -9036 178954 592960 178986
rect -9036 178718 -9004 178954
rect -8768 178718 -8684 178954
rect -8448 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592372 178954
rect 592608 178718 592692 178954
rect 592928 178718 592960 178954
rect -9036 178634 592960 178718
rect -9036 178398 -9004 178634
rect -8768 178398 -8684 178634
rect -8448 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592372 178634
rect 592608 178398 592692 178634
rect 592928 178398 592960 178634
rect -9036 178366 592960 178398
rect -9036 174454 592960 174486
rect -9036 174218 -8044 174454
rect -7808 174218 -7724 174454
rect -7488 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591412 174454
rect 591648 174218 591732 174454
rect 591968 174218 592960 174454
rect -9036 174134 592960 174218
rect -9036 173898 -8044 174134
rect -7808 173898 -7724 174134
rect -7488 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591412 174134
rect 591648 173898 591732 174134
rect 591968 173898 592960 174134
rect -9036 173866 592960 173898
rect -9036 169954 592960 169986
rect -9036 169718 -7084 169954
rect -6848 169718 -6764 169954
rect -6528 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590452 169954
rect 590688 169718 590772 169954
rect 591008 169718 592960 169954
rect -9036 169634 592960 169718
rect -9036 169398 -7084 169634
rect -6848 169398 -6764 169634
rect -6528 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590452 169634
rect 590688 169398 590772 169634
rect 591008 169398 592960 169634
rect -9036 169366 592960 169398
rect -9036 165454 592960 165486
rect -9036 165218 -6124 165454
rect -5888 165218 -5804 165454
rect -5568 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589492 165454
rect 589728 165218 589812 165454
rect 590048 165218 592960 165454
rect -9036 165134 592960 165218
rect -9036 164898 -6124 165134
rect -5888 164898 -5804 165134
rect -5568 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589492 165134
rect 589728 164898 589812 165134
rect 590048 164898 592960 165134
rect -9036 164866 592960 164898
rect -9036 160954 592960 160986
rect -9036 160718 -5164 160954
rect -4928 160718 -4844 160954
rect -4608 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588532 160954
rect 588768 160718 588852 160954
rect 589088 160718 592960 160954
rect -9036 160634 592960 160718
rect -9036 160398 -5164 160634
rect -4928 160398 -4844 160634
rect -4608 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588532 160634
rect 588768 160398 588852 160634
rect 589088 160398 592960 160634
rect -9036 160366 592960 160398
rect -9036 156454 592960 156486
rect -9036 156218 -4204 156454
rect -3968 156218 -3884 156454
rect -3648 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587572 156454
rect 587808 156218 587892 156454
rect 588128 156218 592960 156454
rect -9036 156134 592960 156218
rect -9036 155898 -4204 156134
rect -3968 155898 -3884 156134
rect -3648 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587572 156134
rect 587808 155898 587892 156134
rect 588128 155898 592960 156134
rect -9036 155866 592960 155898
rect -9036 151954 592960 151986
rect -9036 151718 -3244 151954
rect -3008 151718 -2924 151954
rect -2688 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586612 151954
rect 586848 151718 586932 151954
rect 587168 151718 592960 151954
rect -9036 151634 592960 151718
rect -9036 151398 -3244 151634
rect -3008 151398 -2924 151634
rect -2688 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586612 151634
rect 586848 151398 586932 151634
rect 587168 151398 592960 151634
rect -9036 151366 592960 151398
rect -9036 147454 592960 147486
rect -9036 147218 -2284 147454
rect -2048 147218 -1964 147454
rect -1728 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585652 147454
rect 585888 147218 585972 147454
rect 586208 147218 592960 147454
rect -9036 147134 592960 147218
rect -9036 146898 -2284 147134
rect -2048 146898 -1964 147134
rect -1728 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585652 147134
rect 585888 146898 585972 147134
rect 586208 146898 592960 147134
rect -9036 146866 592960 146898
rect -9036 142954 592960 142986
rect -9036 142718 -9004 142954
rect -8768 142718 -8684 142954
rect -8448 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592372 142954
rect 592608 142718 592692 142954
rect 592928 142718 592960 142954
rect -9036 142634 592960 142718
rect -9036 142398 -9004 142634
rect -8768 142398 -8684 142634
rect -8448 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592372 142634
rect 592608 142398 592692 142634
rect 592928 142398 592960 142634
rect -9036 142366 592960 142398
rect -9036 138454 592960 138486
rect -9036 138218 -8044 138454
rect -7808 138218 -7724 138454
rect -7488 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591412 138454
rect 591648 138218 591732 138454
rect 591968 138218 592960 138454
rect -9036 138134 592960 138218
rect -9036 137898 -8044 138134
rect -7808 137898 -7724 138134
rect -7488 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591412 138134
rect 591648 137898 591732 138134
rect 591968 137898 592960 138134
rect -9036 137866 592960 137898
rect -9036 133954 592960 133986
rect -9036 133718 -7084 133954
rect -6848 133718 -6764 133954
rect -6528 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590452 133954
rect 590688 133718 590772 133954
rect 591008 133718 592960 133954
rect -9036 133634 592960 133718
rect -9036 133398 -7084 133634
rect -6848 133398 -6764 133634
rect -6528 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590452 133634
rect 590688 133398 590772 133634
rect 591008 133398 592960 133634
rect -9036 133366 592960 133398
rect -9036 129454 592960 129486
rect -9036 129218 -6124 129454
rect -5888 129218 -5804 129454
rect -5568 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589492 129454
rect 589728 129218 589812 129454
rect 590048 129218 592960 129454
rect -9036 129134 592960 129218
rect -9036 128898 -6124 129134
rect -5888 128898 -5804 129134
rect -5568 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589492 129134
rect 589728 128898 589812 129134
rect 590048 128898 592960 129134
rect -9036 128866 592960 128898
rect -9036 124954 592960 124986
rect -9036 124718 -5164 124954
rect -4928 124718 -4844 124954
rect -4608 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 123326 124954
rect 123562 124718 123646 124954
rect 123882 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588532 124954
rect 588768 124718 588852 124954
rect 589088 124718 592960 124954
rect -9036 124634 592960 124718
rect -9036 124398 -5164 124634
rect -4928 124398 -4844 124634
rect -4608 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 123326 124634
rect 123562 124398 123646 124634
rect 123882 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588532 124634
rect 588768 124398 588852 124634
rect 589088 124398 592960 124634
rect -9036 124366 592960 124398
rect -9036 120454 592960 120486
rect -9036 120218 -4204 120454
rect -3968 120218 -3884 120454
rect -3648 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587572 120454
rect 587808 120218 587892 120454
rect 588128 120218 592960 120454
rect -9036 120134 592960 120218
rect -9036 119898 -4204 120134
rect -3968 119898 -3884 120134
rect -3648 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587572 120134
rect 587808 119898 587892 120134
rect 588128 119898 592960 120134
rect -9036 119866 592960 119898
rect -9036 115954 592960 115986
rect -9036 115718 -3244 115954
rect -3008 115718 -2924 115954
rect -2688 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586612 115954
rect 586848 115718 586932 115954
rect 587168 115718 592960 115954
rect -9036 115634 592960 115718
rect -9036 115398 -3244 115634
rect -3008 115398 -2924 115634
rect -2688 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586612 115634
rect 586848 115398 586932 115634
rect 587168 115398 592960 115634
rect -9036 115366 592960 115398
rect -9036 111454 592960 111486
rect -9036 111218 -2284 111454
rect -2048 111218 -1964 111454
rect -1728 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585652 111454
rect 585888 111218 585972 111454
rect 586208 111218 592960 111454
rect -9036 111134 592960 111218
rect -9036 110898 -2284 111134
rect -2048 110898 -1964 111134
rect -1728 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585652 111134
rect 585888 110898 585972 111134
rect 586208 110898 592960 111134
rect -9036 110866 592960 110898
rect -9036 106954 592960 106986
rect -9036 106718 -9004 106954
rect -8768 106718 -8684 106954
rect -8448 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592372 106954
rect 592608 106718 592692 106954
rect 592928 106718 592960 106954
rect -9036 106634 592960 106718
rect -9036 106398 -9004 106634
rect -8768 106398 -8684 106634
rect -8448 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592372 106634
rect 592608 106398 592692 106634
rect 592928 106398 592960 106634
rect -9036 106366 592960 106398
rect -9036 102454 592960 102486
rect -9036 102218 -8044 102454
rect -7808 102218 -7724 102454
rect -7488 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591412 102454
rect 591648 102218 591732 102454
rect 591968 102218 592960 102454
rect -9036 102134 592960 102218
rect -9036 101898 -8044 102134
rect -7808 101898 -7724 102134
rect -7488 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591412 102134
rect 591648 101898 591732 102134
rect 591968 101898 592960 102134
rect -9036 101866 592960 101898
rect -9036 97954 592960 97986
rect -9036 97718 -7084 97954
rect -6848 97718 -6764 97954
rect -6528 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590452 97954
rect 590688 97718 590772 97954
rect 591008 97718 592960 97954
rect -9036 97634 592960 97718
rect -9036 97398 -7084 97634
rect -6848 97398 -6764 97634
rect -6528 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590452 97634
rect 590688 97398 590772 97634
rect 591008 97398 592960 97634
rect -9036 97366 592960 97398
rect -9036 93454 592960 93486
rect -9036 93218 -6124 93454
rect -5888 93218 -5804 93454
rect -5568 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589492 93454
rect 589728 93218 589812 93454
rect 590048 93218 592960 93454
rect -9036 93134 592960 93218
rect -9036 92898 -6124 93134
rect -5888 92898 -5804 93134
rect -5568 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589492 93134
rect 589728 92898 589812 93134
rect 590048 92898 592960 93134
rect -9036 92866 592960 92898
rect -9036 88954 592960 88986
rect -9036 88718 -5164 88954
rect -4928 88718 -4844 88954
rect -4608 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588532 88954
rect 588768 88718 588852 88954
rect 589088 88718 592960 88954
rect -9036 88634 592960 88718
rect -9036 88398 -5164 88634
rect -4928 88398 -4844 88634
rect -4608 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588532 88634
rect 588768 88398 588852 88634
rect 589088 88398 592960 88634
rect -9036 88366 592960 88398
rect -9036 84454 592960 84486
rect -9036 84218 -4204 84454
rect -3968 84218 -3884 84454
rect -3648 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587572 84454
rect 587808 84218 587892 84454
rect 588128 84218 592960 84454
rect -9036 84134 592960 84218
rect -9036 83898 -4204 84134
rect -3968 83898 -3884 84134
rect -3648 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587572 84134
rect 587808 83898 587892 84134
rect 588128 83898 592960 84134
rect -9036 83866 592960 83898
rect -9036 79954 592960 79986
rect -9036 79718 -3244 79954
rect -3008 79718 -2924 79954
rect -2688 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586612 79954
rect 586848 79718 586932 79954
rect 587168 79718 592960 79954
rect -9036 79634 592960 79718
rect -9036 79398 -3244 79634
rect -3008 79398 -2924 79634
rect -2688 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586612 79634
rect 586848 79398 586932 79634
rect 587168 79398 592960 79634
rect -9036 79366 592960 79398
rect -9036 75454 592960 75486
rect -9036 75218 -2284 75454
rect -2048 75218 -1964 75454
rect -1728 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585652 75454
rect 585888 75218 585972 75454
rect 586208 75218 592960 75454
rect -9036 75134 592960 75218
rect -9036 74898 -2284 75134
rect -2048 74898 -1964 75134
rect -1728 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585652 75134
rect 585888 74898 585972 75134
rect 586208 74898 592960 75134
rect -9036 74866 592960 74898
rect -9036 70954 592960 70986
rect -9036 70718 -9004 70954
rect -8768 70718 -8684 70954
rect -8448 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592372 70954
rect 592608 70718 592692 70954
rect 592928 70718 592960 70954
rect -9036 70634 592960 70718
rect -9036 70398 -9004 70634
rect -8768 70398 -8684 70634
rect -8448 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592372 70634
rect 592608 70398 592692 70634
rect 592928 70398 592960 70634
rect -9036 70366 592960 70398
rect -9036 66454 592960 66486
rect -9036 66218 -8044 66454
rect -7808 66218 -7724 66454
rect -7488 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591412 66454
rect 591648 66218 591732 66454
rect 591968 66218 592960 66454
rect -9036 66134 592960 66218
rect -9036 65898 -8044 66134
rect -7808 65898 -7724 66134
rect -7488 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591412 66134
rect 591648 65898 591732 66134
rect 591968 65898 592960 66134
rect -9036 65866 592960 65898
rect -9036 61954 592960 61986
rect -9036 61718 -7084 61954
rect -6848 61718 -6764 61954
rect -6528 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590452 61954
rect 590688 61718 590772 61954
rect 591008 61718 592960 61954
rect -9036 61634 592960 61718
rect -9036 61398 -7084 61634
rect -6848 61398 -6764 61634
rect -6528 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590452 61634
rect 590688 61398 590772 61634
rect 591008 61398 592960 61634
rect -9036 61366 592960 61398
rect -9036 57454 592960 57486
rect -9036 57218 -6124 57454
rect -5888 57218 -5804 57454
rect -5568 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589492 57454
rect 589728 57218 589812 57454
rect 590048 57218 592960 57454
rect -9036 57134 592960 57218
rect -9036 56898 -6124 57134
rect -5888 56898 -5804 57134
rect -5568 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589492 57134
rect 589728 56898 589812 57134
rect 590048 56898 592960 57134
rect -9036 56866 592960 56898
rect -9036 52954 592960 52986
rect -9036 52718 -5164 52954
rect -4928 52718 -4844 52954
rect -4608 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588532 52954
rect 588768 52718 588852 52954
rect 589088 52718 592960 52954
rect -9036 52634 592960 52718
rect -9036 52398 -5164 52634
rect -4928 52398 -4844 52634
rect -4608 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588532 52634
rect 588768 52398 588852 52634
rect 589088 52398 592960 52634
rect -9036 52366 592960 52398
rect -9036 48454 592960 48486
rect -9036 48218 -4204 48454
rect -3968 48218 -3884 48454
rect -3648 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587572 48454
rect 587808 48218 587892 48454
rect 588128 48218 592960 48454
rect -9036 48134 592960 48218
rect -9036 47898 -4204 48134
rect -3968 47898 -3884 48134
rect -3648 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587572 48134
rect 587808 47898 587892 48134
rect 588128 47898 592960 48134
rect -9036 47866 592960 47898
rect -9036 43954 592960 43986
rect -9036 43718 -3244 43954
rect -3008 43718 -2924 43954
rect -2688 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586612 43954
rect 586848 43718 586932 43954
rect 587168 43718 592960 43954
rect -9036 43634 592960 43718
rect -9036 43398 -3244 43634
rect -3008 43398 -2924 43634
rect -2688 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586612 43634
rect 586848 43398 586932 43634
rect 587168 43398 592960 43634
rect -9036 43366 592960 43398
rect -9036 39454 592960 39486
rect -9036 39218 -2284 39454
rect -2048 39218 -1964 39454
rect -1728 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585652 39454
rect 585888 39218 585972 39454
rect 586208 39218 592960 39454
rect -9036 39134 592960 39218
rect -9036 38898 -2284 39134
rect -2048 38898 -1964 39134
rect -1728 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585652 39134
rect 585888 38898 585972 39134
rect 586208 38898 592960 39134
rect -9036 38866 592960 38898
rect -9036 34954 592960 34986
rect -9036 34718 -9004 34954
rect -8768 34718 -8684 34954
rect -8448 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592372 34954
rect 592608 34718 592692 34954
rect 592928 34718 592960 34954
rect -9036 34634 592960 34718
rect -9036 34398 -9004 34634
rect -8768 34398 -8684 34634
rect -8448 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592372 34634
rect 592608 34398 592692 34634
rect 592928 34398 592960 34634
rect -9036 34366 592960 34398
rect -9036 30454 592960 30486
rect -9036 30218 -8044 30454
rect -7808 30218 -7724 30454
rect -7488 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591412 30454
rect 591648 30218 591732 30454
rect 591968 30218 592960 30454
rect -9036 30134 592960 30218
rect -9036 29898 -8044 30134
rect -7808 29898 -7724 30134
rect -7488 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591412 30134
rect 591648 29898 591732 30134
rect 591968 29898 592960 30134
rect -9036 29866 592960 29898
rect -9036 25954 592960 25986
rect -9036 25718 -7084 25954
rect -6848 25718 -6764 25954
rect -6528 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590452 25954
rect 590688 25718 590772 25954
rect 591008 25718 592960 25954
rect -9036 25634 592960 25718
rect -9036 25398 -7084 25634
rect -6848 25398 -6764 25634
rect -6528 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590452 25634
rect 590688 25398 590772 25634
rect 591008 25398 592960 25634
rect -9036 25366 592960 25398
rect -9036 21454 592960 21486
rect -9036 21218 -6124 21454
rect -5888 21218 -5804 21454
rect -5568 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589492 21454
rect 589728 21218 589812 21454
rect 590048 21218 592960 21454
rect -9036 21134 592960 21218
rect -9036 20898 -6124 21134
rect -5888 20898 -5804 21134
rect -5568 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589492 21134
rect 589728 20898 589812 21134
rect 590048 20898 592960 21134
rect -9036 20866 592960 20898
rect -9036 16954 592960 16986
rect -9036 16718 -5164 16954
rect -4928 16718 -4844 16954
rect -4608 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588532 16954
rect 588768 16718 588852 16954
rect 589088 16718 592960 16954
rect -9036 16634 592960 16718
rect -9036 16398 -5164 16634
rect -4928 16398 -4844 16634
rect -4608 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588532 16634
rect 588768 16398 588852 16634
rect 589088 16398 592960 16634
rect -9036 16366 592960 16398
rect -9036 12454 592960 12486
rect -9036 12218 -4204 12454
rect -3968 12218 -3884 12454
rect -3648 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587572 12454
rect 587808 12218 587892 12454
rect 588128 12218 592960 12454
rect -9036 12134 592960 12218
rect -9036 11898 -4204 12134
rect -3968 11898 -3884 12134
rect -3648 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587572 12134
rect 587808 11898 587892 12134
rect 588128 11898 592960 12134
rect -9036 11866 592960 11898
rect -9036 7954 592960 7986
rect -9036 7718 -3244 7954
rect -3008 7718 -2924 7954
rect -2688 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586612 7954
rect 586848 7718 586932 7954
rect 587168 7718 592960 7954
rect -9036 7634 592960 7718
rect -9036 7398 -3244 7634
rect -3008 7398 -2924 7634
rect -2688 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586612 7634
rect 586848 7398 586932 7634
rect 587168 7398 592960 7634
rect -9036 7366 592960 7398
rect -9036 3454 592960 3486
rect -9036 3218 -2284 3454
rect -2048 3218 -1964 3454
rect -1728 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585652 3454
rect 585888 3218 585972 3454
rect 586208 3218 592960 3454
rect -9036 3134 592960 3218
rect -9036 2898 -2284 3134
rect -2048 2898 -1964 3134
rect -1728 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585652 3134
rect 585888 2898 585972 3134
rect 586208 2898 592960 3134
rect -9036 2866 592960 2898
rect -2316 -656 586240 -624
rect -2316 -892 -2284 -656
rect -2048 -892 -1964 -656
rect -1728 -892 1826 -656
rect 2062 -892 2146 -656
rect 2382 -892 37826 -656
rect 38062 -892 38146 -656
rect 38382 -892 73826 -656
rect 74062 -892 74146 -656
rect 74382 -892 109826 -656
rect 110062 -892 110146 -656
rect 110382 -892 145826 -656
rect 146062 -892 146146 -656
rect 146382 -892 181826 -656
rect 182062 -892 182146 -656
rect 182382 -892 217826 -656
rect 218062 -892 218146 -656
rect 218382 -892 253826 -656
rect 254062 -892 254146 -656
rect 254382 -892 289826 -656
rect 290062 -892 290146 -656
rect 290382 -892 325826 -656
rect 326062 -892 326146 -656
rect 326382 -892 361826 -656
rect 362062 -892 362146 -656
rect 362382 -892 397826 -656
rect 398062 -892 398146 -656
rect 398382 -892 433826 -656
rect 434062 -892 434146 -656
rect 434382 -892 469826 -656
rect 470062 -892 470146 -656
rect 470382 -892 505826 -656
rect 506062 -892 506146 -656
rect 506382 -892 541826 -656
rect 542062 -892 542146 -656
rect 542382 -892 577826 -656
rect 578062 -892 578146 -656
rect 578382 -892 585652 -656
rect 585888 -892 585972 -656
rect 586208 -892 586240 -656
rect -2316 -976 586240 -892
rect -2316 -1212 -2284 -976
rect -2048 -1212 -1964 -976
rect -1728 -1212 1826 -976
rect 2062 -1212 2146 -976
rect 2382 -1212 37826 -976
rect 38062 -1212 38146 -976
rect 38382 -1212 73826 -976
rect 74062 -1212 74146 -976
rect 74382 -1212 109826 -976
rect 110062 -1212 110146 -976
rect 110382 -1212 145826 -976
rect 146062 -1212 146146 -976
rect 146382 -1212 181826 -976
rect 182062 -1212 182146 -976
rect 182382 -1212 217826 -976
rect 218062 -1212 218146 -976
rect 218382 -1212 253826 -976
rect 254062 -1212 254146 -976
rect 254382 -1212 289826 -976
rect 290062 -1212 290146 -976
rect 290382 -1212 325826 -976
rect 326062 -1212 326146 -976
rect 326382 -1212 361826 -976
rect 362062 -1212 362146 -976
rect 362382 -1212 397826 -976
rect 398062 -1212 398146 -976
rect 398382 -1212 433826 -976
rect 434062 -1212 434146 -976
rect 434382 -1212 469826 -976
rect 470062 -1212 470146 -976
rect 470382 -1212 505826 -976
rect 506062 -1212 506146 -976
rect 506382 -1212 541826 -976
rect 542062 -1212 542146 -976
rect 542382 -1212 577826 -976
rect 578062 -1212 578146 -976
rect 578382 -1212 585652 -976
rect 585888 -1212 585972 -976
rect 586208 -1212 586240 -976
rect -2316 -1244 586240 -1212
rect -3276 -1616 587200 -1584
rect -3276 -1852 -3244 -1616
rect -3008 -1852 -2924 -1616
rect -2688 -1852 6326 -1616
rect 6562 -1852 6646 -1616
rect 6882 -1852 42326 -1616
rect 42562 -1852 42646 -1616
rect 42882 -1852 78326 -1616
rect 78562 -1852 78646 -1616
rect 78882 -1852 114326 -1616
rect 114562 -1852 114646 -1616
rect 114882 -1852 150326 -1616
rect 150562 -1852 150646 -1616
rect 150882 -1852 186326 -1616
rect 186562 -1852 186646 -1616
rect 186882 -1852 222326 -1616
rect 222562 -1852 222646 -1616
rect 222882 -1852 258326 -1616
rect 258562 -1852 258646 -1616
rect 258882 -1852 294326 -1616
rect 294562 -1852 294646 -1616
rect 294882 -1852 330326 -1616
rect 330562 -1852 330646 -1616
rect 330882 -1852 366326 -1616
rect 366562 -1852 366646 -1616
rect 366882 -1852 402326 -1616
rect 402562 -1852 402646 -1616
rect 402882 -1852 438326 -1616
rect 438562 -1852 438646 -1616
rect 438882 -1852 474326 -1616
rect 474562 -1852 474646 -1616
rect 474882 -1852 510326 -1616
rect 510562 -1852 510646 -1616
rect 510882 -1852 546326 -1616
rect 546562 -1852 546646 -1616
rect 546882 -1852 582326 -1616
rect 582562 -1852 582646 -1616
rect 582882 -1852 586612 -1616
rect 586848 -1852 586932 -1616
rect 587168 -1852 587200 -1616
rect -3276 -1936 587200 -1852
rect -3276 -2172 -3244 -1936
rect -3008 -2172 -2924 -1936
rect -2688 -2172 6326 -1936
rect 6562 -2172 6646 -1936
rect 6882 -2172 42326 -1936
rect 42562 -2172 42646 -1936
rect 42882 -2172 78326 -1936
rect 78562 -2172 78646 -1936
rect 78882 -2172 114326 -1936
rect 114562 -2172 114646 -1936
rect 114882 -2172 150326 -1936
rect 150562 -2172 150646 -1936
rect 150882 -2172 186326 -1936
rect 186562 -2172 186646 -1936
rect 186882 -2172 222326 -1936
rect 222562 -2172 222646 -1936
rect 222882 -2172 258326 -1936
rect 258562 -2172 258646 -1936
rect 258882 -2172 294326 -1936
rect 294562 -2172 294646 -1936
rect 294882 -2172 330326 -1936
rect 330562 -2172 330646 -1936
rect 330882 -2172 366326 -1936
rect 366562 -2172 366646 -1936
rect 366882 -2172 402326 -1936
rect 402562 -2172 402646 -1936
rect 402882 -2172 438326 -1936
rect 438562 -2172 438646 -1936
rect 438882 -2172 474326 -1936
rect 474562 -2172 474646 -1936
rect 474882 -2172 510326 -1936
rect 510562 -2172 510646 -1936
rect 510882 -2172 546326 -1936
rect 546562 -2172 546646 -1936
rect 546882 -2172 582326 -1936
rect 582562 -2172 582646 -1936
rect 582882 -2172 586612 -1936
rect 586848 -2172 586932 -1936
rect 587168 -2172 587200 -1936
rect -3276 -2204 587200 -2172
rect -4236 -2576 588160 -2544
rect -4236 -2812 -4204 -2576
rect -3968 -2812 -3884 -2576
rect -3648 -2812 10826 -2576
rect 11062 -2812 11146 -2576
rect 11382 -2812 46826 -2576
rect 47062 -2812 47146 -2576
rect 47382 -2812 82826 -2576
rect 83062 -2812 83146 -2576
rect 83382 -2812 118826 -2576
rect 119062 -2812 119146 -2576
rect 119382 -2812 154826 -2576
rect 155062 -2812 155146 -2576
rect 155382 -2812 190826 -2576
rect 191062 -2812 191146 -2576
rect 191382 -2812 226826 -2576
rect 227062 -2812 227146 -2576
rect 227382 -2812 262826 -2576
rect 263062 -2812 263146 -2576
rect 263382 -2812 298826 -2576
rect 299062 -2812 299146 -2576
rect 299382 -2812 334826 -2576
rect 335062 -2812 335146 -2576
rect 335382 -2812 370826 -2576
rect 371062 -2812 371146 -2576
rect 371382 -2812 406826 -2576
rect 407062 -2812 407146 -2576
rect 407382 -2812 442826 -2576
rect 443062 -2812 443146 -2576
rect 443382 -2812 478826 -2576
rect 479062 -2812 479146 -2576
rect 479382 -2812 514826 -2576
rect 515062 -2812 515146 -2576
rect 515382 -2812 550826 -2576
rect 551062 -2812 551146 -2576
rect 551382 -2812 587572 -2576
rect 587808 -2812 587892 -2576
rect 588128 -2812 588160 -2576
rect -4236 -2896 588160 -2812
rect -4236 -3132 -4204 -2896
rect -3968 -3132 -3884 -2896
rect -3648 -3132 10826 -2896
rect 11062 -3132 11146 -2896
rect 11382 -3132 46826 -2896
rect 47062 -3132 47146 -2896
rect 47382 -3132 82826 -2896
rect 83062 -3132 83146 -2896
rect 83382 -3132 118826 -2896
rect 119062 -3132 119146 -2896
rect 119382 -3132 154826 -2896
rect 155062 -3132 155146 -2896
rect 155382 -3132 190826 -2896
rect 191062 -3132 191146 -2896
rect 191382 -3132 226826 -2896
rect 227062 -3132 227146 -2896
rect 227382 -3132 262826 -2896
rect 263062 -3132 263146 -2896
rect 263382 -3132 298826 -2896
rect 299062 -3132 299146 -2896
rect 299382 -3132 334826 -2896
rect 335062 -3132 335146 -2896
rect 335382 -3132 370826 -2896
rect 371062 -3132 371146 -2896
rect 371382 -3132 406826 -2896
rect 407062 -3132 407146 -2896
rect 407382 -3132 442826 -2896
rect 443062 -3132 443146 -2896
rect 443382 -3132 478826 -2896
rect 479062 -3132 479146 -2896
rect 479382 -3132 514826 -2896
rect 515062 -3132 515146 -2896
rect 515382 -3132 550826 -2896
rect 551062 -3132 551146 -2896
rect 551382 -3132 587572 -2896
rect 587808 -3132 587892 -2896
rect 588128 -3132 588160 -2896
rect -4236 -3164 588160 -3132
rect -5196 -3536 589120 -3504
rect -5196 -3772 -5164 -3536
rect -4928 -3772 -4844 -3536
rect -4608 -3772 15326 -3536
rect 15562 -3772 15646 -3536
rect 15882 -3772 51326 -3536
rect 51562 -3772 51646 -3536
rect 51882 -3772 87326 -3536
rect 87562 -3772 87646 -3536
rect 87882 -3772 123326 -3536
rect 123562 -3772 123646 -3536
rect 123882 -3772 159326 -3536
rect 159562 -3772 159646 -3536
rect 159882 -3772 195326 -3536
rect 195562 -3772 195646 -3536
rect 195882 -3772 231326 -3536
rect 231562 -3772 231646 -3536
rect 231882 -3772 267326 -3536
rect 267562 -3772 267646 -3536
rect 267882 -3772 303326 -3536
rect 303562 -3772 303646 -3536
rect 303882 -3772 339326 -3536
rect 339562 -3772 339646 -3536
rect 339882 -3772 375326 -3536
rect 375562 -3772 375646 -3536
rect 375882 -3772 411326 -3536
rect 411562 -3772 411646 -3536
rect 411882 -3772 447326 -3536
rect 447562 -3772 447646 -3536
rect 447882 -3772 483326 -3536
rect 483562 -3772 483646 -3536
rect 483882 -3772 519326 -3536
rect 519562 -3772 519646 -3536
rect 519882 -3772 555326 -3536
rect 555562 -3772 555646 -3536
rect 555882 -3772 588532 -3536
rect 588768 -3772 588852 -3536
rect 589088 -3772 589120 -3536
rect -5196 -3856 589120 -3772
rect -5196 -4092 -5164 -3856
rect -4928 -4092 -4844 -3856
rect -4608 -4092 15326 -3856
rect 15562 -4092 15646 -3856
rect 15882 -4092 51326 -3856
rect 51562 -4092 51646 -3856
rect 51882 -4092 87326 -3856
rect 87562 -4092 87646 -3856
rect 87882 -4092 123326 -3856
rect 123562 -4092 123646 -3856
rect 123882 -4092 159326 -3856
rect 159562 -4092 159646 -3856
rect 159882 -4092 195326 -3856
rect 195562 -4092 195646 -3856
rect 195882 -4092 231326 -3856
rect 231562 -4092 231646 -3856
rect 231882 -4092 267326 -3856
rect 267562 -4092 267646 -3856
rect 267882 -4092 303326 -3856
rect 303562 -4092 303646 -3856
rect 303882 -4092 339326 -3856
rect 339562 -4092 339646 -3856
rect 339882 -4092 375326 -3856
rect 375562 -4092 375646 -3856
rect 375882 -4092 411326 -3856
rect 411562 -4092 411646 -3856
rect 411882 -4092 447326 -3856
rect 447562 -4092 447646 -3856
rect 447882 -4092 483326 -3856
rect 483562 -4092 483646 -3856
rect 483882 -4092 519326 -3856
rect 519562 -4092 519646 -3856
rect 519882 -4092 555326 -3856
rect 555562 -4092 555646 -3856
rect 555882 -4092 588532 -3856
rect 588768 -4092 588852 -3856
rect 589088 -4092 589120 -3856
rect -5196 -4124 589120 -4092
rect -6156 -4496 590080 -4464
rect -6156 -4732 -6124 -4496
rect -5888 -4732 -5804 -4496
rect -5568 -4732 19826 -4496
rect 20062 -4732 20146 -4496
rect 20382 -4732 55826 -4496
rect 56062 -4732 56146 -4496
rect 56382 -4732 91826 -4496
rect 92062 -4732 92146 -4496
rect 92382 -4732 127826 -4496
rect 128062 -4732 128146 -4496
rect 128382 -4732 163826 -4496
rect 164062 -4732 164146 -4496
rect 164382 -4732 199826 -4496
rect 200062 -4732 200146 -4496
rect 200382 -4732 235826 -4496
rect 236062 -4732 236146 -4496
rect 236382 -4732 271826 -4496
rect 272062 -4732 272146 -4496
rect 272382 -4732 307826 -4496
rect 308062 -4732 308146 -4496
rect 308382 -4732 343826 -4496
rect 344062 -4732 344146 -4496
rect 344382 -4732 379826 -4496
rect 380062 -4732 380146 -4496
rect 380382 -4732 415826 -4496
rect 416062 -4732 416146 -4496
rect 416382 -4732 451826 -4496
rect 452062 -4732 452146 -4496
rect 452382 -4732 487826 -4496
rect 488062 -4732 488146 -4496
rect 488382 -4732 523826 -4496
rect 524062 -4732 524146 -4496
rect 524382 -4732 559826 -4496
rect 560062 -4732 560146 -4496
rect 560382 -4732 589492 -4496
rect 589728 -4732 589812 -4496
rect 590048 -4732 590080 -4496
rect -6156 -4816 590080 -4732
rect -6156 -5052 -6124 -4816
rect -5888 -5052 -5804 -4816
rect -5568 -5052 19826 -4816
rect 20062 -5052 20146 -4816
rect 20382 -5052 55826 -4816
rect 56062 -5052 56146 -4816
rect 56382 -5052 91826 -4816
rect 92062 -5052 92146 -4816
rect 92382 -5052 127826 -4816
rect 128062 -5052 128146 -4816
rect 128382 -5052 163826 -4816
rect 164062 -5052 164146 -4816
rect 164382 -5052 199826 -4816
rect 200062 -5052 200146 -4816
rect 200382 -5052 235826 -4816
rect 236062 -5052 236146 -4816
rect 236382 -5052 271826 -4816
rect 272062 -5052 272146 -4816
rect 272382 -5052 307826 -4816
rect 308062 -5052 308146 -4816
rect 308382 -5052 343826 -4816
rect 344062 -5052 344146 -4816
rect 344382 -5052 379826 -4816
rect 380062 -5052 380146 -4816
rect 380382 -5052 415826 -4816
rect 416062 -5052 416146 -4816
rect 416382 -5052 451826 -4816
rect 452062 -5052 452146 -4816
rect 452382 -5052 487826 -4816
rect 488062 -5052 488146 -4816
rect 488382 -5052 523826 -4816
rect 524062 -5052 524146 -4816
rect 524382 -5052 559826 -4816
rect 560062 -5052 560146 -4816
rect 560382 -5052 589492 -4816
rect 589728 -5052 589812 -4816
rect 590048 -5052 590080 -4816
rect -6156 -5084 590080 -5052
rect -7116 -5456 591040 -5424
rect -7116 -5692 -7084 -5456
rect -6848 -5692 -6764 -5456
rect -6528 -5692 24326 -5456
rect 24562 -5692 24646 -5456
rect 24882 -5692 60326 -5456
rect 60562 -5692 60646 -5456
rect 60882 -5692 96326 -5456
rect 96562 -5692 96646 -5456
rect 96882 -5692 132326 -5456
rect 132562 -5692 132646 -5456
rect 132882 -5692 168326 -5456
rect 168562 -5692 168646 -5456
rect 168882 -5692 204326 -5456
rect 204562 -5692 204646 -5456
rect 204882 -5692 240326 -5456
rect 240562 -5692 240646 -5456
rect 240882 -5692 276326 -5456
rect 276562 -5692 276646 -5456
rect 276882 -5692 312326 -5456
rect 312562 -5692 312646 -5456
rect 312882 -5692 348326 -5456
rect 348562 -5692 348646 -5456
rect 348882 -5692 384326 -5456
rect 384562 -5692 384646 -5456
rect 384882 -5692 420326 -5456
rect 420562 -5692 420646 -5456
rect 420882 -5692 456326 -5456
rect 456562 -5692 456646 -5456
rect 456882 -5692 492326 -5456
rect 492562 -5692 492646 -5456
rect 492882 -5692 528326 -5456
rect 528562 -5692 528646 -5456
rect 528882 -5692 564326 -5456
rect 564562 -5692 564646 -5456
rect 564882 -5692 590452 -5456
rect 590688 -5692 590772 -5456
rect 591008 -5692 591040 -5456
rect -7116 -5776 591040 -5692
rect -7116 -6012 -7084 -5776
rect -6848 -6012 -6764 -5776
rect -6528 -6012 24326 -5776
rect 24562 -6012 24646 -5776
rect 24882 -6012 60326 -5776
rect 60562 -6012 60646 -5776
rect 60882 -6012 96326 -5776
rect 96562 -6012 96646 -5776
rect 96882 -6012 132326 -5776
rect 132562 -6012 132646 -5776
rect 132882 -6012 168326 -5776
rect 168562 -6012 168646 -5776
rect 168882 -6012 204326 -5776
rect 204562 -6012 204646 -5776
rect 204882 -6012 240326 -5776
rect 240562 -6012 240646 -5776
rect 240882 -6012 276326 -5776
rect 276562 -6012 276646 -5776
rect 276882 -6012 312326 -5776
rect 312562 -6012 312646 -5776
rect 312882 -6012 348326 -5776
rect 348562 -6012 348646 -5776
rect 348882 -6012 384326 -5776
rect 384562 -6012 384646 -5776
rect 384882 -6012 420326 -5776
rect 420562 -6012 420646 -5776
rect 420882 -6012 456326 -5776
rect 456562 -6012 456646 -5776
rect 456882 -6012 492326 -5776
rect 492562 -6012 492646 -5776
rect 492882 -6012 528326 -5776
rect 528562 -6012 528646 -5776
rect 528882 -6012 564326 -5776
rect 564562 -6012 564646 -5776
rect 564882 -6012 590452 -5776
rect 590688 -6012 590772 -5776
rect 591008 -6012 591040 -5776
rect -7116 -6044 591040 -6012
rect -8076 -6416 592000 -6384
rect -8076 -6652 -8044 -6416
rect -7808 -6652 -7724 -6416
rect -7488 -6652 28826 -6416
rect 29062 -6652 29146 -6416
rect 29382 -6652 64826 -6416
rect 65062 -6652 65146 -6416
rect 65382 -6652 100826 -6416
rect 101062 -6652 101146 -6416
rect 101382 -6652 136826 -6416
rect 137062 -6652 137146 -6416
rect 137382 -6652 172826 -6416
rect 173062 -6652 173146 -6416
rect 173382 -6652 208826 -6416
rect 209062 -6652 209146 -6416
rect 209382 -6652 244826 -6416
rect 245062 -6652 245146 -6416
rect 245382 -6652 280826 -6416
rect 281062 -6652 281146 -6416
rect 281382 -6652 316826 -6416
rect 317062 -6652 317146 -6416
rect 317382 -6652 352826 -6416
rect 353062 -6652 353146 -6416
rect 353382 -6652 388826 -6416
rect 389062 -6652 389146 -6416
rect 389382 -6652 424826 -6416
rect 425062 -6652 425146 -6416
rect 425382 -6652 460826 -6416
rect 461062 -6652 461146 -6416
rect 461382 -6652 496826 -6416
rect 497062 -6652 497146 -6416
rect 497382 -6652 532826 -6416
rect 533062 -6652 533146 -6416
rect 533382 -6652 568826 -6416
rect 569062 -6652 569146 -6416
rect 569382 -6652 591412 -6416
rect 591648 -6652 591732 -6416
rect 591968 -6652 592000 -6416
rect -8076 -6736 592000 -6652
rect -8076 -6972 -8044 -6736
rect -7808 -6972 -7724 -6736
rect -7488 -6972 28826 -6736
rect 29062 -6972 29146 -6736
rect 29382 -6972 64826 -6736
rect 65062 -6972 65146 -6736
rect 65382 -6972 100826 -6736
rect 101062 -6972 101146 -6736
rect 101382 -6972 136826 -6736
rect 137062 -6972 137146 -6736
rect 137382 -6972 172826 -6736
rect 173062 -6972 173146 -6736
rect 173382 -6972 208826 -6736
rect 209062 -6972 209146 -6736
rect 209382 -6972 244826 -6736
rect 245062 -6972 245146 -6736
rect 245382 -6972 280826 -6736
rect 281062 -6972 281146 -6736
rect 281382 -6972 316826 -6736
rect 317062 -6972 317146 -6736
rect 317382 -6972 352826 -6736
rect 353062 -6972 353146 -6736
rect 353382 -6972 388826 -6736
rect 389062 -6972 389146 -6736
rect 389382 -6972 424826 -6736
rect 425062 -6972 425146 -6736
rect 425382 -6972 460826 -6736
rect 461062 -6972 461146 -6736
rect 461382 -6972 496826 -6736
rect 497062 -6972 497146 -6736
rect 497382 -6972 532826 -6736
rect 533062 -6972 533146 -6736
rect 533382 -6972 568826 -6736
rect 569062 -6972 569146 -6736
rect 569382 -6972 591412 -6736
rect 591648 -6972 591732 -6736
rect 591968 -6972 592000 -6736
rect -8076 -7004 592000 -6972
rect -9036 -7376 592960 -7344
rect -9036 -7612 -9004 -7376
rect -8768 -7612 -8684 -7376
rect -8448 -7612 33326 -7376
rect 33562 -7612 33646 -7376
rect 33882 -7612 69326 -7376
rect 69562 -7612 69646 -7376
rect 69882 -7612 105326 -7376
rect 105562 -7612 105646 -7376
rect 105882 -7612 141326 -7376
rect 141562 -7612 141646 -7376
rect 141882 -7612 177326 -7376
rect 177562 -7612 177646 -7376
rect 177882 -7612 213326 -7376
rect 213562 -7612 213646 -7376
rect 213882 -7612 249326 -7376
rect 249562 -7612 249646 -7376
rect 249882 -7612 285326 -7376
rect 285562 -7612 285646 -7376
rect 285882 -7612 321326 -7376
rect 321562 -7612 321646 -7376
rect 321882 -7612 357326 -7376
rect 357562 -7612 357646 -7376
rect 357882 -7612 393326 -7376
rect 393562 -7612 393646 -7376
rect 393882 -7612 429326 -7376
rect 429562 -7612 429646 -7376
rect 429882 -7612 465326 -7376
rect 465562 -7612 465646 -7376
rect 465882 -7612 501326 -7376
rect 501562 -7612 501646 -7376
rect 501882 -7612 537326 -7376
rect 537562 -7612 537646 -7376
rect 537882 -7612 573326 -7376
rect 573562 -7612 573646 -7376
rect 573882 -7612 592372 -7376
rect 592608 -7612 592692 -7376
rect 592928 -7612 592960 -7376
rect -9036 -7696 592960 -7612
rect -9036 -7932 -9004 -7696
rect -8768 -7932 -8684 -7696
rect -8448 -7932 33326 -7696
rect 33562 -7932 33646 -7696
rect 33882 -7932 69326 -7696
rect 69562 -7932 69646 -7696
rect 69882 -7932 105326 -7696
rect 105562 -7932 105646 -7696
rect 105882 -7932 141326 -7696
rect 141562 -7932 141646 -7696
rect 141882 -7932 177326 -7696
rect 177562 -7932 177646 -7696
rect 177882 -7932 213326 -7696
rect 213562 -7932 213646 -7696
rect 213882 -7932 249326 -7696
rect 249562 -7932 249646 -7696
rect 249882 -7932 285326 -7696
rect 285562 -7932 285646 -7696
rect 285882 -7932 321326 -7696
rect 321562 -7932 321646 -7696
rect 321882 -7932 357326 -7696
rect 357562 -7932 357646 -7696
rect 357882 -7932 393326 -7696
rect 393562 -7932 393646 -7696
rect 393882 -7932 429326 -7696
rect 429562 -7932 429646 -7696
rect 429882 -7932 465326 -7696
rect 465562 -7932 465646 -7696
rect 465882 -7932 501326 -7696
rect 501562 -7932 501646 -7696
rect 501882 -7932 537326 -7696
rect 537562 -7932 537646 -7696
rect 537882 -7932 573326 -7696
rect 573562 -7932 573646 -7696
rect 573882 -7932 592372 -7696
rect 592608 -7932 592692 -7696
rect 592928 -7932 592960 -7696
rect -9036 -7964 592960 -7932
use sky130_sram_2kbyte_1rw1r_32x512_8  dram_inst
timestamp 0
transform 1 0 220000 0 1 480000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  iram_inst
timestamp 0
transform 1 0 220000 0 1 160000
box 0 0 136620 83308
use rvj1_caravel_soc  rvj1_soc
timestamp 0
transform 1 0 232400 0 1 310400
box 13 0 119678 121902
use wbuart_wrap  uart_inst
timestamp 0
transform 1 0 100000 0 1 300000
box 0 0 70020 72164
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal4 s -2316 -1244 -1696 705180 4 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2316 -1244 586240 -624 8 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2316 704560 586240 705180 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 585620 -1244 586240 705180 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 1794 -7964 2414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 37794 -7964 38414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 73794 -7964 74414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 109794 -7964 110414 298000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 109794 374164 110414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 145794 -7964 146414 298000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 145794 374164 146414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 181794 -7964 182414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 217794 -7964 218414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 217794 245308 218414 478000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 217794 565308 218414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 253794 -7964 254414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 253794 245308 254414 308400 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 253794 434302 254414 478000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 253794 565308 254414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 289794 -7964 290414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 289794 245308 290414 308400 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 289794 434302 290414 478000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 289794 565308 290414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 -7964 326414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 245308 326414 308400 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 434302 326414 478000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 565308 326414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 361794 -7964 362414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 397794 -7964 398414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 433794 -7964 434414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 469794 -7964 470414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 505794 -7964 506414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 541794 -7964 542414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 577794 -7964 578414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 2866 592960 3486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 38866 592960 39486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 74866 592960 75486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 110866 592960 111486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 146866 592960 147486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 182866 592960 183486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 218866 592960 219486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 254866 592960 255486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 290866 592960 291486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 326866 592960 327486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 362866 592960 363486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 398866 592960 399486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 434866 592960 435486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 470866 592960 471486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 506866 592960 507486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 542866 592960 543486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 578866 592960 579486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 614866 592960 615486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 650866 592960 651486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 686866 592960 687486 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s -4236 -3164 -3616 707100 4 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -4236 -3164 588160 -2544 8 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -4236 706480 588160 707100 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 587540 -3164 588160 707100 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 10794 -7964 11414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 46794 -7964 47414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 82794 -7964 83414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 118794 -7964 119414 298000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 118794 374164 119414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 154794 -7964 155414 298000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 154794 374164 155414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 190794 -7964 191414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 226794 -7964 227414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 226794 245308 227414 478000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 226794 565308 227414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 262794 -7964 263414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 262794 245308 263414 308400 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 262794 565308 263414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 298794 -7964 299414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 298794 245308 299414 308400 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 298794 565308 299414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 334794 -7964 335414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 334794 245308 335414 308400 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 334794 565308 335414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 370794 -7964 371414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 406794 -7964 407414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 442794 -7964 443414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 478794 -7964 479414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 514794 -7964 515414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 550794 -7964 551414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 11866 592960 12486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 47866 592960 48486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 83866 592960 84486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 119866 592960 120486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 155866 592960 156486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 191866 592960 192486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 227866 592960 228486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 263866 592960 264486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 299866 592960 300486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 335866 592960 336486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 371866 592960 372486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 407866 592960 408486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 443866 592960 444486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 479866 592960 480486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 515866 592960 516486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 551866 592960 552486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 587866 592960 588486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 623866 592960 624486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 659866 592960 660486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 695866 592960 696486 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s -5196 -4124 -4576 708060 4 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -5196 -4124 589120 -3504 8 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -5196 707440 589120 708060 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 588500 -4124 589120 708060 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 15294 -7964 15914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 51294 -7964 51914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 87294 -7964 87914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 123294 -7964 123914 298000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 123294 374164 123914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 159294 -7964 159914 298000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 159294 374164 159914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 195294 -7964 195914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 231294 -7964 231914 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 231294 245308 231914 308400 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 231294 565308 231914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 267294 -7964 267914 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 267294 245308 267914 308400 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 267294 565308 267914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 303294 -7964 303914 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 303294 245308 303914 308400 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 303294 565308 303914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 339294 -7964 339914 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 339294 245308 339914 308400 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 339294 565308 339914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 375294 -7964 375914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 411294 -7964 411914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 447294 -7964 447914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 483294 -7964 483914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 519294 -7964 519914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 555294 -7964 555914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 16366 592960 16986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 52366 592960 52986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 88366 592960 88986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 124366 592960 124986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 160366 592960 160986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 196366 592960 196986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 232366 592960 232986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 268366 592960 268986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 304366 592960 304986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 340366 592960 340986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 376366 592960 376986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 412366 592960 412986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 448366 592960 448986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 484366 592960 484986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 520366 592960 520986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 556366 592960 556986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 592366 592960 592986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 628366 592960 628986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 664366 592960 664986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 700366 592960 700986 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s -6156 -5084 -5536 709020 4 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -6156 -5084 590080 -4464 8 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -6156 708400 590080 709020 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 589460 -5084 590080 709020 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 19794 -7964 20414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 55794 -7964 56414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 91794 -7964 92414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 127794 -7964 128414 298000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 127794 374164 128414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 163794 -7964 164414 298000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 163794 374164 164414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 199794 -7964 200414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 235794 -7964 236414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 235794 565308 236414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 271794 -7964 272414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 271794 565308 272414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 307794 -7964 308414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 307794 565308 308414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 343794 -7964 344414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 343794 565308 344414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 379794 -7964 380414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 415794 -7964 416414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 451794 -7964 452414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 487794 -7964 488414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 523794 -7964 524414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 559794 -7964 560414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 20866 592960 21486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 56866 592960 57486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 92866 592960 93486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 128866 592960 129486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 164866 592960 165486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 200866 592960 201486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 236866 592960 237486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 272866 592960 273486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 308866 592960 309486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 344866 592960 345486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 380866 592960 381486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 416866 592960 417486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 452866 592960 453486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 488866 592960 489486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 524866 592960 525486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 560866 592960 561486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 596866 592960 597486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 632866 592960 633486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 668866 592960 669486 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s -8076 -7004 -7456 710940 4 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8076 -7004 592000 -6384 8 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8076 710320 592000 710940 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 591380 -7004 592000 710940 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 28794 -7964 29414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 64794 -7964 65414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 100794 -7964 101414 298000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 100794 374164 101414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 136794 -7964 137414 298000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 136794 374164 137414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 172794 -7964 173414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 208794 -7964 209414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 244794 -7964 245414 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 244794 245308 245414 308400 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 244794 565308 245414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 280794 -7964 281414 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 280794 245308 281414 308400 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 280794 565308 281414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 316794 -7964 317414 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 316794 245308 317414 308400 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 316794 565308 317414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 352794 -7964 353414 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 352794 245308 353414 308400 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 352794 565308 353414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 388794 -7964 389414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 424794 -7964 425414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 460794 -7964 461414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 496794 -7964 497414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 532794 -7964 533414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 568794 -7964 569414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 29866 592960 30486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 65866 592960 66486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 101866 592960 102486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 137866 592960 138486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 173866 592960 174486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 209866 592960 210486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 245866 592960 246486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 281866 592960 282486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 317866 592960 318486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 353866 592960 354486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 389866 592960 390486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 425866 592960 426486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 461866 592960 462486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 497866 592960 498486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 533866 592960 534486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 569866 592960 570486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 605866 592960 606486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 641866 592960 642486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 677866 592960 678486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s -9036 -7964 -8416 711900 4 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 -7964 592960 -7344 8 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 711280 592960 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 592340 -7964 592960 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 33294 -7964 33914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 69294 -7964 69914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 105294 -7964 105914 298000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 105294 374164 105914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 141294 -7964 141914 298000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 141294 374164 141914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 177294 -7964 177914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 213294 -7964 213914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 249294 -7964 249914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 249294 245308 249914 308400 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 249294 565308 249914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 285294 -7964 285914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 285294 245308 285914 308400 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 285294 565308 285914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 321294 -7964 321914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 321294 245308 321914 308400 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 321294 565308 321914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 357294 -7964 357914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 357294 245308 357914 478000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 357294 565308 357914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 393294 -7964 393914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 429294 -7964 429914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 465294 -7964 465914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 501294 -7964 501914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 537294 -7964 537914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 573294 -7964 573914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 34366 592960 34986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 70366 592960 70986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 106366 592960 106986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 142366 592960 142986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 178366 592960 178986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 214366 592960 214986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 250366 592960 250986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 286366 592960 286986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 322366 592960 322986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 358366 592960 358986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 394366 592960 394986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 430366 592960 430986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 466366 592960 466986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 502366 592960 502986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 538366 592960 538986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 574366 592960 574986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 610366 592960 610986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 646366 592960 646986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 682366 592960 682986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s -3276 -2204 -2656 706140 4 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -3276 -2204 587200 -1584 8 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -3276 705520 587200 706140 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 586580 -2204 587200 706140 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 6294 -7964 6914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 42294 -7964 42914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 78294 -7964 78914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 114294 -7964 114914 298000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 114294 374164 114914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 150294 -7964 150914 298000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 150294 374164 150914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 186294 -7964 186914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 222294 -7964 222914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 222294 245308 222914 478000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 222294 565308 222914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 258294 -7964 258914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 258294 245308 258914 308400 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 258294 434302 258914 478000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 258294 565308 258914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 294294 -7964 294914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 294294 245308 294914 308400 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 294294 434302 294914 478000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 294294 565308 294914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 330294 -7964 330914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 330294 245308 330914 308400 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 330294 434302 330914 478000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 330294 565308 330914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 366294 -7964 366914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 402294 -7964 402914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 438294 -7964 438914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 474294 -7964 474914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 510294 -7964 510914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 546294 -7964 546914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 582294 -7964 582914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 7366 592960 7986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 43366 592960 43986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 79366 592960 79986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 115366 592960 115986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 151366 592960 151986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 187366 592960 187986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 223366 592960 223986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 259366 592960 259986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 295366 592960 295986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 331366 592960 331986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 367366 592960 367986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 403366 592960 403986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 439366 592960 439986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 475366 592960 475986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 511366 592960 511986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 547366 592960 547986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 583366 592960 583986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 619366 592960 619986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 655366 592960 655986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 691366 592960 691986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s -7116 -6044 -6496 709980 4 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -7116 -6044 591040 -5424 8 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -7116 709360 591040 709980 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 590420 -6044 591040 709980 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 24294 -7964 24914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 60294 -7964 60914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 96294 -7964 96914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 132294 -7964 132914 298000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 132294 374164 132914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 168294 -7964 168914 298000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 168294 374164 168914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 204294 -7964 204914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 240294 -7964 240914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 240294 565308 240914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 276294 -7964 276914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 276294 565308 276914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 312294 -7964 312914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 312294 565308 312914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 348294 -7964 348914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 348294 565308 348914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 384294 -7964 384914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 420294 -7964 420914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 456294 -7964 456914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 492294 -7964 492914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 528294 -7964 528914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 564294 -7964 564914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 25366 592960 25986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 61366 592960 61986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 97366 592960 97986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 133366 592960 133986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 169366 592960 169986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 205366 592960 205986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 241366 592960 241986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 277366 592960 277986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 313366 592960 313986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 349366 592960 349986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 385366 592960 385986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 421366 592960 421986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 457366 592960 457986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 493366 592960 493986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 529366 592960 529986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 565366 592960 565986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 601366 592960 601986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 637366 592960 637986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 673366 592960 673986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
