magic
tech sky130A
magscale 1 2
timestamp 1654158136
<< obsli1 >>
rect 1104 2159 69276 70193
<< obsm1 >>
rect 14 1844 69630 70224
<< metal2 >>
rect 662 71755 718 72555
rect 3238 71755 3294 72555
rect 5814 71755 5870 72555
rect 8390 71755 8446 72555
rect 10966 71755 11022 72555
rect 13542 71755 13598 72555
rect 16118 71755 16174 72555
rect 18694 71755 18750 72555
rect 21270 71755 21326 72555
rect 23846 71755 23902 72555
rect 26422 71755 26478 72555
rect 28998 71755 29054 72555
rect 31574 71755 31630 72555
rect 34150 71755 34206 72555
rect 36726 71755 36782 72555
rect 39302 71755 39358 72555
rect 41878 71755 41934 72555
rect 44454 71755 44510 72555
rect 47030 71755 47086 72555
rect 49606 71755 49662 72555
rect 52182 71755 52238 72555
rect 54758 71755 54814 72555
rect 57334 71755 57390 72555
rect 59910 71755 59966 72555
rect 62486 71755 62542 72555
rect 65062 71755 65118 72555
rect 67638 71755 67694 72555
rect 18 0 74 800
rect 2594 0 2650 800
rect 5170 0 5226 800
rect 7746 0 7802 800
rect 10322 0 10378 800
rect 12898 0 12954 800
rect 15474 0 15530 800
rect 18050 0 18106 800
rect 20626 0 20682 800
rect 23202 0 23258 800
rect 25778 0 25834 800
rect 28354 0 28410 800
rect 30930 0 30986 800
rect 33506 0 33562 800
rect 36082 0 36138 800
rect 38658 0 38714 800
rect 41234 0 41290 800
rect 43810 0 43866 800
rect 46386 0 46442 800
rect 48962 0 49018 800
rect 51538 0 51594 800
rect 54114 0 54170 800
rect 56690 0 56746 800
rect 59266 0 59322 800
rect 61842 0 61898 800
rect 64418 0 64474 800
rect 66994 0 67050 800
rect 69570 0 69626 800
<< obsm2 >>
rect 20 71699 606 72185
rect 774 71699 3182 72185
rect 3350 71699 5758 72185
rect 5926 71699 8334 72185
rect 8502 71699 10910 72185
rect 11078 71699 13486 72185
rect 13654 71699 16062 72185
rect 16230 71699 18638 72185
rect 18806 71699 21214 72185
rect 21382 71699 23790 72185
rect 23958 71699 26366 72185
rect 26534 71699 28942 72185
rect 29110 71699 31518 72185
rect 31686 71699 34094 72185
rect 34262 71699 36670 72185
rect 36838 71699 39246 72185
rect 39414 71699 41822 72185
rect 41990 71699 44398 72185
rect 44566 71699 46974 72185
rect 47142 71699 49550 72185
rect 49718 71699 52126 72185
rect 52294 71699 54702 72185
rect 54870 71699 57278 72185
rect 57446 71699 59854 72185
rect 60022 71699 62430 72185
rect 62598 71699 65006 72185
rect 65174 71699 67582 72185
rect 67750 71699 69624 72185
rect 20 856 69624 71699
rect 130 734 2538 856
rect 2706 734 5114 856
rect 5282 734 7690 856
rect 7858 734 10266 856
rect 10434 734 12842 856
rect 13010 734 15418 856
rect 15586 734 17994 856
rect 18162 734 20570 856
rect 20738 734 23146 856
rect 23314 734 25722 856
rect 25890 734 28298 856
rect 28466 734 30874 856
rect 31042 734 33450 856
rect 33618 734 36026 856
rect 36194 734 38602 856
rect 38770 734 41178 856
rect 41346 734 43754 856
rect 43922 734 46330 856
rect 46498 734 48906 856
rect 49074 734 51482 856
rect 51650 734 54058 856
rect 54226 734 56634 856
rect 56802 734 59210 856
rect 59378 734 61786 856
rect 61954 734 64362 856
rect 64530 734 66938 856
rect 67106 734 69514 856
<< metal3 >>
rect 69611 72088 70411 72208
rect 0 70728 800 70848
rect 69611 69368 70411 69488
rect 0 68008 800 68128
rect 69611 66648 70411 66768
rect 0 65288 800 65408
rect 69611 63928 70411 64048
rect 0 62568 800 62688
rect 69611 61208 70411 61328
rect 0 59848 800 59968
rect 69611 58488 70411 58608
rect 0 57128 800 57248
rect 69611 55768 70411 55888
rect 0 54408 800 54528
rect 69611 53048 70411 53168
rect 0 51688 800 51808
rect 69611 50328 70411 50448
rect 0 48968 800 49088
rect 69611 47608 70411 47728
rect 0 46248 800 46368
rect 69611 44888 70411 45008
rect 0 43528 800 43648
rect 69611 42168 70411 42288
rect 0 40808 800 40928
rect 69611 39448 70411 39568
rect 0 38088 800 38208
rect 69611 36728 70411 36848
rect 0 35368 800 35488
rect 69611 34008 70411 34128
rect 0 32648 800 32768
rect 69611 31288 70411 31408
rect 0 29928 800 30048
rect 69611 28568 70411 28688
rect 0 27208 800 27328
rect 69611 25848 70411 25968
rect 0 24488 800 24608
rect 69611 23128 70411 23248
rect 0 21768 800 21888
rect 69611 20408 70411 20528
rect 0 19048 800 19168
rect 69611 17688 70411 17808
rect 0 16328 800 16448
rect 69611 14968 70411 15088
rect 0 13608 800 13728
rect 69611 12248 70411 12368
rect 0 10888 800 11008
rect 69611 9528 70411 9648
rect 0 8168 800 8288
rect 69611 6808 70411 6928
rect 0 5448 800 5568
rect 69611 4088 70411 4208
rect 0 2728 800 2848
rect 69611 1368 70411 1488
<< obsm3 >>
rect 800 72008 69531 72181
rect 800 70928 69611 72008
rect 880 70648 69611 70928
rect 800 69568 69611 70648
rect 800 69288 69531 69568
rect 800 68208 69611 69288
rect 880 67928 69611 68208
rect 800 66848 69611 67928
rect 800 66568 69531 66848
rect 800 65488 69611 66568
rect 880 65208 69611 65488
rect 800 64128 69611 65208
rect 800 63848 69531 64128
rect 800 62768 69611 63848
rect 880 62488 69611 62768
rect 800 61408 69611 62488
rect 800 61128 69531 61408
rect 800 60048 69611 61128
rect 880 59768 69611 60048
rect 800 58688 69611 59768
rect 800 58408 69531 58688
rect 800 57328 69611 58408
rect 880 57048 69611 57328
rect 800 55968 69611 57048
rect 800 55688 69531 55968
rect 800 54608 69611 55688
rect 880 54328 69611 54608
rect 800 53248 69611 54328
rect 800 52968 69531 53248
rect 800 51888 69611 52968
rect 880 51608 69611 51888
rect 800 50528 69611 51608
rect 800 50248 69531 50528
rect 800 49168 69611 50248
rect 880 48888 69611 49168
rect 800 47808 69611 48888
rect 800 47528 69531 47808
rect 800 46448 69611 47528
rect 880 46168 69611 46448
rect 800 45088 69611 46168
rect 800 44808 69531 45088
rect 800 43728 69611 44808
rect 880 43448 69611 43728
rect 800 42368 69611 43448
rect 800 42088 69531 42368
rect 800 41008 69611 42088
rect 880 40728 69611 41008
rect 800 39648 69611 40728
rect 800 39368 69531 39648
rect 800 38288 69611 39368
rect 880 38008 69611 38288
rect 800 36928 69611 38008
rect 800 36648 69531 36928
rect 800 35568 69611 36648
rect 880 35288 69611 35568
rect 800 34208 69611 35288
rect 800 33928 69531 34208
rect 800 32848 69611 33928
rect 880 32568 69611 32848
rect 800 31488 69611 32568
rect 800 31208 69531 31488
rect 800 30128 69611 31208
rect 880 29848 69611 30128
rect 800 28768 69611 29848
rect 800 28488 69531 28768
rect 800 27408 69611 28488
rect 880 27128 69611 27408
rect 800 26048 69611 27128
rect 800 25768 69531 26048
rect 800 24688 69611 25768
rect 880 24408 69611 24688
rect 800 23328 69611 24408
rect 800 23048 69531 23328
rect 800 21968 69611 23048
rect 880 21688 69611 21968
rect 800 20608 69611 21688
rect 800 20328 69531 20608
rect 800 19248 69611 20328
rect 880 18968 69611 19248
rect 800 17888 69611 18968
rect 800 17608 69531 17888
rect 800 16528 69611 17608
rect 880 16248 69611 16528
rect 800 15168 69611 16248
rect 800 14888 69531 15168
rect 800 13808 69611 14888
rect 880 13528 69611 13808
rect 800 12448 69611 13528
rect 800 12168 69531 12448
rect 800 11088 69611 12168
rect 880 10808 69611 11088
rect 800 9728 69611 10808
rect 800 9448 69531 9728
rect 800 8368 69611 9448
rect 880 8088 69611 8368
rect 800 7008 69611 8088
rect 800 6728 69531 7008
rect 800 5648 69611 6728
rect 880 5368 69611 5648
rect 800 4288 69611 5368
rect 800 4008 69531 4288
rect 800 2928 69611 4008
rect 880 2648 69611 2928
rect 800 1568 69611 2648
rect 800 1395 69531 1568
<< metal4 >>
rect 4208 2128 4528 70224
rect 19568 2128 19888 70224
rect 34928 2128 35248 70224
rect 50288 2128 50608 70224
rect 65648 2128 65968 70224
<< obsm4 >>
rect 9627 2347 19488 69053
rect 19968 2347 34848 69053
rect 35328 2347 50208 69053
rect 50688 2347 61029 69053
<< labels >>
rlabel metal3 s 69611 50328 70411 50448 6 clk_i
port 1 nsew signal input
rlabel metal2 s 65062 71755 65118 72555 6 rst_i
port 2 nsew signal input
rlabel metal2 s 41878 71755 41934 72555 6 uart_rx_i
port 3 nsew signal input
rlabel metal3 s 0 51688 800 51808 6 uart_tx_o
port 4 nsew signal output
rlabel metal4 s 4208 2128 4528 70224 6 vccd1
port 5 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 70224 6 vccd1
port 5 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 70224 6 vccd1
port 5 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 70224 6 vssd1
port 6 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 70224 6 vssd1
port 6 nsew ground bidirectional
rlabel metal2 s 39302 71755 39358 72555 6 wbs_ack_o
port 7 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 wbs_adr_i[0]
port 8 nsew signal input
rlabel metal3 s 69611 1368 70411 1488 6 wbs_adr_i[10]
port 9 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 wbs_adr_i[11]
port 10 nsew signal input
rlabel metal3 s 69611 61208 70411 61328 6 wbs_adr_i[12]
port 11 nsew signal input
rlabel metal2 s 28998 71755 29054 72555 6 wbs_adr_i[13]
port 12 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 wbs_adr_i[14]
port 13 nsew signal input
rlabel metal2 s 34150 71755 34206 72555 6 wbs_adr_i[15]
port 14 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 wbs_adr_i[16]
port 15 nsew signal input
rlabel metal3 s 69611 25848 70411 25968 6 wbs_adr_i[17]
port 16 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 wbs_adr_i[18]
port 17 nsew signal input
rlabel metal3 s 0 59848 800 59968 6 wbs_adr_i[19]
port 18 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 wbs_adr_i[1]
port 19 nsew signal input
rlabel metal3 s 0 46248 800 46368 6 wbs_adr_i[20]
port 20 nsew signal input
rlabel metal2 s 49606 71755 49662 72555 6 wbs_adr_i[21]
port 21 nsew signal input
rlabel metal2 s 59910 71755 59966 72555 6 wbs_adr_i[22]
port 22 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wbs_adr_i[23]
port 23 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 wbs_adr_i[24]
port 24 nsew signal input
rlabel metal3 s 69611 69368 70411 69488 6 wbs_adr_i[25]
port 25 nsew signal input
rlabel metal3 s 69611 17688 70411 17808 6 wbs_adr_i[26]
port 26 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 wbs_adr_i[27]
port 27 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 wbs_adr_i[28]
port 28 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 wbs_adr_i[29]
port 29 nsew signal input
rlabel metal3 s 69611 14968 70411 15088 6 wbs_adr_i[2]
port 30 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 wbs_adr_i[30]
port 31 nsew signal input
rlabel metal3 s 0 48968 800 49088 6 wbs_adr_i[31]
port 32 nsew signal input
rlabel metal3 s 69611 12248 70411 12368 6 wbs_adr_i[3]
port 33 nsew signal input
rlabel metal2 s 36726 71755 36782 72555 6 wbs_adr_i[4]
port 34 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 wbs_adr_i[5]
port 35 nsew signal input
rlabel metal2 s 44454 71755 44510 72555 6 wbs_adr_i[6]
port 36 nsew signal input
rlabel metal3 s 69611 55768 70411 55888 6 wbs_adr_i[7]
port 37 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 wbs_adr_i[8]
port 38 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 wbs_adr_i[9]
port 39 nsew signal input
rlabel metal3 s 69611 63928 70411 64048 6 wbs_cyc_i
port 40 nsew signal input
rlabel metal3 s 69611 72088 70411 72208 6 wbs_dat_i[0]
port 41 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 wbs_dat_i[10]
port 42 nsew signal input
rlabel metal2 s 21270 71755 21326 72555 6 wbs_dat_i[11]
port 43 nsew signal input
rlabel metal3 s 69611 31288 70411 31408 6 wbs_dat_i[12]
port 44 nsew signal input
rlabel metal2 s 23846 71755 23902 72555 6 wbs_dat_i[13]
port 45 nsew signal input
rlabel metal3 s 69611 58488 70411 58608 6 wbs_dat_i[14]
port 46 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 wbs_dat_i[15]
port 47 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_dat_i[16]
port 48 nsew signal input
rlabel metal2 s 26422 71755 26478 72555 6 wbs_dat_i[17]
port 49 nsew signal input
rlabel metal3 s 69611 4088 70411 4208 6 wbs_dat_i[18]
port 50 nsew signal input
rlabel metal3 s 69611 39448 70411 39568 6 wbs_dat_i[19]
port 51 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_dat_i[1]
port 52 nsew signal input
rlabel metal2 s 16118 71755 16174 72555 6 wbs_dat_i[20]
port 53 nsew signal input
rlabel metal3 s 69611 6808 70411 6928 6 wbs_dat_i[21]
port 54 nsew signal input
rlabel metal3 s 69611 66648 70411 66768 6 wbs_dat_i[22]
port 55 nsew signal input
rlabel metal2 s 57334 71755 57390 72555 6 wbs_dat_i[23]
port 56 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 wbs_dat_i[24]
port 57 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 wbs_dat_i[25]
port 58 nsew signal input
rlabel metal3 s 69611 20408 70411 20528 6 wbs_dat_i[26]
port 59 nsew signal input
rlabel metal2 s 18694 71755 18750 72555 6 wbs_dat_i[27]
port 60 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 wbs_dat_i[28]
port 61 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 wbs_dat_i[29]
port 62 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 wbs_dat_i[2]
port 63 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 wbs_dat_i[30]
port 64 nsew signal input
rlabel metal3 s 0 65288 800 65408 6 wbs_dat_i[31]
port 65 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 wbs_dat_i[3]
port 66 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_dat_i[4]
port 67 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 wbs_dat_i[5]
port 68 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 wbs_dat_i[6]
port 69 nsew signal input
rlabel metal3 s 69611 36728 70411 36848 6 wbs_dat_i[7]
port 70 nsew signal input
rlabel metal3 s 69611 23128 70411 23248 6 wbs_dat_i[8]
port 71 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 wbs_dat_i[9]
port 72 nsew signal input
rlabel metal3 s 0 57128 800 57248 6 wbs_dat_o[0]
port 73 nsew signal output
rlabel metal3 s 0 43528 800 43648 6 wbs_dat_o[10]
port 74 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 wbs_dat_o[11]
port 75 nsew signal output
rlabel metal3 s 69611 28568 70411 28688 6 wbs_dat_o[12]
port 76 nsew signal output
rlabel metal3 s 69611 47608 70411 47728 6 wbs_dat_o[13]
port 77 nsew signal output
rlabel metal2 s 59266 0 59322 800 6 wbs_dat_o[14]
port 78 nsew signal output
rlabel metal3 s 69611 53048 70411 53168 6 wbs_dat_o[15]
port 79 nsew signal output
rlabel metal2 s 5814 71755 5870 72555 6 wbs_dat_o[16]
port 80 nsew signal output
rlabel metal2 s 8390 71755 8446 72555 6 wbs_dat_o[17]
port 81 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 wbs_dat_o[18]
port 82 nsew signal output
rlabel metal2 s 18 0 74 800 6 wbs_dat_o[19]
port 83 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 wbs_dat_o[1]
port 84 nsew signal output
rlabel metal2 s 10966 71755 11022 72555 6 wbs_dat_o[20]
port 85 nsew signal output
rlabel metal2 s 31574 71755 31630 72555 6 wbs_dat_o[21]
port 86 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 wbs_dat_o[22]
port 87 nsew signal output
rlabel metal3 s 0 68008 800 68128 6 wbs_dat_o[23]
port 88 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 wbs_dat_o[24]
port 89 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_o[25]
port 90 nsew signal output
rlabel metal2 s 62486 71755 62542 72555 6 wbs_dat_o[26]
port 91 nsew signal output
rlabel metal2 s 47030 71755 47086 72555 6 wbs_dat_o[27]
port 92 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 wbs_dat_o[28]
port 93 nsew signal output
rlabel metal2 s 67638 71755 67694 72555 6 wbs_dat_o[29]
port 94 nsew signal output
rlabel metal3 s 69611 9528 70411 9648 6 wbs_dat_o[2]
port 95 nsew signal output
rlabel metal2 s 662 71755 718 72555 6 wbs_dat_o[30]
port 96 nsew signal output
rlabel metal3 s 69611 42168 70411 42288 6 wbs_dat_o[31]
port 97 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 wbs_dat_o[3]
port 98 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 wbs_dat_o[4]
port 99 nsew signal output
rlabel metal3 s 0 24488 800 24608 6 wbs_dat_o[5]
port 100 nsew signal output
rlabel metal3 s 69611 44888 70411 45008 6 wbs_dat_o[6]
port 101 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 wbs_dat_o[7]
port 102 nsew signal output
rlabel metal2 s 54758 71755 54814 72555 6 wbs_dat_o[8]
port 103 nsew signal output
rlabel metal2 s 52182 71755 52238 72555 6 wbs_dat_o[9]
port 104 nsew signal output
rlabel metal2 s 3238 71755 3294 72555 6 wbs_sel_i[0]
port 105 nsew signal input
rlabel metal2 s 13542 71755 13598 72555 6 wbs_sel_i[1]
port 106 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 wbs_sel_i[2]
port 107 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 wbs_sel_i[3]
port 108 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 wbs_stb_i
port 109 nsew signal input
rlabel metal3 s 69611 34008 70411 34128 6 wbs_we_i
port 110 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 70411 72555
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 11520518
string GDS_FILE /home/jure/Projekti/rvj1-caravel-soc/openlane/wbuart32/runs/wbuart32/results/signoff/wbuart_wrap.magic.gds
string GDS_START 1116912
<< end >>

