magic
tech sky130A
magscale 1 2
timestamp 1654186225
<< obsli1 >>
rect 1104 2159 129168 130033
<< obsm1 >>
rect 14 348 130166 130416
<< metal2 >>
rect 386 131635 442 132435
rect 1122 131635 1178 132435
rect 1858 131635 1914 132435
rect 2686 131635 2742 132435
rect 3422 131635 3478 132435
rect 4158 131635 4214 132435
rect 4986 131635 5042 132435
rect 5722 131635 5778 132435
rect 6550 131635 6606 132435
rect 7286 131635 7342 132435
rect 8022 131635 8078 132435
rect 8850 131635 8906 132435
rect 9586 131635 9642 132435
rect 10322 131635 10378 132435
rect 11150 131635 11206 132435
rect 11886 131635 11942 132435
rect 12714 131635 12770 132435
rect 13450 131635 13506 132435
rect 14186 131635 14242 132435
rect 15014 131635 15070 132435
rect 15750 131635 15806 132435
rect 16486 131635 16542 132435
rect 17314 131635 17370 132435
rect 18050 131635 18106 132435
rect 18878 131635 18934 132435
rect 19614 131635 19670 132435
rect 20350 131635 20406 132435
rect 21178 131635 21234 132435
rect 21914 131635 21970 132435
rect 22650 131635 22706 132435
rect 23478 131635 23534 132435
rect 24214 131635 24270 132435
rect 25042 131635 25098 132435
rect 25778 131635 25834 132435
rect 26514 131635 26570 132435
rect 27342 131635 27398 132435
rect 28078 131635 28134 132435
rect 28906 131635 28962 132435
rect 29642 131635 29698 132435
rect 30378 131635 30434 132435
rect 31206 131635 31262 132435
rect 31942 131635 31998 132435
rect 32678 131635 32734 132435
rect 33506 131635 33562 132435
rect 34242 131635 34298 132435
rect 35070 131635 35126 132435
rect 35806 131635 35862 132435
rect 36542 131635 36598 132435
rect 37370 131635 37426 132435
rect 38106 131635 38162 132435
rect 38842 131635 38898 132435
rect 39670 131635 39726 132435
rect 40406 131635 40462 132435
rect 41234 131635 41290 132435
rect 41970 131635 42026 132435
rect 42706 131635 42762 132435
rect 43534 131635 43590 132435
rect 44270 131635 44326 132435
rect 45006 131635 45062 132435
rect 45834 131635 45890 132435
rect 46570 131635 46626 132435
rect 47398 131635 47454 132435
rect 48134 131635 48190 132435
rect 48870 131635 48926 132435
rect 49698 131635 49754 132435
rect 50434 131635 50490 132435
rect 51170 131635 51226 132435
rect 51998 131635 52054 132435
rect 52734 131635 52790 132435
rect 53562 131635 53618 132435
rect 54298 131635 54354 132435
rect 55034 131635 55090 132435
rect 55862 131635 55918 132435
rect 56598 131635 56654 132435
rect 57426 131635 57482 132435
rect 58162 131635 58218 132435
rect 58898 131635 58954 132435
rect 59726 131635 59782 132435
rect 60462 131635 60518 132435
rect 61198 131635 61254 132435
rect 62026 131635 62082 132435
rect 62762 131635 62818 132435
rect 63590 131635 63646 132435
rect 64326 131635 64382 132435
rect 65062 131635 65118 132435
rect 65890 131635 65946 132435
rect 66626 131635 66682 132435
rect 67362 131635 67418 132435
rect 68190 131635 68246 132435
rect 68926 131635 68982 132435
rect 69754 131635 69810 132435
rect 70490 131635 70546 132435
rect 71226 131635 71282 132435
rect 72054 131635 72110 132435
rect 72790 131635 72846 132435
rect 73526 131635 73582 132435
rect 74354 131635 74410 132435
rect 75090 131635 75146 132435
rect 75918 131635 75974 132435
rect 76654 131635 76710 132435
rect 77390 131635 77446 132435
rect 78218 131635 78274 132435
rect 78954 131635 79010 132435
rect 79782 131635 79838 132435
rect 80518 131635 80574 132435
rect 81254 131635 81310 132435
rect 82082 131635 82138 132435
rect 82818 131635 82874 132435
rect 83554 131635 83610 132435
rect 84382 131635 84438 132435
rect 85118 131635 85174 132435
rect 85946 131635 86002 132435
rect 86682 131635 86738 132435
rect 87418 131635 87474 132435
rect 88246 131635 88302 132435
rect 88982 131635 89038 132435
rect 89718 131635 89774 132435
rect 90546 131635 90602 132435
rect 91282 131635 91338 132435
rect 92110 131635 92166 132435
rect 92846 131635 92902 132435
rect 93582 131635 93638 132435
rect 94410 131635 94466 132435
rect 95146 131635 95202 132435
rect 95882 131635 95938 132435
rect 96710 131635 96766 132435
rect 97446 131635 97502 132435
rect 98274 131635 98330 132435
rect 99010 131635 99066 132435
rect 99746 131635 99802 132435
rect 100574 131635 100630 132435
rect 101310 131635 101366 132435
rect 102046 131635 102102 132435
rect 102874 131635 102930 132435
rect 103610 131635 103666 132435
rect 104438 131635 104494 132435
rect 105174 131635 105230 132435
rect 105910 131635 105966 132435
rect 106738 131635 106794 132435
rect 107474 131635 107530 132435
rect 108302 131635 108358 132435
rect 109038 131635 109094 132435
rect 109774 131635 109830 132435
rect 110602 131635 110658 132435
rect 111338 131635 111394 132435
rect 112074 131635 112130 132435
rect 112902 131635 112958 132435
rect 113638 131635 113694 132435
rect 114466 131635 114522 132435
rect 115202 131635 115258 132435
rect 115938 131635 115994 132435
rect 116766 131635 116822 132435
rect 117502 131635 117558 132435
rect 118238 131635 118294 132435
rect 119066 131635 119122 132435
rect 119802 131635 119858 132435
rect 120630 131635 120686 132435
rect 121366 131635 121422 132435
rect 122102 131635 122158 132435
rect 122930 131635 122986 132435
rect 123666 131635 123722 132435
rect 124402 131635 124458 132435
rect 125230 131635 125286 132435
rect 125966 131635 126022 132435
rect 126794 131635 126850 132435
rect 127530 131635 127586 132435
rect 128266 131635 128322 132435
rect 129094 131635 129150 132435
rect 129830 131635 129886 132435
rect 110 0 166 800
rect 294 0 350 800
rect 478 0 534 800
rect 754 0 810 800
rect 938 0 994 800
rect 1214 0 1270 800
rect 1398 0 1454 800
rect 1674 0 1730 800
rect 1858 0 1914 800
rect 2134 0 2190 800
rect 2318 0 2374 800
rect 2594 0 2650 800
rect 2778 0 2834 800
rect 3054 0 3110 800
rect 3238 0 3294 800
rect 3514 0 3570 800
rect 3698 0 3754 800
rect 3974 0 4030 800
rect 4158 0 4214 800
rect 4434 0 4490 800
rect 4618 0 4674 800
rect 4894 0 4950 800
rect 5078 0 5134 800
rect 5354 0 5410 800
rect 5538 0 5594 800
rect 5814 0 5870 800
rect 5998 0 6054 800
rect 6274 0 6330 800
rect 6458 0 6514 800
rect 6734 0 6790 800
rect 6918 0 6974 800
rect 7194 0 7250 800
rect 7378 0 7434 800
rect 7562 0 7618 800
rect 7838 0 7894 800
rect 8022 0 8078 800
rect 8298 0 8354 800
rect 8482 0 8538 800
rect 8758 0 8814 800
rect 8942 0 8998 800
rect 9218 0 9274 800
rect 9402 0 9458 800
rect 9678 0 9734 800
rect 9862 0 9918 800
rect 10138 0 10194 800
rect 10322 0 10378 800
rect 10598 0 10654 800
rect 10782 0 10838 800
rect 11058 0 11114 800
rect 11242 0 11298 800
rect 11518 0 11574 800
rect 11702 0 11758 800
rect 11978 0 12034 800
rect 12162 0 12218 800
rect 12438 0 12494 800
rect 12622 0 12678 800
rect 12898 0 12954 800
rect 13082 0 13138 800
rect 13358 0 13414 800
rect 13542 0 13598 800
rect 13818 0 13874 800
rect 14002 0 14058 800
rect 14278 0 14334 800
rect 14462 0 14518 800
rect 14646 0 14702 800
rect 14922 0 14978 800
rect 15106 0 15162 800
rect 15382 0 15438 800
rect 15566 0 15622 800
rect 15842 0 15898 800
rect 16026 0 16082 800
rect 16302 0 16358 800
rect 16486 0 16542 800
rect 16762 0 16818 800
rect 16946 0 17002 800
rect 17222 0 17278 800
rect 17406 0 17462 800
rect 17682 0 17738 800
rect 17866 0 17922 800
rect 18142 0 18198 800
rect 18326 0 18382 800
rect 18602 0 18658 800
rect 18786 0 18842 800
rect 19062 0 19118 800
rect 19246 0 19302 800
rect 19522 0 19578 800
rect 19706 0 19762 800
rect 19982 0 20038 800
rect 20166 0 20222 800
rect 20442 0 20498 800
rect 20626 0 20682 800
rect 20902 0 20958 800
rect 21086 0 21142 800
rect 21362 0 21418 800
rect 21546 0 21602 800
rect 21822 0 21878 800
rect 22006 0 22062 800
rect 22190 0 22246 800
rect 22466 0 22522 800
rect 22650 0 22706 800
rect 22926 0 22982 800
rect 23110 0 23166 800
rect 23386 0 23442 800
rect 23570 0 23626 800
rect 23846 0 23902 800
rect 24030 0 24086 800
rect 24306 0 24362 800
rect 24490 0 24546 800
rect 24766 0 24822 800
rect 24950 0 25006 800
rect 25226 0 25282 800
rect 25410 0 25466 800
rect 25686 0 25742 800
rect 25870 0 25926 800
rect 26146 0 26202 800
rect 26330 0 26386 800
rect 26606 0 26662 800
rect 26790 0 26846 800
rect 27066 0 27122 800
rect 27250 0 27306 800
rect 27526 0 27582 800
rect 27710 0 27766 800
rect 27986 0 28042 800
rect 28170 0 28226 800
rect 28446 0 28502 800
rect 28630 0 28686 800
rect 28906 0 28962 800
rect 29090 0 29146 800
rect 29274 0 29330 800
rect 29550 0 29606 800
rect 29734 0 29790 800
rect 30010 0 30066 800
rect 30194 0 30250 800
rect 30470 0 30526 800
rect 30654 0 30710 800
rect 30930 0 30986 800
rect 31114 0 31170 800
rect 31390 0 31446 800
rect 31574 0 31630 800
rect 31850 0 31906 800
rect 32034 0 32090 800
rect 32310 0 32366 800
rect 32494 0 32550 800
rect 32770 0 32826 800
rect 32954 0 33010 800
rect 33230 0 33286 800
rect 33414 0 33470 800
rect 33690 0 33746 800
rect 33874 0 33930 800
rect 34150 0 34206 800
rect 34334 0 34390 800
rect 34610 0 34666 800
rect 34794 0 34850 800
rect 35070 0 35126 800
rect 35254 0 35310 800
rect 35530 0 35586 800
rect 35714 0 35770 800
rect 35990 0 36046 800
rect 36174 0 36230 800
rect 36358 0 36414 800
rect 36634 0 36690 800
rect 36818 0 36874 800
rect 37094 0 37150 800
rect 37278 0 37334 800
rect 37554 0 37610 800
rect 37738 0 37794 800
rect 38014 0 38070 800
rect 38198 0 38254 800
rect 38474 0 38530 800
rect 38658 0 38714 800
rect 38934 0 38990 800
rect 39118 0 39174 800
rect 39394 0 39450 800
rect 39578 0 39634 800
rect 39854 0 39910 800
rect 40038 0 40094 800
rect 40314 0 40370 800
rect 40498 0 40554 800
rect 40774 0 40830 800
rect 40958 0 41014 800
rect 41234 0 41290 800
rect 41418 0 41474 800
rect 41694 0 41750 800
rect 41878 0 41934 800
rect 42154 0 42210 800
rect 42338 0 42394 800
rect 42614 0 42670 800
rect 42798 0 42854 800
rect 43074 0 43130 800
rect 43258 0 43314 800
rect 43534 0 43590 800
rect 43718 0 43774 800
rect 43902 0 43958 800
rect 44178 0 44234 800
rect 44362 0 44418 800
rect 44638 0 44694 800
rect 44822 0 44878 800
rect 45098 0 45154 800
rect 45282 0 45338 800
rect 45558 0 45614 800
rect 45742 0 45798 800
rect 46018 0 46074 800
rect 46202 0 46258 800
rect 46478 0 46534 800
rect 46662 0 46718 800
rect 46938 0 46994 800
rect 47122 0 47178 800
rect 47398 0 47454 800
rect 47582 0 47638 800
rect 47858 0 47914 800
rect 48042 0 48098 800
rect 48318 0 48374 800
rect 48502 0 48558 800
rect 48778 0 48834 800
rect 48962 0 49018 800
rect 49238 0 49294 800
rect 49422 0 49478 800
rect 49698 0 49754 800
rect 49882 0 49938 800
rect 50158 0 50214 800
rect 50342 0 50398 800
rect 50618 0 50674 800
rect 50802 0 50858 800
rect 50986 0 51042 800
rect 51262 0 51318 800
rect 51446 0 51502 800
rect 51722 0 51778 800
rect 51906 0 51962 800
rect 52182 0 52238 800
rect 52366 0 52422 800
rect 52642 0 52698 800
rect 52826 0 52882 800
rect 53102 0 53158 800
rect 53286 0 53342 800
rect 53562 0 53618 800
rect 53746 0 53802 800
rect 54022 0 54078 800
rect 54206 0 54262 800
rect 54482 0 54538 800
rect 54666 0 54722 800
rect 54942 0 54998 800
rect 55126 0 55182 800
rect 55402 0 55458 800
rect 55586 0 55642 800
rect 55862 0 55918 800
rect 56046 0 56102 800
rect 56322 0 56378 800
rect 56506 0 56562 800
rect 56782 0 56838 800
rect 56966 0 57022 800
rect 57242 0 57298 800
rect 57426 0 57482 800
rect 57702 0 57758 800
rect 57886 0 57942 800
rect 58070 0 58126 800
rect 58346 0 58402 800
rect 58530 0 58586 800
rect 58806 0 58862 800
rect 58990 0 59046 800
rect 59266 0 59322 800
rect 59450 0 59506 800
rect 59726 0 59782 800
rect 59910 0 59966 800
rect 60186 0 60242 800
rect 60370 0 60426 800
rect 60646 0 60702 800
rect 60830 0 60886 800
rect 61106 0 61162 800
rect 61290 0 61346 800
rect 61566 0 61622 800
rect 61750 0 61806 800
rect 62026 0 62082 800
rect 62210 0 62266 800
rect 62486 0 62542 800
rect 62670 0 62726 800
rect 62946 0 63002 800
rect 63130 0 63186 800
rect 63406 0 63462 800
rect 63590 0 63646 800
rect 63866 0 63922 800
rect 64050 0 64106 800
rect 64326 0 64382 800
rect 64510 0 64566 800
rect 64786 0 64842 800
rect 64970 0 65026 800
rect 65246 0 65302 800
rect 65430 0 65486 800
rect 65614 0 65670 800
rect 65890 0 65946 800
rect 66074 0 66130 800
rect 66350 0 66406 800
rect 66534 0 66590 800
rect 66810 0 66866 800
rect 66994 0 67050 800
rect 67270 0 67326 800
rect 67454 0 67510 800
rect 67730 0 67786 800
rect 67914 0 67970 800
rect 68190 0 68246 800
rect 68374 0 68430 800
rect 68650 0 68706 800
rect 68834 0 68890 800
rect 69110 0 69166 800
rect 69294 0 69350 800
rect 69570 0 69626 800
rect 69754 0 69810 800
rect 70030 0 70086 800
rect 70214 0 70270 800
rect 70490 0 70546 800
rect 70674 0 70730 800
rect 70950 0 71006 800
rect 71134 0 71190 800
rect 71410 0 71466 800
rect 71594 0 71650 800
rect 71870 0 71926 800
rect 72054 0 72110 800
rect 72330 0 72386 800
rect 72514 0 72570 800
rect 72698 0 72754 800
rect 72974 0 73030 800
rect 73158 0 73214 800
rect 73434 0 73490 800
rect 73618 0 73674 800
rect 73894 0 73950 800
rect 74078 0 74134 800
rect 74354 0 74410 800
rect 74538 0 74594 800
rect 74814 0 74870 800
rect 74998 0 75054 800
rect 75274 0 75330 800
rect 75458 0 75514 800
rect 75734 0 75790 800
rect 75918 0 75974 800
rect 76194 0 76250 800
rect 76378 0 76434 800
rect 76654 0 76710 800
rect 76838 0 76894 800
rect 77114 0 77170 800
rect 77298 0 77354 800
rect 77574 0 77630 800
rect 77758 0 77814 800
rect 78034 0 78090 800
rect 78218 0 78274 800
rect 78494 0 78550 800
rect 78678 0 78734 800
rect 78954 0 79010 800
rect 79138 0 79194 800
rect 79414 0 79470 800
rect 79598 0 79654 800
rect 79782 0 79838 800
rect 80058 0 80114 800
rect 80242 0 80298 800
rect 80518 0 80574 800
rect 80702 0 80758 800
rect 80978 0 81034 800
rect 81162 0 81218 800
rect 81438 0 81494 800
rect 81622 0 81678 800
rect 81898 0 81954 800
rect 82082 0 82138 800
rect 82358 0 82414 800
rect 82542 0 82598 800
rect 82818 0 82874 800
rect 83002 0 83058 800
rect 83278 0 83334 800
rect 83462 0 83518 800
rect 83738 0 83794 800
rect 83922 0 83978 800
rect 84198 0 84254 800
rect 84382 0 84438 800
rect 84658 0 84714 800
rect 84842 0 84898 800
rect 85118 0 85174 800
rect 85302 0 85358 800
rect 85578 0 85634 800
rect 85762 0 85818 800
rect 86038 0 86094 800
rect 86222 0 86278 800
rect 86498 0 86554 800
rect 86682 0 86738 800
rect 86958 0 87014 800
rect 87142 0 87198 800
rect 87326 0 87382 800
rect 87602 0 87658 800
rect 87786 0 87842 800
rect 88062 0 88118 800
rect 88246 0 88302 800
rect 88522 0 88578 800
rect 88706 0 88762 800
rect 88982 0 89038 800
rect 89166 0 89222 800
rect 89442 0 89498 800
rect 89626 0 89682 800
rect 89902 0 89958 800
rect 90086 0 90142 800
rect 90362 0 90418 800
rect 90546 0 90602 800
rect 90822 0 90878 800
rect 91006 0 91062 800
rect 91282 0 91338 800
rect 91466 0 91522 800
rect 91742 0 91798 800
rect 91926 0 91982 800
rect 92202 0 92258 800
rect 92386 0 92442 800
rect 92662 0 92718 800
rect 92846 0 92902 800
rect 93122 0 93178 800
rect 93306 0 93362 800
rect 93582 0 93638 800
rect 93766 0 93822 800
rect 94042 0 94098 800
rect 94226 0 94282 800
rect 94410 0 94466 800
rect 94686 0 94742 800
rect 94870 0 94926 800
rect 95146 0 95202 800
rect 95330 0 95386 800
rect 95606 0 95662 800
rect 95790 0 95846 800
rect 96066 0 96122 800
rect 96250 0 96306 800
rect 96526 0 96582 800
rect 96710 0 96766 800
rect 96986 0 97042 800
rect 97170 0 97226 800
rect 97446 0 97502 800
rect 97630 0 97686 800
rect 97906 0 97962 800
rect 98090 0 98146 800
rect 98366 0 98422 800
rect 98550 0 98606 800
rect 98826 0 98882 800
rect 99010 0 99066 800
rect 99286 0 99342 800
rect 99470 0 99526 800
rect 99746 0 99802 800
rect 99930 0 99986 800
rect 100206 0 100262 800
rect 100390 0 100446 800
rect 100666 0 100722 800
rect 100850 0 100906 800
rect 101126 0 101182 800
rect 101310 0 101366 800
rect 101494 0 101550 800
rect 101770 0 101826 800
rect 101954 0 102010 800
rect 102230 0 102286 800
rect 102414 0 102470 800
rect 102690 0 102746 800
rect 102874 0 102930 800
rect 103150 0 103206 800
rect 103334 0 103390 800
rect 103610 0 103666 800
rect 103794 0 103850 800
rect 104070 0 104126 800
rect 104254 0 104310 800
rect 104530 0 104586 800
rect 104714 0 104770 800
rect 104990 0 105046 800
rect 105174 0 105230 800
rect 105450 0 105506 800
rect 105634 0 105690 800
rect 105910 0 105966 800
rect 106094 0 106150 800
rect 106370 0 106426 800
rect 106554 0 106610 800
rect 106830 0 106886 800
rect 107014 0 107070 800
rect 107290 0 107346 800
rect 107474 0 107530 800
rect 107750 0 107806 800
rect 107934 0 107990 800
rect 108210 0 108266 800
rect 108394 0 108450 800
rect 108670 0 108726 800
rect 108854 0 108910 800
rect 109038 0 109094 800
rect 109314 0 109370 800
rect 109498 0 109554 800
rect 109774 0 109830 800
rect 109958 0 110014 800
rect 110234 0 110290 800
rect 110418 0 110474 800
rect 110694 0 110750 800
rect 110878 0 110934 800
rect 111154 0 111210 800
rect 111338 0 111394 800
rect 111614 0 111670 800
rect 111798 0 111854 800
rect 112074 0 112130 800
rect 112258 0 112314 800
rect 112534 0 112590 800
rect 112718 0 112774 800
rect 112994 0 113050 800
rect 113178 0 113234 800
rect 113454 0 113510 800
rect 113638 0 113694 800
rect 113914 0 113970 800
rect 114098 0 114154 800
rect 114374 0 114430 800
rect 114558 0 114614 800
rect 114834 0 114890 800
rect 115018 0 115074 800
rect 115294 0 115350 800
rect 115478 0 115534 800
rect 115754 0 115810 800
rect 115938 0 115994 800
rect 116122 0 116178 800
rect 116398 0 116454 800
rect 116582 0 116638 800
rect 116858 0 116914 800
rect 117042 0 117098 800
rect 117318 0 117374 800
rect 117502 0 117558 800
rect 117778 0 117834 800
rect 117962 0 118018 800
rect 118238 0 118294 800
rect 118422 0 118478 800
rect 118698 0 118754 800
rect 118882 0 118938 800
rect 119158 0 119214 800
rect 119342 0 119398 800
rect 119618 0 119674 800
rect 119802 0 119858 800
rect 120078 0 120134 800
rect 120262 0 120318 800
rect 120538 0 120594 800
rect 120722 0 120778 800
rect 120998 0 121054 800
rect 121182 0 121238 800
rect 121458 0 121514 800
rect 121642 0 121698 800
rect 121918 0 121974 800
rect 122102 0 122158 800
rect 122378 0 122434 800
rect 122562 0 122618 800
rect 122838 0 122894 800
rect 123022 0 123078 800
rect 123206 0 123262 800
rect 123482 0 123538 800
rect 123666 0 123722 800
rect 123942 0 123998 800
rect 124126 0 124182 800
rect 124402 0 124458 800
rect 124586 0 124642 800
rect 124862 0 124918 800
rect 125046 0 125102 800
rect 125322 0 125378 800
rect 125506 0 125562 800
rect 125782 0 125838 800
rect 125966 0 126022 800
rect 126242 0 126298 800
rect 126426 0 126482 800
rect 126702 0 126758 800
rect 126886 0 126942 800
rect 127162 0 127218 800
rect 127346 0 127402 800
rect 127622 0 127678 800
rect 127806 0 127862 800
rect 128082 0 128138 800
rect 128266 0 128322 800
rect 128542 0 128598 800
rect 128726 0 128782 800
rect 129002 0 129058 800
rect 129186 0 129242 800
rect 129462 0 129518 800
rect 129646 0 129702 800
rect 129922 0 129978 800
rect 130106 0 130162 800
<< obsm2 >>
rect 20 131579 330 131730
rect 498 131579 1066 131730
rect 1234 131579 1802 131730
rect 1970 131579 2630 131730
rect 2798 131579 3366 131730
rect 3534 131579 4102 131730
rect 4270 131579 4930 131730
rect 5098 131579 5666 131730
rect 5834 131579 6494 131730
rect 6662 131579 7230 131730
rect 7398 131579 7966 131730
rect 8134 131579 8794 131730
rect 8962 131579 9530 131730
rect 9698 131579 10266 131730
rect 10434 131579 11094 131730
rect 11262 131579 11830 131730
rect 11998 131579 12658 131730
rect 12826 131579 13394 131730
rect 13562 131579 14130 131730
rect 14298 131579 14958 131730
rect 15126 131579 15694 131730
rect 15862 131579 16430 131730
rect 16598 131579 17258 131730
rect 17426 131579 17994 131730
rect 18162 131579 18822 131730
rect 18990 131579 19558 131730
rect 19726 131579 20294 131730
rect 20462 131579 21122 131730
rect 21290 131579 21858 131730
rect 22026 131579 22594 131730
rect 22762 131579 23422 131730
rect 23590 131579 24158 131730
rect 24326 131579 24986 131730
rect 25154 131579 25722 131730
rect 25890 131579 26458 131730
rect 26626 131579 27286 131730
rect 27454 131579 28022 131730
rect 28190 131579 28850 131730
rect 29018 131579 29586 131730
rect 29754 131579 30322 131730
rect 30490 131579 31150 131730
rect 31318 131579 31886 131730
rect 32054 131579 32622 131730
rect 32790 131579 33450 131730
rect 33618 131579 34186 131730
rect 34354 131579 35014 131730
rect 35182 131579 35750 131730
rect 35918 131579 36486 131730
rect 36654 131579 37314 131730
rect 37482 131579 38050 131730
rect 38218 131579 38786 131730
rect 38954 131579 39614 131730
rect 39782 131579 40350 131730
rect 40518 131579 41178 131730
rect 41346 131579 41914 131730
rect 42082 131579 42650 131730
rect 42818 131579 43478 131730
rect 43646 131579 44214 131730
rect 44382 131579 44950 131730
rect 45118 131579 45778 131730
rect 45946 131579 46514 131730
rect 46682 131579 47342 131730
rect 47510 131579 48078 131730
rect 48246 131579 48814 131730
rect 48982 131579 49642 131730
rect 49810 131579 50378 131730
rect 50546 131579 51114 131730
rect 51282 131579 51942 131730
rect 52110 131579 52678 131730
rect 52846 131579 53506 131730
rect 53674 131579 54242 131730
rect 54410 131579 54978 131730
rect 55146 131579 55806 131730
rect 55974 131579 56542 131730
rect 56710 131579 57370 131730
rect 57538 131579 58106 131730
rect 58274 131579 58842 131730
rect 59010 131579 59670 131730
rect 59838 131579 60406 131730
rect 60574 131579 61142 131730
rect 61310 131579 61970 131730
rect 62138 131579 62706 131730
rect 62874 131579 63534 131730
rect 63702 131579 64270 131730
rect 64438 131579 65006 131730
rect 65174 131579 65834 131730
rect 66002 131579 66570 131730
rect 66738 131579 67306 131730
rect 67474 131579 68134 131730
rect 68302 131579 68870 131730
rect 69038 131579 69698 131730
rect 69866 131579 70434 131730
rect 70602 131579 71170 131730
rect 71338 131579 71998 131730
rect 72166 131579 72734 131730
rect 72902 131579 73470 131730
rect 73638 131579 74298 131730
rect 74466 131579 75034 131730
rect 75202 131579 75862 131730
rect 76030 131579 76598 131730
rect 76766 131579 77334 131730
rect 77502 131579 78162 131730
rect 78330 131579 78898 131730
rect 79066 131579 79726 131730
rect 79894 131579 80462 131730
rect 80630 131579 81198 131730
rect 81366 131579 82026 131730
rect 82194 131579 82762 131730
rect 82930 131579 83498 131730
rect 83666 131579 84326 131730
rect 84494 131579 85062 131730
rect 85230 131579 85890 131730
rect 86058 131579 86626 131730
rect 86794 131579 87362 131730
rect 87530 131579 88190 131730
rect 88358 131579 88926 131730
rect 89094 131579 89662 131730
rect 89830 131579 90490 131730
rect 90658 131579 91226 131730
rect 91394 131579 92054 131730
rect 92222 131579 92790 131730
rect 92958 131579 93526 131730
rect 93694 131579 94354 131730
rect 94522 131579 95090 131730
rect 95258 131579 95826 131730
rect 95994 131579 96654 131730
rect 96822 131579 97390 131730
rect 97558 131579 98218 131730
rect 98386 131579 98954 131730
rect 99122 131579 99690 131730
rect 99858 131579 100518 131730
rect 100686 131579 101254 131730
rect 101422 131579 101990 131730
rect 102158 131579 102818 131730
rect 102986 131579 103554 131730
rect 103722 131579 104382 131730
rect 104550 131579 105118 131730
rect 105286 131579 105854 131730
rect 106022 131579 106682 131730
rect 106850 131579 107418 131730
rect 107586 131579 108246 131730
rect 108414 131579 108982 131730
rect 109150 131579 109718 131730
rect 109886 131579 110546 131730
rect 110714 131579 111282 131730
rect 111450 131579 112018 131730
rect 112186 131579 112846 131730
rect 113014 131579 113582 131730
rect 113750 131579 114410 131730
rect 114578 131579 115146 131730
rect 115314 131579 115882 131730
rect 116050 131579 116710 131730
rect 116878 131579 117446 131730
rect 117614 131579 118182 131730
rect 118350 131579 119010 131730
rect 119178 131579 119746 131730
rect 119914 131579 120574 131730
rect 120742 131579 121310 131730
rect 121478 131579 122046 131730
rect 122214 131579 122874 131730
rect 123042 131579 123610 131730
rect 123778 131579 124346 131730
rect 124514 131579 125174 131730
rect 125342 131579 125910 131730
rect 126078 131579 126738 131730
rect 126906 131579 127474 131730
rect 127642 131579 128210 131730
rect 128378 131579 129038 131730
rect 129206 131579 129774 131730
rect 129942 131579 130160 131730
rect 20 856 130160 131579
rect 20 303 54 856
rect 222 303 238 856
rect 406 303 422 856
rect 590 303 698 856
rect 866 303 882 856
rect 1050 303 1158 856
rect 1326 303 1342 856
rect 1510 303 1618 856
rect 1786 303 1802 856
rect 1970 303 2078 856
rect 2246 303 2262 856
rect 2430 303 2538 856
rect 2706 303 2722 856
rect 2890 303 2998 856
rect 3166 303 3182 856
rect 3350 303 3458 856
rect 3626 303 3642 856
rect 3810 303 3918 856
rect 4086 303 4102 856
rect 4270 303 4378 856
rect 4546 303 4562 856
rect 4730 303 4838 856
rect 5006 303 5022 856
rect 5190 303 5298 856
rect 5466 303 5482 856
rect 5650 303 5758 856
rect 5926 303 5942 856
rect 6110 303 6218 856
rect 6386 303 6402 856
rect 6570 303 6678 856
rect 6846 303 6862 856
rect 7030 303 7138 856
rect 7306 303 7322 856
rect 7490 303 7506 856
rect 7674 303 7782 856
rect 7950 303 7966 856
rect 8134 303 8242 856
rect 8410 303 8426 856
rect 8594 303 8702 856
rect 8870 303 8886 856
rect 9054 303 9162 856
rect 9330 303 9346 856
rect 9514 303 9622 856
rect 9790 303 9806 856
rect 9974 303 10082 856
rect 10250 303 10266 856
rect 10434 303 10542 856
rect 10710 303 10726 856
rect 10894 303 11002 856
rect 11170 303 11186 856
rect 11354 303 11462 856
rect 11630 303 11646 856
rect 11814 303 11922 856
rect 12090 303 12106 856
rect 12274 303 12382 856
rect 12550 303 12566 856
rect 12734 303 12842 856
rect 13010 303 13026 856
rect 13194 303 13302 856
rect 13470 303 13486 856
rect 13654 303 13762 856
rect 13930 303 13946 856
rect 14114 303 14222 856
rect 14390 303 14406 856
rect 14574 303 14590 856
rect 14758 303 14866 856
rect 15034 303 15050 856
rect 15218 303 15326 856
rect 15494 303 15510 856
rect 15678 303 15786 856
rect 15954 303 15970 856
rect 16138 303 16246 856
rect 16414 303 16430 856
rect 16598 303 16706 856
rect 16874 303 16890 856
rect 17058 303 17166 856
rect 17334 303 17350 856
rect 17518 303 17626 856
rect 17794 303 17810 856
rect 17978 303 18086 856
rect 18254 303 18270 856
rect 18438 303 18546 856
rect 18714 303 18730 856
rect 18898 303 19006 856
rect 19174 303 19190 856
rect 19358 303 19466 856
rect 19634 303 19650 856
rect 19818 303 19926 856
rect 20094 303 20110 856
rect 20278 303 20386 856
rect 20554 303 20570 856
rect 20738 303 20846 856
rect 21014 303 21030 856
rect 21198 303 21306 856
rect 21474 303 21490 856
rect 21658 303 21766 856
rect 21934 303 21950 856
rect 22118 303 22134 856
rect 22302 303 22410 856
rect 22578 303 22594 856
rect 22762 303 22870 856
rect 23038 303 23054 856
rect 23222 303 23330 856
rect 23498 303 23514 856
rect 23682 303 23790 856
rect 23958 303 23974 856
rect 24142 303 24250 856
rect 24418 303 24434 856
rect 24602 303 24710 856
rect 24878 303 24894 856
rect 25062 303 25170 856
rect 25338 303 25354 856
rect 25522 303 25630 856
rect 25798 303 25814 856
rect 25982 303 26090 856
rect 26258 303 26274 856
rect 26442 303 26550 856
rect 26718 303 26734 856
rect 26902 303 27010 856
rect 27178 303 27194 856
rect 27362 303 27470 856
rect 27638 303 27654 856
rect 27822 303 27930 856
rect 28098 303 28114 856
rect 28282 303 28390 856
rect 28558 303 28574 856
rect 28742 303 28850 856
rect 29018 303 29034 856
rect 29202 303 29218 856
rect 29386 303 29494 856
rect 29662 303 29678 856
rect 29846 303 29954 856
rect 30122 303 30138 856
rect 30306 303 30414 856
rect 30582 303 30598 856
rect 30766 303 30874 856
rect 31042 303 31058 856
rect 31226 303 31334 856
rect 31502 303 31518 856
rect 31686 303 31794 856
rect 31962 303 31978 856
rect 32146 303 32254 856
rect 32422 303 32438 856
rect 32606 303 32714 856
rect 32882 303 32898 856
rect 33066 303 33174 856
rect 33342 303 33358 856
rect 33526 303 33634 856
rect 33802 303 33818 856
rect 33986 303 34094 856
rect 34262 303 34278 856
rect 34446 303 34554 856
rect 34722 303 34738 856
rect 34906 303 35014 856
rect 35182 303 35198 856
rect 35366 303 35474 856
rect 35642 303 35658 856
rect 35826 303 35934 856
rect 36102 303 36118 856
rect 36286 303 36302 856
rect 36470 303 36578 856
rect 36746 303 36762 856
rect 36930 303 37038 856
rect 37206 303 37222 856
rect 37390 303 37498 856
rect 37666 303 37682 856
rect 37850 303 37958 856
rect 38126 303 38142 856
rect 38310 303 38418 856
rect 38586 303 38602 856
rect 38770 303 38878 856
rect 39046 303 39062 856
rect 39230 303 39338 856
rect 39506 303 39522 856
rect 39690 303 39798 856
rect 39966 303 39982 856
rect 40150 303 40258 856
rect 40426 303 40442 856
rect 40610 303 40718 856
rect 40886 303 40902 856
rect 41070 303 41178 856
rect 41346 303 41362 856
rect 41530 303 41638 856
rect 41806 303 41822 856
rect 41990 303 42098 856
rect 42266 303 42282 856
rect 42450 303 42558 856
rect 42726 303 42742 856
rect 42910 303 43018 856
rect 43186 303 43202 856
rect 43370 303 43478 856
rect 43646 303 43662 856
rect 43830 303 43846 856
rect 44014 303 44122 856
rect 44290 303 44306 856
rect 44474 303 44582 856
rect 44750 303 44766 856
rect 44934 303 45042 856
rect 45210 303 45226 856
rect 45394 303 45502 856
rect 45670 303 45686 856
rect 45854 303 45962 856
rect 46130 303 46146 856
rect 46314 303 46422 856
rect 46590 303 46606 856
rect 46774 303 46882 856
rect 47050 303 47066 856
rect 47234 303 47342 856
rect 47510 303 47526 856
rect 47694 303 47802 856
rect 47970 303 47986 856
rect 48154 303 48262 856
rect 48430 303 48446 856
rect 48614 303 48722 856
rect 48890 303 48906 856
rect 49074 303 49182 856
rect 49350 303 49366 856
rect 49534 303 49642 856
rect 49810 303 49826 856
rect 49994 303 50102 856
rect 50270 303 50286 856
rect 50454 303 50562 856
rect 50730 303 50746 856
rect 50914 303 50930 856
rect 51098 303 51206 856
rect 51374 303 51390 856
rect 51558 303 51666 856
rect 51834 303 51850 856
rect 52018 303 52126 856
rect 52294 303 52310 856
rect 52478 303 52586 856
rect 52754 303 52770 856
rect 52938 303 53046 856
rect 53214 303 53230 856
rect 53398 303 53506 856
rect 53674 303 53690 856
rect 53858 303 53966 856
rect 54134 303 54150 856
rect 54318 303 54426 856
rect 54594 303 54610 856
rect 54778 303 54886 856
rect 55054 303 55070 856
rect 55238 303 55346 856
rect 55514 303 55530 856
rect 55698 303 55806 856
rect 55974 303 55990 856
rect 56158 303 56266 856
rect 56434 303 56450 856
rect 56618 303 56726 856
rect 56894 303 56910 856
rect 57078 303 57186 856
rect 57354 303 57370 856
rect 57538 303 57646 856
rect 57814 303 57830 856
rect 57998 303 58014 856
rect 58182 303 58290 856
rect 58458 303 58474 856
rect 58642 303 58750 856
rect 58918 303 58934 856
rect 59102 303 59210 856
rect 59378 303 59394 856
rect 59562 303 59670 856
rect 59838 303 59854 856
rect 60022 303 60130 856
rect 60298 303 60314 856
rect 60482 303 60590 856
rect 60758 303 60774 856
rect 60942 303 61050 856
rect 61218 303 61234 856
rect 61402 303 61510 856
rect 61678 303 61694 856
rect 61862 303 61970 856
rect 62138 303 62154 856
rect 62322 303 62430 856
rect 62598 303 62614 856
rect 62782 303 62890 856
rect 63058 303 63074 856
rect 63242 303 63350 856
rect 63518 303 63534 856
rect 63702 303 63810 856
rect 63978 303 63994 856
rect 64162 303 64270 856
rect 64438 303 64454 856
rect 64622 303 64730 856
rect 64898 303 64914 856
rect 65082 303 65190 856
rect 65358 303 65374 856
rect 65542 303 65558 856
rect 65726 303 65834 856
rect 66002 303 66018 856
rect 66186 303 66294 856
rect 66462 303 66478 856
rect 66646 303 66754 856
rect 66922 303 66938 856
rect 67106 303 67214 856
rect 67382 303 67398 856
rect 67566 303 67674 856
rect 67842 303 67858 856
rect 68026 303 68134 856
rect 68302 303 68318 856
rect 68486 303 68594 856
rect 68762 303 68778 856
rect 68946 303 69054 856
rect 69222 303 69238 856
rect 69406 303 69514 856
rect 69682 303 69698 856
rect 69866 303 69974 856
rect 70142 303 70158 856
rect 70326 303 70434 856
rect 70602 303 70618 856
rect 70786 303 70894 856
rect 71062 303 71078 856
rect 71246 303 71354 856
rect 71522 303 71538 856
rect 71706 303 71814 856
rect 71982 303 71998 856
rect 72166 303 72274 856
rect 72442 303 72458 856
rect 72626 303 72642 856
rect 72810 303 72918 856
rect 73086 303 73102 856
rect 73270 303 73378 856
rect 73546 303 73562 856
rect 73730 303 73838 856
rect 74006 303 74022 856
rect 74190 303 74298 856
rect 74466 303 74482 856
rect 74650 303 74758 856
rect 74926 303 74942 856
rect 75110 303 75218 856
rect 75386 303 75402 856
rect 75570 303 75678 856
rect 75846 303 75862 856
rect 76030 303 76138 856
rect 76306 303 76322 856
rect 76490 303 76598 856
rect 76766 303 76782 856
rect 76950 303 77058 856
rect 77226 303 77242 856
rect 77410 303 77518 856
rect 77686 303 77702 856
rect 77870 303 77978 856
rect 78146 303 78162 856
rect 78330 303 78438 856
rect 78606 303 78622 856
rect 78790 303 78898 856
rect 79066 303 79082 856
rect 79250 303 79358 856
rect 79526 303 79542 856
rect 79710 303 79726 856
rect 79894 303 80002 856
rect 80170 303 80186 856
rect 80354 303 80462 856
rect 80630 303 80646 856
rect 80814 303 80922 856
rect 81090 303 81106 856
rect 81274 303 81382 856
rect 81550 303 81566 856
rect 81734 303 81842 856
rect 82010 303 82026 856
rect 82194 303 82302 856
rect 82470 303 82486 856
rect 82654 303 82762 856
rect 82930 303 82946 856
rect 83114 303 83222 856
rect 83390 303 83406 856
rect 83574 303 83682 856
rect 83850 303 83866 856
rect 84034 303 84142 856
rect 84310 303 84326 856
rect 84494 303 84602 856
rect 84770 303 84786 856
rect 84954 303 85062 856
rect 85230 303 85246 856
rect 85414 303 85522 856
rect 85690 303 85706 856
rect 85874 303 85982 856
rect 86150 303 86166 856
rect 86334 303 86442 856
rect 86610 303 86626 856
rect 86794 303 86902 856
rect 87070 303 87086 856
rect 87254 303 87270 856
rect 87438 303 87546 856
rect 87714 303 87730 856
rect 87898 303 88006 856
rect 88174 303 88190 856
rect 88358 303 88466 856
rect 88634 303 88650 856
rect 88818 303 88926 856
rect 89094 303 89110 856
rect 89278 303 89386 856
rect 89554 303 89570 856
rect 89738 303 89846 856
rect 90014 303 90030 856
rect 90198 303 90306 856
rect 90474 303 90490 856
rect 90658 303 90766 856
rect 90934 303 90950 856
rect 91118 303 91226 856
rect 91394 303 91410 856
rect 91578 303 91686 856
rect 91854 303 91870 856
rect 92038 303 92146 856
rect 92314 303 92330 856
rect 92498 303 92606 856
rect 92774 303 92790 856
rect 92958 303 93066 856
rect 93234 303 93250 856
rect 93418 303 93526 856
rect 93694 303 93710 856
rect 93878 303 93986 856
rect 94154 303 94170 856
rect 94338 303 94354 856
rect 94522 303 94630 856
rect 94798 303 94814 856
rect 94982 303 95090 856
rect 95258 303 95274 856
rect 95442 303 95550 856
rect 95718 303 95734 856
rect 95902 303 96010 856
rect 96178 303 96194 856
rect 96362 303 96470 856
rect 96638 303 96654 856
rect 96822 303 96930 856
rect 97098 303 97114 856
rect 97282 303 97390 856
rect 97558 303 97574 856
rect 97742 303 97850 856
rect 98018 303 98034 856
rect 98202 303 98310 856
rect 98478 303 98494 856
rect 98662 303 98770 856
rect 98938 303 98954 856
rect 99122 303 99230 856
rect 99398 303 99414 856
rect 99582 303 99690 856
rect 99858 303 99874 856
rect 100042 303 100150 856
rect 100318 303 100334 856
rect 100502 303 100610 856
rect 100778 303 100794 856
rect 100962 303 101070 856
rect 101238 303 101254 856
rect 101422 303 101438 856
rect 101606 303 101714 856
rect 101882 303 101898 856
rect 102066 303 102174 856
rect 102342 303 102358 856
rect 102526 303 102634 856
rect 102802 303 102818 856
rect 102986 303 103094 856
rect 103262 303 103278 856
rect 103446 303 103554 856
rect 103722 303 103738 856
rect 103906 303 104014 856
rect 104182 303 104198 856
rect 104366 303 104474 856
rect 104642 303 104658 856
rect 104826 303 104934 856
rect 105102 303 105118 856
rect 105286 303 105394 856
rect 105562 303 105578 856
rect 105746 303 105854 856
rect 106022 303 106038 856
rect 106206 303 106314 856
rect 106482 303 106498 856
rect 106666 303 106774 856
rect 106942 303 106958 856
rect 107126 303 107234 856
rect 107402 303 107418 856
rect 107586 303 107694 856
rect 107862 303 107878 856
rect 108046 303 108154 856
rect 108322 303 108338 856
rect 108506 303 108614 856
rect 108782 303 108798 856
rect 108966 303 108982 856
rect 109150 303 109258 856
rect 109426 303 109442 856
rect 109610 303 109718 856
rect 109886 303 109902 856
rect 110070 303 110178 856
rect 110346 303 110362 856
rect 110530 303 110638 856
rect 110806 303 110822 856
rect 110990 303 111098 856
rect 111266 303 111282 856
rect 111450 303 111558 856
rect 111726 303 111742 856
rect 111910 303 112018 856
rect 112186 303 112202 856
rect 112370 303 112478 856
rect 112646 303 112662 856
rect 112830 303 112938 856
rect 113106 303 113122 856
rect 113290 303 113398 856
rect 113566 303 113582 856
rect 113750 303 113858 856
rect 114026 303 114042 856
rect 114210 303 114318 856
rect 114486 303 114502 856
rect 114670 303 114778 856
rect 114946 303 114962 856
rect 115130 303 115238 856
rect 115406 303 115422 856
rect 115590 303 115698 856
rect 115866 303 115882 856
rect 116050 303 116066 856
rect 116234 303 116342 856
rect 116510 303 116526 856
rect 116694 303 116802 856
rect 116970 303 116986 856
rect 117154 303 117262 856
rect 117430 303 117446 856
rect 117614 303 117722 856
rect 117890 303 117906 856
rect 118074 303 118182 856
rect 118350 303 118366 856
rect 118534 303 118642 856
rect 118810 303 118826 856
rect 118994 303 119102 856
rect 119270 303 119286 856
rect 119454 303 119562 856
rect 119730 303 119746 856
rect 119914 303 120022 856
rect 120190 303 120206 856
rect 120374 303 120482 856
rect 120650 303 120666 856
rect 120834 303 120942 856
rect 121110 303 121126 856
rect 121294 303 121402 856
rect 121570 303 121586 856
rect 121754 303 121862 856
rect 122030 303 122046 856
rect 122214 303 122322 856
rect 122490 303 122506 856
rect 122674 303 122782 856
rect 122950 303 122966 856
rect 123134 303 123150 856
rect 123318 303 123426 856
rect 123594 303 123610 856
rect 123778 303 123886 856
rect 124054 303 124070 856
rect 124238 303 124346 856
rect 124514 303 124530 856
rect 124698 303 124806 856
rect 124974 303 124990 856
rect 125158 303 125266 856
rect 125434 303 125450 856
rect 125618 303 125726 856
rect 125894 303 125910 856
rect 126078 303 126186 856
rect 126354 303 126370 856
rect 126538 303 126646 856
rect 126814 303 126830 856
rect 126998 303 127106 856
rect 127274 303 127290 856
rect 127458 303 127566 856
rect 127734 303 127750 856
rect 127918 303 128026 856
rect 128194 303 128210 856
rect 128378 303 128486 856
rect 128654 303 128670 856
rect 128838 303 128946 856
rect 129114 303 129130 856
rect 129298 303 129406 856
rect 129574 303 129590 856
rect 129758 303 129866 856
rect 130034 303 130050 856
<< obsm3 >>
rect 1025 307 128603 130049
<< metal4 >>
rect 4208 2128 4528 130064
rect 19568 2128 19888 130064
rect 34928 2128 35248 130064
rect 50288 2128 50608 130064
rect 65648 2128 65968 130064
rect 81008 2128 81328 130064
rect 96368 2128 96688 130064
rect 111728 2128 112048 130064
rect 127088 2128 127408 130064
<< obsm4 >>
rect 1163 2048 4128 129981
rect 4608 2048 19488 129981
rect 19968 2048 34848 129981
rect 35328 2048 50208 129981
rect 50688 2048 65568 129981
rect 66048 2048 80928 129981
rect 81408 2048 96288 129981
rect 96768 2048 111648 129981
rect 112128 2048 127008 129981
rect 127488 2048 127821 129981
rect 1163 307 127821 2048
<< labels >>
rlabel metal2 s 2686 131635 2742 132435 6 dram_addr0[0]
port 1 nsew signal output
rlabel metal2 s 5722 131635 5778 132435 6 dram_addr0[1]
port 2 nsew signal output
rlabel metal2 s 8850 131635 8906 132435 6 dram_addr0[2]
port 3 nsew signal output
rlabel metal2 s 11886 131635 11942 132435 6 dram_addr0[3]
port 4 nsew signal output
rlabel metal2 s 15014 131635 15070 132435 6 dram_addr0[4]
port 5 nsew signal output
rlabel metal2 s 17314 131635 17370 132435 6 dram_addr0[5]
port 6 nsew signal output
rlabel metal2 s 19614 131635 19670 132435 6 dram_addr0[6]
port 7 nsew signal output
rlabel metal2 s 21914 131635 21970 132435 6 dram_addr0[7]
port 8 nsew signal output
rlabel metal2 s 24214 131635 24270 132435 6 dram_addr0[8]
port 9 nsew signal output
rlabel metal2 s 386 131635 442 132435 6 dram_clk0
port 10 nsew signal output
rlabel metal2 s 1122 131635 1178 132435 6 dram_csb0
port 11 nsew signal output
rlabel metal2 s 3422 131635 3478 132435 6 dram_din0[0]
port 12 nsew signal output
rlabel metal2 s 28078 131635 28134 132435 6 dram_din0[10]
port 13 nsew signal output
rlabel metal2 s 29642 131635 29698 132435 6 dram_din0[11]
port 14 nsew signal output
rlabel metal2 s 31206 131635 31262 132435 6 dram_din0[12]
port 15 nsew signal output
rlabel metal2 s 32678 131635 32734 132435 6 dram_din0[13]
port 16 nsew signal output
rlabel metal2 s 34242 131635 34298 132435 6 dram_din0[14]
port 17 nsew signal output
rlabel metal2 s 35806 131635 35862 132435 6 dram_din0[15]
port 18 nsew signal output
rlabel metal2 s 37370 131635 37426 132435 6 dram_din0[16]
port 19 nsew signal output
rlabel metal2 s 38842 131635 38898 132435 6 dram_din0[17]
port 20 nsew signal output
rlabel metal2 s 40406 131635 40462 132435 6 dram_din0[18]
port 21 nsew signal output
rlabel metal2 s 41970 131635 42026 132435 6 dram_din0[19]
port 22 nsew signal output
rlabel metal2 s 6550 131635 6606 132435 6 dram_din0[1]
port 23 nsew signal output
rlabel metal2 s 43534 131635 43590 132435 6 dram_din0[20]
port 24 nsew signal output
rlabel metal2 s 45006 131635 45062 132435 6 dram_din0[21]
port 25 nsew signal output
rlabel metal2 s 46570 131635 46626 132435 6 dram_din0[22]
port 26 nsew signal output
rlabel metal2 s 48134 131635 48190 132435 6 dram_din0[23]
port 27 nsew signal output
rlabel metal2 s 49698 131635 49754 132435 6 dram_din0[24]
port 28 nsew signal output
rlabel metal2 s 51170 131635 51226 132435 6 dram_din0[25]
port 29 nsew signal output
rlabel metal2 s 52734 131635 52790 132435 6 dram_din0[26]
port 30 nsew signal output
rlabel metal2 s 54298 131635 54354 132435 6 dram_din0[27]
port 31 nsew signal output
rlabel metal2 s 55862 131635 55918 132435 6 dram_din0[28]
port 32 nsew signal output
rlabel metal2 s 57426 131635 57482 132435 6 dram_din0[29]
port 33 nsew signal output
rlabel metal2 s 9586 131635 9642 132435 6 dram_din0[2]
port 34 nsew signal output
rlabel metal2 s 58898 131635 58954 132435 6 dram_din0[30]
port 35 nsew signal output
rlabel metal2 s 60462 131635 60518 132435 6 dram_din0[31]
port 36 nsew signal output
rlabel metal2 s 12714 131635 12770 132435 6 dram_din0[3]
port 37 nsew signal output
rlabel metal2 s 15750 131635 15806 132435 6 dram_din0[4]
port 38 nsew signal output
rlabel metal2 s 18050 131635 18106 132435 6 dram_din0[5]
port 39 nsew signal output
rlabel metal2 s 20350 131635 20406 132435 6 dram_din0[6]
port 40 nsew signal output
rlabel metal2 s 22650 131635 22706 132435 6 dram_din0[7]
port 41 nsew signal output
rlabel metal2 s 25042 131635 25098 132435 6 dram_din0[8]
port 42 nsew signal output
rlabel metal2 s 26514 131635 26570 132435 6 dram_din0[9]
port 43 nsew signal output
rlabel metal2 s 4158 131635 4214 132435 6 dram_dout0[0]
port 44 nsew signal input
rlabel metal2 s 28906 131635 28962 132435 6 dram_dout0[10]
port 45 nsew signal input
rlabel metal2 s 30378 131635 30434 132435 6 dram_dout0[11]
port 46 nsew signal input
rlabel metal2 s 31942 131635 31998 132435 6 dram_dout0[12]
port 47 nsew signal input
rlabel metal2 s 33506 131635 33562 132435 6 dram_dout0[13]
port 48 nsew signal input
rlabel metal2 s 35070 131635 35126 132435 6 dram_dout0[14]
port 49 nsew signal input
rlabel metal2 s 36542 131635 36598 132435 6 dram_dout0[15]
port 50 nsew signal input
rlabel metal2 s 38106 131635 38162 132435 6 dram_dout0[16]
port 51 nsew signal input
rlabel metal2 s 39670 131635 39726 132435 6 dram_dout0[17]
port 52 nsew signal input
rlabel metal2 s 41234 131635 41290 132435 6 dram_dout0[18]
port 53 nsew signal input
rlabel metal2 s 42706 131635 42762 132435 6 dram_dout0[19]
port 54 nsew signal input
rlabel metal2 s 7286 131635 7342 132435 6 dram_dout0[1]
port 55 nsew signal input
rlabel metal2 s 44270 131635 44326 132435 6 dram_dout0[20]
port 56 nsew signal input
rlabel metal2 s 45834 131635 45890 132435 6 dram_dout0[21]
port 57 nsew signal input
rlabel metal2 s 47398 131635 47454 132435 6 dram_dout0[22]
port 58 nsew signal input
rlabel metal2 s 48870 131635 48926 132435 6 dram_dout0[23]
port 59 nsew signal input
rlabel metal2 s 50434 131635 50490 132435 6 dram_dout0[24]
port 60 nsew signal input
rlabel metal2 s 51998 131635 52054 132435 6 dram_dout0[25]
port 61 nsew signal input
rlabel metal2 s 53562 131635 53618 132435 6 dram_dout0[26]
port 62 nsew signal input
rlabel metal2 s 55034 131635 55090 132435 6 dram_dout0[27]
port 63 nsew signal input
rlabel metal2 s 56598 131635 56654 132435 6 dram_dout0[28]
port 64 nsew signal input
rlabel metal2 s 58162 131635 58218 132435 6 dram_dout0[29]
port 65 nsew signal input
rlabel metal2 s 10322 131635 10378 132435 6 dram_dout0[2]
port 66 nsew signal input
rlabel metal2 s 59726 131635 59782 132435 6 dram_dout0[30]
port 67 nsew signal input
rlabel metal2 s 61198 131635 61254 132435 6 dram_dout0[31]
port 68 nsew signal input
rlabel metal2 s 13450 131635 13506 132435 6 dram_dout0[3]
port 69 nsew signal input
rlabel metal2 s 16486 131635 16542 132435 6 dram_dout0[4]
port 70 nsew signal input
rlabel metal2 s 18878 131635 18934 132435 6 dram_dout0[5]
port 71 nsew signal input
rlabel metal2 s 21178 131635 21234 132435 6 dram_dout0[6]
port 72 nsew signal input
rlabel metal2 s 23478 131635 23534 132435 6 dram_dout0[7]
port 73 nsew signal input
rlabel metal2 s 25778 131635 25834 132435 6 dram_dout0[8]
port 74 nsew signal input
rlabel metal2 s 27342 131635 27398 132435 6 dram_dout0[9]
port 75 nsew signal input
rlabel metal2 s 1858 131635 1914 132435 6 dram_web0
port 76 nsew signal output
rlabel metal2 s 4986 131635 5042 132435 6 dram_wmask0[0]
port 77 nsew signal output
rlabel metal2 s 8022 131635 8078 132435 6 dram_wmask0[1]
port 78 nsew signal output
rlabel metal2 s 11150 131635 11206 132435 6 dram_wmask0[2]
port 79 nsew signal output
rlabel metal2 s 14186 131635 14242 132435 6 dram_wmask0[3]
port 80 nsew signal output
rlabel metal2 s 64326 131635 64382 132435 6 gpio_in[0]
port 81 nsew signal input
rlabel metal2 s 87418 131635 87474 132435 6 gpio_in[10]
port 82 nsew signal input
rlabel metal2 s 89718 131635 89774 132435 6 gpio_in[11]
port 83 nsew signal input
rlabel metal2 s 92110 131635 92166 132435 6 gpio_in[12]
port 84 nsew signal input
rlabel metal2 s 94410 131635 94466 132435 6 gpio_in[13]
port 85 nsew signal input
rlabel metal2 s 96710 131635 96766 132435 6 gpio_in[14]
port 86 nsew signal input
rlabel metal2 s 99010 131635 99066 132435 6 gpio_in[15]
port 87 nsew signal input
rlabel metal2 s 101310 131635 101366 132435 6 gpio_in[16]
port 88 nsew signal input
rlabel metal2 s 103610 131635 103666 132435 6 gpio_in[17]
port 89 nsew signal input
rlabel metal2 s 105910 131635 105966 132435 6 gpio_in[18]
port 90 nsew signal input
rlabel metal2 s 108302 131635 108358 132435 6 gpio_in[19]
port 91 nsew signal input
rlabel metal2 s 66626 131635 66682 132435 6 gpio_in[1]
port 92 nsew signal input
rlabel metal2 s 110602 131635 110658 132435 6 gpio_in[20]
port 93 nsew signal input
rlabel metal2 s 112902 131635 112958 132435 6 gpio_in[21]
port 94 nsew signal input
rlabel metal2 s 115202 131635 115258 132435 6 gpio_in[22]
port 95 nsew signal input
rlabel metal2 s 117502 131635 117558 132435 6 gpio_in[23]
port 96 nsew signal input
rlabel metal2 s 68926 131635 68982 132435 6 gpio_in[2]
port 97 nsew signal input
rlabel metal2 s 71226 131635 71282 132435 6 gpio_in[3]
port 98 nsew signal input
rlabel metal2 s 73526 131635 73582 132435 6 gpio_in[4]
port 99 nsew signal input
rlabel metal2 s 75918 131635 75974 132435 6 gpio_in[5]
port 100 nsew signal input
rlabel metal2 s 78218 131635 78274 132435 6 gpio_in[6]
port 101 nsew signal input
rlabel metal2 s 80518 131635 80574 132435 6 gpio_in[7]
port 102 nsew signal input
rlabel metal2 s 82818 131635 82874 132435 6 gpio_in[8]
port 103 nsew signal input
rlabel metal2 s 85118 131635 85174 132435 6 gpio_in[9]
port 104 nsew signal input
rlabel metal2 s 65062 131635 65118 132435 6 gpio_oeb[0]
port 105 nsew signal output
rlabel metal2 s 88246 131635 88302 132435 6 gpio_oeb[10]
port 106 nsew signal output
rlabel metal2 s 90546 131635 90602 132435 6 gpio_oeb[11]
port 107 nsew signal output
rlabel metal2 s 92846 131635 92902 132435 6 gpio_oeb[12]
port 108 nsew signal output
rlabel metal2 s 95146 131635 95202 132435 6 gpio_oeb[13]
port 109 nsew signal output
rlabel metal2 s 97446 131635 97502 132435 6 gpio_oeb[14]
port 110 nsew signal output
rlabel metal2 s 99746 131635 99802 132435 6 gpio_oeb[15]
port 111 nsew signal output
rlabel metal2 s 102046 131635 102102 132435 6 gpio_oeb[16]
port 112 nsew signal output
rlabel metal2 s 104438 131635 104494 132435 6 gpio_oeb[17]
port 113 nsew signal output
rlabel metal2 s 106738 131635 106794 132435 6 gpio_oeb[18]
port 114 nsew signal output
rlabel metal2 s 109038 131635 109094 132435 6 gpio_oeb[19]
port 115 nsew signal output
rlabel metal2 s 67362 131635 67418 132435 6 gpio_oeb[1]
port 116 nsew signal output
rlabel metal2 s 111338 131635 111394 132435 6 gpio_oeb[20]
port 117 nsew signal output
rlabel metal2 s 113638 131635 113694 132435 6 gpio_oeb[21]
port 118 nsew signal output
rlabel metal2 s 115938 131635 115994 132435 6 gpio_oeb[22]
port 119 nsew signal output
rlabel metal2 s 118238 131635 118294 132435 6 gpio_oeb[23]
port 120 nsew signal output
rlabel metal2 s 119802 131635 119858 132435 6 gpio_oeb[24]
port 121 nsew signal output
rlabel metal2 s 120630 131635 120686 132435 6 gpio_oeb[25]
port 122 nsew signal output
rlabel metal2 s 121366 131635 121422 132435 6 gpio_oeb[26]
port 123 nsew signal output
rlabel metal2 s 122102 131635 122158 132435 6 gpio_oeb[27]
port 124 nsew signal output
rlabel metal2 s 122930 131635 122986 132435 6 gpio_oeb[28]
port 125 nsew signal output
rlabel metal2 s 123666 131635 123722 132435 6 gpio_oeb[29]
port 126 nsew signal output
rlabel metal2 s 69754 131635 69810 132435 6 gpio_oeb[2]
port 127 nsew signal output
rlabel metal2 s 124402 131635 124458 132435 6 gpio_oeb[30]
port 128 nsew signal output
rlabel metal2 s 125230 131635 125286 132435 6 gpio_oeb[31]
port 129 nsew signal output
rlabel metal2 s 125966 131635 126022 132435 6 gpio_oeb[32]
port 130 nsew signal output
rlabel metal2 s 126794 131635 126850 132435 6 gpio_oeb[33]
port 131 nsew signal output
rlabel metal2 s 127530 131635 127586 132435 6 gpio_oeb[34]
port 132 nsew signal output
rlabel metal2 s 128266 131635 128322 132435 6 gpio_oeb[35]
port 133 nsew signal output
rlabel metal2 s 129094 131635 129150 132435 6 gpio_oeb[36]
port 134 nsew signal output
rlabel metal2 s 129830 131635 129886 132435 6 gpio_oeb[37]
port 135 nsew signal output
rlabel metal2 s 72054 131635 72110 132435 6 gpio_oeb[3]
port 136 nsew signal output
rlabel metal2 s 74354 131635 74410 132435 6 gpio_oeb[4]
port 137 nsew signal output
rlabel metal2 s 76654 131635 76710 132435 6 gpio_oeb[5]
port 138 nsew signal output
rlabel metal2 s 78954 131635 79010 132435 6 gpio_oeb[6]
port 139 nsew signal output
rlabel metal2 s 81254 131635 81310 132435 6 gpio_oeb[7]
port 140 nsew signal output
rlabel metal2 s 83554 131635 83610 132435 6 gpio_oeb[8]
port 141 nsew signal output
rlabel metal2 s 85946 131635 86002 132435 6 gpio_oeb[9]
port 142 nsew signal output
rlabel metal2 s 65890 131635 65946 132435 6 gpio_out[0]
port 143 nsew signal output
rlabel metal2 s 88982 131635 89038 132435 6 gpio_out[10]
port 144 nsew signal output
rlabel metal2 s 91282 131635 91338 132435 6 gpio_out[11]
port 145 nsew signal output
rlabel metal2 s 93582 131635 93638 132435 6 gpio_out[12]
port 146 nsew signal output
rlabel metal2 s 95882 131635 95938 132435 6 gpio_out[13]
port 147 nsew signal output
rlabel metal2 s 98274 131635 98330 132435 6 gpio_out[14]
port 148 nsew signal output
rlabel metal2 s 100574 131635 100630 132435 6 gpio_out[15]
port 149 nsew signal output
rlabel metal2 s 102874 131635 102930 132435 6 gpio_out[16]
port 150 nsew signal output
rlabel metal2 s 105174 131635 105230 132435 6 gpio_out[17]
port 151 nsew signal output
rlabel metal2 s 107474 131635 107530 132435 6 gpio_out[18]
port 152 nsew signal output
rlabel metal2 s 109774 131635 109830 132435 6 gpio_out[19]
port 153 nsew signal output
rlabel metal2 s 68190 131635 68246 132435 6 gpio_out[1]
port 154 nsew signal output
rlabel metal2 s 112074 131635 112130 132435 6 gpio_out[20]
port 155 nsew signal output
rlabel metal2 s 114466 131635 114522 132435 6 gpio_out[21]
port 156 nsew signal output
rlabel metal2 s 116766 131635 116822 132435 6 gpio_out[22]
port 157 nsew signal output
rlabel metal2 s 119066 131635 119122 132435 6 gpio_out[23]
port 158 nsew signal output
rlabel metal2 s 70490 131635 70546 132435 6 gpio_out[2]
port 159 nsew signal output
rlabel metal2 s 72790 131635 72846 132435 6 gpio_out[3]
port 160 nsew signal output
rlabel metal2 s 75090 131635 75146 132435 6 gpio_out[4]
port 161 nsew signal output
rlabel metal2 s 77390 131635 77446 132435 6 gpio_out[5]
port 162 nsew signal output
rlabel metal2 s 79782 131635 79838 132435 6 gpio_out[6]
port 163 nsew signal output
rlabel metal2 s 82082 131635 82138 132435 6 gpio_out[7]
port 164 nsew signal output
rlabel metal2 s 84382 131635 84438 132435 6 gpio_out[8]
port 165 nsew signal output
rlabel metal2 s 86682 131635 86738 132435 6 gpio_out[9]
port 166 nsew signal output
rlabel metal2 s 112718 0 112774 800 6 iram_addr0[0]
port 167 nsew signal output
rlabel metal2 s 113638 0 113694 800 6 iram_addr0[1]
port 168 nsew signal output
rlabel metal2 s 114558 0 114614 800 6 iram_addr0[2]
port 169 nsew signal output
rlabel metal2 s 115478 0 115534 800 6 iram_addr0[3]
port 170 nsew signal output
rlabel metal2 s 116398 0 116454 800 6 iram_addr0[4]
port 171 nsew signal output
rlabel metal2 s 117042 0 117098 800 6 iram_addr0[5]
port 172 nsew signal output
rlabel metal2 s 117778 0 117834 800 6 iram_addr0[6]
port 173 nsew signal output
rlabel metal2 s 118422 0 118478 800 6 iram_addr0[7]
port 174 nsew signal output
rlabel metal2 s 119158 0 119214 800 6 iram_addr0[8]
port 175 nsew signal output
rlabel metal2 s 112074 0 112130 800 6 iram_clk0
port 176 nsew signal output
rlabel metal2 s 112258 0 112314 800 6 iram_csb0
port 177 nsew signal output
rlabel metal2 s 112994 0 113050 800 6 iram_din0[0]
port 178 nsew signal output
rlabel metal2 s 120262 0 120318 800 6 iram_din0[10]
port 179 nsew signal output
rlabel metal2 s 120722 0 120778 800 6 iram_din0[11]
port 180 nsew signal output
rlabel metal2 s 121182 0 121238 800 6 iram_din0[12]
port 181 nsew signal output
rlabel metal2 s 121642 0 121698 800 6 iram_din0[13]
port 182 nsew signal output
rlabel metal2 s 122102 0 122158 800 6 iram_din0[14]
port 183 nsew signal output
rlabel metal2 s 122562 0 122618 800 6 iram_din0[15]
port 184 nsew signal output
rlabel metal2 s 123022 0 123078 800 6 iram_din0[16]
port 185 nsew signal output
rlabel metal2 s 123482 0 123538 800 6 iram_din0[17]
port 186 nsew signal output
rlabel metal2 s 123942 0 123998 800 6 iram_din0[18]
port 187 nsew signal output
rlabel metal2 s 124402 0 124458 800 6 iram_din0[19]
port 188 nsew signal output
rlabel metal2 s 113914 0 113970 800 6 iram_din0[1]
port 189 nsew signal output
rlabel metal2 s 124862 0 124918 800 6 iram_din0[20]
port 190 nsew signal output
rlabel metal2 s 125322 0 125378 800 6 iram_din0[21]
port 191 nsew signal output
rlabel metal2 s 125782 0 125838 800 6 iram_din0[22]
port 192 nsew signal output
rlabel metal2 s 126242 0 126298 800 6 iram_din0[23]
port 193 nsew signal output
rlabel metal2 s 126702 0 126758 800 6 iram_din0[24]
port 194 nsew signal output
rlabel metal2 s 127162 0 127218 800 6 iram_din0[25]
port 195 nsew signal output
rlabel metal2 s 127622 0 127678 800 6 iram_din0[26]
port 196 nsew signal output
rlabel metal2 s 128082 0 128138 800 6 iram_din0[27]
port 197 nsew signal output
rlabel metal2 s 128542 0 128598 800 6 iram_din0[28]
port 198 nsew signal output
rlabel metal2 s 129002 0 129058 800 6 iram_din0[29]
port 199 nsew signal output
rlabel metal2 s 114834 0 114890 800 6 iram_din0[2]
port 200 nsew signal output
rlabel metal2 s 129462 0 129518 800 6 iram_din0[30]
port 201 nsew signal output
rlabel metal2 s 129922 0 129978 800 6 iram_din0[31]
port 202 nsew signal output
rlabel metal2 s 115754 0 115810 800 6 iram_din0[3]
port 203 nsew signal output
rlabel metal2 s 116582 0 116638 800 6 iram_din0[4]
port 204 nsew signal output
rlabel metal2 s 117318 0 117374 800 6 iram_din0[5]
port 205 nsew signal output
rlabel metal2 s 117962 0 118018 800 6 iram_din0[6]
port 206 nsew signal output
rlabel metal2 s 118698 0 118754 800 6 iram_din0[7]
port 207 nsew signal output
rlabel metal2 s 119342 0 119398 800 6 iram_din0[8]
port 208 nsew signal output
rlabel metal2 s 119802 0 119858 800 6 iram_din0[9]
port 209 nsew signal output
rlabel metal2 s 113178 0 113234 800 6 iram_dout0[0]
port 210 nsew signal input
rlabel metal2 s 120538 0 120594 800 6 iram_dout0[10]
port 211 nsew signal input
rlabel metal2 s 120998 0 121054 800 6 iram_dout0[11]
port 212 nsew signal input
rlabel metal2 s 121458 0 121514 800 6 iram_dout0[12]
port 213 nsew signal input
rlabel metal2 s 121918 0 121974 800 6 iram_dout0[13]
port 214 nsew signal input
rlabel metal2 s 122378 0 122434 800 6 iram_dout0[14]
port 215 nsew signal input
rlabel metal2 s 122838 0 122894 800 6 iram_dout0[15]
port 216 nsew signal input
rlabel metal2 s 123206 0 123262 800 6 iram_dout0[16]
port 217 nsew signal input
rlabel metal2 s 123666 0 123722 800 6 iram_dout0[17]
port 218 nsew signal input
rlabel metal2 s 124126 0 124182 800 6 iram_dout0[18]
port 219 nsew signal input
rlabel metal2 s 124586 0 124642 800 6 iram_dout0[19]
port 220 nsew signal input
rlabel metal2 s 114098 0 114154 800 6 iram_dout0[1]
port 221 nsew signal input
rlabel metal2 s 125046 0 125102 800 6 iram_dout0[20]
port 222 nsew signal input
rlabel metal2 s 125506 0 125562 800 6 iram_dout0[21]
port 223 nsew signal input
rlabel metal2 s 125966 0 126022 800 6 iram_dout0[22]
port 224 nsew signal input
rlabel metal2 s 126426 0 126482 800 6 iram_dout0[23]
port 225 nsew signal input
rlabel metal2 s 126886 0 126942 800 6 iram_dout0[24]
port 226 nsew signal input
rlabel metal2 s 127346 0 127402 800 6 iram_dout0[25]
port 227 nsew signal input
rlabel metal2 s 127806 0 127862 800 6 iram_dout0[26]
port 228 nsew signal input
rlabel metal2 s 128266 0 128322 800 6 iram_dout0[27]
port 229 nsew signal input
rlabel metal2 s 128726 0 128782 800 6 iram_dout0[28]
port 230 nsew signal input
rlabel metal2 s 129186 0 129242 800 6 iram_dout0[29]
port 231 nsew signal input
rlabel metal2 s 115018 0 115074 800 6 iram_dout0[2]
port 232 nsew signal input
rlabel metal2 s 129646 0 129702 800 6 iram_dout0[30]
port 233 nsew signal input
rlabel metal2 s 130106 0 130162 800 6 iram_dout0[31]
port 234 nsew signal input
rlabel metal2 s 115938 0 115994 800 6 iram_dout0[3]
port 235 nsew signal input
rlabel metal2 s 116858 0 116914 800 6 iram_dout0[4]
port 236 nsew signal input
rlabel metal2 s 117502 0 117558 800 6 iram_dout0[5]
port 237 nsew signal input
rlabel metal2 s 118238 0 118294 800 6 iram_dout0[6]
port 238 nsew signal input
rlabel metal2 s 118882 0 118938 800 6 iram_dout0[7]
port 239 nsew signal input
rlabel metal2 s 119618 0 119674 800 6 iram_dout0[8]
port 240 nsew signal input
rlabel metal2 s 120078 0 120134 800 6 iram_dout0[9]
port 241 nsew signal input
rlabel metal2 s 112534 0 112590 800 6 iram_web0
port 242 nsew signal output
rlabel metal2 s 113454 0 113510 800 6 iram_wmask0[0]
port 243 nsew signal output
rlabel metal2 s 114374 0 114430 800 6 iram_wmask0[1]
port 244 nsew signal output
rlabel metal2 s 115294 0 115350 800 6 iram_wmask0[2]
port 245 nsew signal output
rlabel metal2 s 116122 0 116178 800 6 iram_wmask0[3]
port 246 nsew signal output
rlabel metal2 s 24306 0 24362 800 6 la_data_in[0]
port 247 nsew signal input
rlabel metal2 s 92846 0 92902 800 6 la_data_in[100]
port 248 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 la_data_in[101]
port 249 nsew signal input
rlabel metal2 s 94226 0 94282 800 6 la_data_in[102]
port 250 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 la_data_in[103]
port 251 nsew signal input
rlabel metal2 s 95606 0 95662 800 6 la_data_in[104]
port 252 nsew signal input
rlabel metal2 s 96250 0 96306 800 6 la_data_in[105]
port 253 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 la_data_in[106]
port 254 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 la_data_in[107]
port 255 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 la_data_in[108]
port 256 nsew signal input
rlabel metal2 s 99010 0 99066 800 6 la_data_in[109]
port 257 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 la_data_in[10]
port 258 nsew signal input
rlabel metal2 s 99746 0 99802 800 6 la_data_in[110]
port 259 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 la_data_in[111]
port 260 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 la_data_in[112]
port 261 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 la_data_in[113]
port 262 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 la_data_in[114]
port 263 nsew signal input
rlabel metal2 s 103150 0 103206 800 6 la_data_in[115]
port 264 nsew signal input
rlabel metal2 s 103794 0 103850 800 6 la_data_in[116]
port 265 nsew signal input
rlabel metal2 s 104530 0 104586 800 6 la_data_in[117]
port 266 nsew signal input
rlabel metal2 s 105174 0 105230 800 6 la_data_in[118]
port 267 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 la_data_in[119]
port 268 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 la_data_in[11]
port 269 nsew signal input
rlabel metal2 s 106554 0 106610 800 6 la_data_in[120]
port 270 nsew signal input
rlabel metal2 s 107290 0 107346 800 6 la_data_in[121]
port 271 nsew signal input
rlabel metal2 s 107934 0 107990 800 6 la_data_in[122]
port 272 nsew signal input
rlabel metal2 s 108670 0 108726 800 6 la_data_in[123]
port 273 nsew signal input
rlabel metal2 s 109314 0 109370 800 6 la_data_in[124]
port 274 nsew signal input
rlabel metal2 s 109958 0 110014 800 6 la_data_in[125]
port 275 nsew signal input
rlabel metal2 s 110694 0 110750 800 6 la_data_in[126]
port 276 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 la_data_in[127]
port 277 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 la_data_in[12]
port 278 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 la_data_in[13]
port 279 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 la_data_in[14]
port 280 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 la_data_in[15]
port 281 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 la_data_in[16]
port 282 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 la_data_in[17]
port 283 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 la_data_in[18]
port 284 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 la_data_in[19]
port 285 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 la_data_in[1]
port 286 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 la_data_in[20]
port 287 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 la_data_in[21]
port 288 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 la_data_in[22]
port 289 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 la_data_in[23]
port 290 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 la_data_in[24]
port 291 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 la_data_in[25]
port 292 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 la_data_in[26]
port 293 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 la_data_in[27]
port 294 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 la_data_in[28]
port 295 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 la_data_in[29]
port 296 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 la_data_in[2]
port 297 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 la_data_in[30]
port 298 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 la_data_in[31]
port 299 nsew signal input
rlabel metal2 s 46202 0 46258 800 6 la_data_in[32]
port 300 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 la_data_in[33]
port 301 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 la_data_in[34]
port 302 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 la_data_in[35]
port 303 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 la_data_in[36]
port 304 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 la_data_in[37]
port 305 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 la_data_in[38]
port 306 nsew signal input
rlabel metal2 s 50986 0 51042 800 6 la_data_in[39]
port 307 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 la_data_in[3]
port 308 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 la_data_in[40]
port 309 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 la_data_in[41]
port 310 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 la_data_in[42]
port 311 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 la_data_in[43]
port 312 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 la_data_in[44]
port 313 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 la_data_in[45]
port 314 nsew signal input
rlabel metal2 s 55862 0 55918 800 6 la_data_in[46]
port 315 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 la_data_in[47]
port 316 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 la_data_in[48]
port 317 nsew signal input
rlabel metal2 s 57886 0 57942 800 6 la_data_in[49]
port 318 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 la_data_in[4]
port 319 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 la_data_in[50]
port 320 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 la_data_in[51]
port 321 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 la_data_in[52]
port 322 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 la_data_in[53]
port 323 nsew signal input
rlabel metal2 s 61290 0 61346 800 6 la_data_in[54]
port 324 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 la_data_in[55]
port 325 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 la_data_in[56]
port 326 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 la_data_in[57]
port 327 nsew signal input
rlabel metal2 s 64050 0 64106 800 6 la_data_in[58]
port 328 nsew signal input
rlabel metal2 s 64786 0 64842 800 6 la_data_in[59]
port 329 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 la_data_in[5]
port 330 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 la_data_in[60]
port 331 nsew signal input
rlabel metal2 s 66074 0 66130 800 6 la_data_in[61]
port 332 nsew signal input
rlabel metal2 s 66810 0 66866 800 6 la_data_in[62]
port 333 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 la_data_in[63]
port 334 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 la_data_in[64]
port 335 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 la_data_in[65]
port 336 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 la_data_in[66]
port 337 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 la_data_in[67]
port 338 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 la_data_in[68]
port 339 nsew signal input
rlabel metal2 s 71594 0 71650 800 6 la_data_in[69]
port 340 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 la_data_in[6]
port 341 nsew signal input
rlabel metal2 s 72330 0 72386 800 6 la_data_in[70]
port 342 nsew signal input
rlabel metal2 s 72974 0 73030 800 6 la_data_in[71]
port 343 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 la_data_in[72]
port 344 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 la_data_in[73]
port 345 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_data_in[74]
port 346 nsew signal input
rlabel metal2 s 75734 0 75790 800 6 la_data_in[75]
port 347 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 la_data_in[76]
port 348 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 la_data_in[77]
port 349 nsew signal input
rlabel metal2 s 77758 0 77814 800 6 la_data_in[78]
port 350 nsew signal input
rlabel metal2 s 78494 0 78550 800 6 la_data_in[79]
port 351 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 la_data_in[7]
port 352 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 la_data_in[80]
port 353 nsew signal input
rlabel metal2 s 79782 0 79838 800 6 la_data_in[81]
port 354 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_data_in[82]
port 355 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 la_data_in[83]
port 356 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 la_data_in[84]
port 357 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 la_data_in[85]
port 358 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 la_data_in[86]
port 359 nsew signal input
rlabel metal2 s 83922 0 83978 800 6 la_data_in[87]
port 360 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 la_data_in[88]
port 361 nsew signal input
rlabel metal2 s 85302 0 85358 800 6 la_data_in[89]
port 362 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 la_data_in[8]
port 363 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 la_data_in[90]
port 364 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 la_data_in[91]
port 365 nsew signal input
rlabel metal2 s 87326 0 87382 800 6 la_data_in[92]
port 366 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 la_data_in[93]
port 367 nsew signal input
rlabel metal2 s 88706 0 88762 800 6 la_data_in[94]
port 368 nsew signal input
rlabel metal2 s 89442 0 89498 800 6 la_data_in[95]
port 369 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 la_data_in[96]
port 370 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 la_data_in[97]
port 371 nsew signal input
rlabel metal2 s 91466 0 91522 800 6 la_data_in[98]
port 372 nsew signal input
rlabel metal2 s 92202 0 92258 800 6 la_data_in[99]
port 373 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 la_data_in[9]
port 374 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 la_data_out[0]
port 375 nsew signal output
rlabel metal2 s 93122 0 93178 800 6 la_data_out[100]
port 376 nsew signal output
rlabel metal2 s 93766 0 93822 800 6 la_data_out[101]
port 377 nsew signal output
rlabel metal2 s 94410 0 94466 800 6 la_data_out[102]
port 378 nsew signal output
rlabel metal2 s 95146 0 95202 800 6 la_data_out[103]
port 379 nsew signal output
rlabel metal2 s 95790 0 95846 800 6 la_data_out[104]
port 380 nsew signal output
rlabel metal2 s 96526 0 96582 800 6 la_data_out[105]
port 381 nsew signal output
rlabel metal2 s 97170 0 97226 800 6 la_data_out[106]
port 382 nsew signal output
rlabel metal2 s 97906 0 97962 800 6 la_data_out[107]
port 383 nsew signal output
rlabel metal2 s 98550 0 98606 800 6 la_data_out[108]
port 384 nsew signal output
rlabel metal2 s 99286 0 99342 800 6 la_data_out[109]
port 385 nsew signal output
rlabel metal2 s 31390 0 31446 800 6 la_data_out[10]
port 386 nsew signal output
rlabel metal2 s 99930 0 99986 800 6 la_data_out[110]
port 387 nsew signal output
rlabel metal2 s 100666 0 100722 800 6 la_data_out[111]
port 388 nsew signal output
rlabel metal2 s 101310 0 101366 800 6 la_data_out[112]
port 389 nsew signal output
rlabel metal2 s 101954 0 102010 800 6 la_data_out[113]
port 390 nsew signal output
rlabel metal2 s 102690 0 102746 800 6 la_data_out[114]
port 391 nsew signal output
rlabel metal2 s 103334 0 103390 800 6 la_data_out[115]
port 392 nsew signal output
rlabel metal2 s 104070 0 104126 800 6 la_data_out[116]
port 393 nsew signal output
rlabel metal2 s 104714 0 104770 800 6 la_data_out[117]
port 394 nsew signal output
rlabel metal2 s 105450 0 105506 800 6 la_data_out[118]
port 395 nsew signal output
rlabel metal2 s 106094 0 106150 800 6 la_data_out[119]
port 396 nsew signal output
rlabel metal2 s 32034 0 32090 800 6 la_data_out[11]
port 397 nsew signal output
rlabel metal2 s 106830 0 106886 800 6 la_data_out[120]
port 398 nsew signal output
rlabel metal2 s 107474 0 107530 800 6 la_data_out[121]
port 399 nsew signal output
rlabel metal2 s 108210 0 108266 800 6 la_data_out[122]
port 400 nsew signal output
rlabel metal2 s 108854 0 108910 800 6 la_data_out[123]
port 401 nsew signal output
rlabel metal2 s 109498 0 109554 800 6 la_data_out[124]
port 402 nsew signal output
rlabel metal2 s 110234 0 110290 800 6 la_data_out[125]
port 403 nsew signal output
rlabel metal2 s 110878 0 110934 800 6 la_data_out[126]
port 404 nsew signal output
rlabel metal2 s 111614 0 111670 800 6 la_data_out[127]
port 405 nsew signal output
rlabel metal2 s 32770 0 32826 800 6 la_data_out[12]
port 406 nsew signal output
rlabel metal2 s 33414 0 33470 800 6 la_data_out[13]
port 407 nsew signal output
rlabel metal2 s 34150 0 34206 800 6 la_data_out[14]
port 408 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 la_data_out[15]
port 409 nsew signal output
rlabel metal2 s 35530 0 35586 800 6 la_data_out[16]
port 410 nsew signal output
rlabel metal2 s 36174 0 36230 800 6 la_data_out[17]
port 411 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 la_data_out[18]
port 412 nsew signal output
rlabel metal2 s 37554 0 37610 800 6 la_data_out[19]
port 413 nsew signal output
rlabel metal2 s 25226 0 25282 800 6 la_data_out[1]
port 414 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 la_data_out[20]
port 415 nsew signal output
rlabel metal2 s 38934 0 38990 800 6 la_data_out[21]
port 416 nsew signal output
rlabel metal2 s 39578 0 39634 800 6 la_data_out[22]
port 417 nsew signal output
rlabel metal2 s 40314 0 40370 800 6 la_data_out[23]
port 418 nsew signal output
rlabel metal2 s 40958 0 41014 800 6 la_data_out[24]
port 419 nsew signal output
rlabel metal2 s 41694 0 41750 800 6 la_data_out[25]
port 420 nsew signal output
rlabel metal2 s 42338 0 42394 800 6 la_data_out[26]
port 421 nsew signal output
rlabel metal2 s 43074 0 43130 800 6 la_data_out[27]
port 422 nsew signal output
rlabel metal2 s 43718 0 43774 800 6 la_data_out[28]
port 423 nsew signal output
rlabel metal2 s 44362 0 44418 800 6 la_data_out[29]
port 424 nsew signal output
rlabel metal2 s 25870 0 25926 800 6 la_data_out[2]
port 425 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 la_data_out[30]
port 426 nsew signal output
rlabel metal2 s 45742 0 45798 800 6 la_data_out[31]
port 427 nsew signal output
rlabel metal2 s 46478 0 46534 800 6 la_data_out[32]
port 428 nsew signal output
rlabel metal2 s 47122 0 47178 800 6 la_data_out[33]
port 429 nsew signal output
rlabel metal2 s 47858 0 47914 800 6 la_data_out[34]
port 430 nsew signal output
rlabel metal2 s 48502 0 48558 800 6 la_data_out[35]
port 431 nsew signal output
rlabel metal2 s 49238 0 49294 800 6 la_data_out[36]
port 432 nsew signal output
rlabel metal2 s 49882 0 49938 800 6 la_data_out[37]
port 433 nsew signal output
rlabel metal2 s 50618 0 50674 800 6 la_data_out[38]
port 434 nsew signal output
rlabel metal2 s 51262 0 51318 800 6 la_data_out[39]
port 435 nsew signal output
rlabel metal2 s 26606 0 26662 800 6 la_data_out[3]
port 436 nsew signal output
rlabel metal2 s 51906 0 51962 800 6 la_data_out[40]
port 437 nsew signal output
rlabel metal2 s 52642 0 52698 800 6 la_data_out[41]
port 438 nsew signal output
rlabel metal2 s 53286 0 53342 800 6 la_data_out[42]
port 439 nsew signal output
rlabel metal2 s 54022 0 54078 800 6 la_data_out[43]
port 440 nsew signal output
rlabel metal2 s 54666 0 54722 800 6 la_data_out[44]
port 441 nsew signal output
rlabel metal2 s 55402 0 55458 800 6 la_data_out[45]
port 442 nsew signal output
rlabel metal2 s 56046 0 56102 800 6 la_data_out[46]
port 443 nsew signal output
rlabel metal2 s 56782 0 56838 800 6 la_data_out[47]
port 444 nsew signal output
rlabel metal2 s 57426 0 57482 800 6 la_data_out[48]
port 445 nsew signal output
rlabel metal2 s 58070 0 58126 800 6 la_data_out[49]
port 446 nsew signal output
rlabel metal2 s 27250 0 27306 800 6 la_data_out[4]
port 447 nsew signal output
rlabel metal2 s 58806 0 58862 800 6 la_data_out[50]
port 448 nsew signal output
rlabel metal2 s 59450 0 59506 800 6 la_data_out[51]
port 449 nsew signal output
rlabel metal2 s 60186 0 60242 800 6 la_data_out[52]
port 450 nsew signal output
rlabel metal2 s 60830 0 60886 800 6 la_data_out[53]
port 451 nsew signal output
rlabel metal2 s 61566 0 61622 800 6 la_data_out[54]
port 452 nsew signal output
rlabel metal2 s 62210 0 62266 800 6 la_data_out[55]
port 453 nsew signal output
rlabel metal2 s 62946 0 63002 800 6 la_data_out[56]
port 454 nsew signal output
rlabel metal2 s 63590 0 63646 800 6 la_data_out[57]
port 455 nsew signal output
rlabel metal2 s 64326 0 64382 800 6 la_data_out[58]
port 456 nsew signal output
rlabel metal2 s 64970 0 65026 800 6 la_data_out[59]
port 457 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 la_data_out[5]
port 458 nsew signal output
rlabel metal2 s 65614 0 65670 800 6 la_data_out[60]
port 459 nsew signal output
rlabel metal2 s 66350 0 66406 800 6 la_data_out[61]
port 460 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 la_data_out[62]
port 461 nsew signal output
rlabel metal2 s 67730 0 67786 800 6 la_data_out[63]
port 462 nsew signal output
rlabel metal2 s 68374 0 68430 800 6 la_data_out[64]
port 463 nsew signal output
rlabel metal2 s 69110 0 69166 800 6 la_data_out[65]
port 464 nsew signal output
rlabel metal2 s 69754 0 69810 800 6 la_data_out[66]
port 465 nsew signal output
rlabel metal2 s 70490 0 70546 800 6 la_data_out[67]
port 466 nsew signal output
rlabel metal2 s 71134 0 71190 800 6 la_data_out[68]
port 467 nsew signal output
rlabel metal2 s 71870 0 71926 800 6 la_data_out[69]
port 468 nsew signal output
rlabel metal2 s 28630 0 28686 800 6 la_data_out[6]
port 469 nsew signal output
rlabel metal2 s 72514 0 72570 800 6 la_data_out[70]
port 470 nsew signal output
rlabel metal2 s 73158 0 73214 800 6 la_data_out[71]
port 471 nsew signal output
rlabel metal2 s 73894 0 73950 800 6 la_data_out[72]
port 472 nsew signal output
rlabel metal2 s 74538 0 74594 800 6 la_data_out[73]
port 473 nsew signal output
rlabel metal2 s 75274 0 75330 800 6 la_data_out[74]
port 474 nsew signal output
rlabel metal2 s 75918 0 75974 800 6 la_data_out[75]
port 475 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 la_data_out[76]
port 476 nsew signal output
rlabel metal2 s 77298 0 77354 800 6 la_data_out[77]
port 477 nsew signal output
rlabel metal2 s 78034 0 78090 800 6 la_data_out[78]
port 478 nsew signal output
rlabel metal2 s 78678 0 78734 800 6 la_data_out[79]
port 479 nsew signal output
rlabel metal2 s 29274 0 29330 800 6 la_data_out[7]
port 480 nsew signal output
rlabel metal2 s 79414 0 79470 800 6 la_data_out[80]
port 481 nsew signal output
rlabel metal2 s 80058 0 80114 800 6 la_data_out[81]
port 482 nsew signal output
rlabel metal2 s 80702 0 80758 800 6 la_data_out[82]
port 483 nsew signal output
rlabel metal2 s 81438 0 81494 800 6 la_data_out[83]
port 484 nsew signal output
rlabel metal2 s 82082 0 82138 800 6 la_data_out[84]
port 485 nsew signal output
rlabel metal2 s 82818 0 82874 800 6 la_data_out[85]
port 486 nsew signal output
rlabel metal2 s 83462 0 83518 800 6 la_data_out[86]
port 487 nsew signal output
rlabel metal2 s 84198 0 84254 800 6 la_data_out[87]
port 488 nsew signal output
rlabel metal2 s 84842 0 84898 800 6 la_data_out[88]
port 489 nsew signal output
rlabel metal2 s 85578 0 85634 800 6 la_data_out[89]
port 490 nsew signal output
rlabel metal2 s 30010 0 30066 800 6 la_data_out[8]
port 491 nsew signal output
rlabel metal2 s 86222 0 86278 800 6 la_data_out[90]
port 492 nsew signal output
rlabel metal2 s 86958 0 87014 800 6 la_data_out[91]
port 493 nsew signal output
rlabel metal2 s 87602 0 87658 800 6 la_data_out[92]
port 494 nsew signal output
rlabel metal2 s 88246 0 88302 800 6 la_data_out[93]
port 495 nsew signal output
rlabel metal2 s 88982 0 89038 800 6 la_data_out[94]
port 496 nsew signal output
rlabel metal2 s 89626 0 89682 800 6 la_data_out[95]
port 497 nsew signal output
rlabel metal2 s 90362 0 90418 800 6 la_data_out[96]
port 498 nsew signal output
rlabel metal2 s 91006 0 91062 800 6 la_data_out[97]
port 499 nsew signal output
rlabel metal2 s 91742 0 91798 800 6 la_data_out[98]
port 500 nsew signal output
rlabel metal2 s 92386 0 92442 800 6 la_data_out[99]
port 501 nsew signal output
rlabel metal2 s 30654 0 30710 800 6 la_data_out[9]
port 502 nsew signal output
rlabel metal2 s 24766 0 24822 800 6 la_oenb[0]
port 503 nsew signal input
rlabel metal2 s 93306 0 93362 800 6 la_oenb[100]
port 504 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 la_oenb[101]
port 505 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 la_oenb[102]
port 506 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 la_oenb[103]
port 507 nsew signal input
rlabel metal2 s 96066 0 96122 800 6 la_oenb[104]
port 508 nsew signal input
rlabel metal2 s 96710 0 96766 800 6 la_oenb[105]
port 509 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_oenb[106]
port 510 nsew signal input
rlabel metal2 s 98090 0 98146 800 6 la_oenb[107]
port 511 nsew signal input
rlabel metal2 s 98826 0 98882 800 6 la_oenb[108]
port 512 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 la_oenb[109]
port 513 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 la_oenb[10]
port 514 nsew signal input
rlabel metal2 s 100206 0 100262 800 6 la_oenb[110]
port 515 nsew signal input
rlabel metal2 s 100850 0 100906 800 6 la_oenb[111]
port 516 nsew signal input
rlabel metal2 s 101494 0 101550 800 6 la_oenb[112]
port 517 nsew signal input
rlabel metal2 s 102230 0 102286 800 6 la_oenb[113]
port 518 nsew signal input
rlabel metal2 s 102874 0 102930 800 6 la_oenb[114]
port 519 nsew signal input
rlabel metal2 s 103610 0 103666 800 6 la_oenb[115]
port 520 nsew signal input
rlabel metal2 s 104254 0 104310 800 6 la_oenb[116]
port 521 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 la_oenb[117]
port 522 nsew signal input
rlabel metal2 s 105634 0 105690 800 6 la_oenb[118]
port 523 nsew signal input
rlabel metal2 s 106370 0 106426 800 6 la_oenb[119]
port 524 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 la_oenb[11]
port 525 nsew signal input
rlabel metal2 s 107014 0 107070 800 6 la_oenb[120]
port 526 nsew signal input
rlabel metal2 s 107750 0 107806 800 6 la_oenb[121]
port 527 nsew signal input
rlabel metal2 s 108394 0 108450 800 6 la_oenb[122]
port 528 nsew signal input
rlabel metal2 s 109038 0 109094 800 6 la_oenb[123]
port 529 nsew signal input
rlabel metal2 s 109774 0 109830 800 6 la_oenb[124]
port 530 nsew signal input
rlabel metal2 s 110418 0 110474 800 6 la_oenb[125]
port 531 nsew signal input
rlabel metal2 s 111154 0 111210 800 6 la_oenb[126]
port 532 nsew signal input
rlabel metal2 s 111798 0 111854 800 6 la_oenb[127]
port 533 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 la_oenb[12]
port 534 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 la_oenb[13]
port 535 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 la_oenb[14]
port 536 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 la_oenb[15]
port 537 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 la_oenb[16]
port 538 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 la_oenb[17]
port 539 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 la_oenb[18]
port 540 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 la_oenb[19]
port 541 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 la_oenb[1]
port 542 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 la_oenb[20]
port 543 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 la_oenb[21]
port 544 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 la_oenb[22]
port 545 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 la_oenb[23]
port 546 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 la_oenb[24]
port 547 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 la_oenb[25]
port 548 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 la_oenb[26]
port 549 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 la_oenb[27]
port 550 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 la_oenb[28]
port 551 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 la_oenb[29]
port 552 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 la_oenb[2]
port 553 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 la_oenb[30]
port 554 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 la_oenb[31]
port 555 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 la_oenb[32]
port 556 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 la_oenb[33]
port 557 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 la_oenb[34]
port 558 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 la_oenb[35]
port 559 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 la_oenb[36]
port 560 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 la_oenb[37]
port 561 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 la_oenb[38]
port 562 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 la_oenb[39]
port 563 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 la_oenb[3]
port 564 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 la_oenb[40]
port 565 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 la_oenb[41]
port 566 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 la_oenb[42]
port 567 nsew signal input
rlabel metal2 s 54206 0 54262 800 6 la_oenb[43]
port 568 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 la_oenb[44]
port 569 nsew signal input
rlabel metal2 s 55586 0 55642 800 6 la_oenb[45]
port 570 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 la_oenb[46]
port 571 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 la_oenb[47]
port 572 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 la_oenb[48]
port 573 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 la_oenb[49]
port 574 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 la_oenb[4]
port 575 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 la_oenb[50]
port 576 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 la_oenb[51]
port 577 nsew signal input
rlabel metal2 s 60370 0 60426 800 6 la_oenb[52]
port 578 nsew signal input
rlabel metal2 s 61106 0 61162 800 6 la_oenb[53]
port 579 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 la_oenb[54]
port 580 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 la_oenb[55]
port 581 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 la_oenb[56]
port 582 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 la_oenb[57]
port 583 nsew signal input
rlabel metal2 s 64510 0 64566 800 6 la_oenb[58]
port 584 nsew signal input
rlabel metal2 s 65246 0 65302 800 6 la_oenb[59]
port 585 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 la_oenb[5]
port 586 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 la_oenb[60]
port 587 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 la_oenb[61]
port 588 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 la_oenb[62]
port 589 nsew signal input
rlabel metal2 s 67914 0 67970 800 6 la_oenb[63]
port 590 nsew signal input
rlabel metal2 s 68650 0 68706 800 6 la_oenb[64]
port 591 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 la_oenb[65]
port 592 nsew signal input
rlabel metal2 s 70030 0 70086 800 6 la_oenb[66]
port 593 nsew signal input
rlabel metal2 s 70674 0 70730 800 6 la_oenb[67]
port 594 nsew signal input
rlabel metal2 s 71410 0 71466 800 6 la_oenb[68]
port 595 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_oenb[69]
port 596 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 la_oenb[6]
port 597 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 la_oenb[70]
port 598 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 la_oenb[71]
port 599 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_oenb[72]
port 600 nsew signal input
rlabel metal2 s 74814 0 74870 800 6 la_oenb[73]
port 601 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 la_oenb[74]
port 602 nsew signal input
rlabel metal2 s 76194 0 76250 800 6 la_oenb[75]
port 603 nsew signal input
rlabel metal2 s 76838 0 76894 800 6 la_oenb[76]
port 604 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 la_oenb[77]
port 605 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 la_oenb[78]
port 606 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 la_oenb[79]
port 607 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 la_oenb[7]
port 608 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 la_oenb[80]
port 609 nsew signal input
rlabel metal2 s 80242 0 80298 800 6 la_oenb[81]
port 610 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 la_oenb[82]
port 611 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 la_oenb[83]
port 612 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 la_oenb[84]
port 613 nsew signal input
rlabel metal2 s 83002 0 83058 800 6 la_oenb[85]
port 614 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 la_oenb[86]
port 615 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 la_oenb[87]
port 616 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 la_oenb[88]
port 617 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 la_oenb[89]
port 618 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 la_oenb[8]
port 619 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 la_oenb[90]
port 620 nsew signal input
rlabel metal2 s 87142 0 87198 800 6 la_oenb[91]
port 621 nsew signal input
rlabel metal2 s 87786 0 87842 800 6 la_oenb[92]
port 622 nsew signal input
rlabel metal2 s 88522 0 88578 800 6 la_oenb[93]
port 623 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 la_oenb[94]
port 624 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 la_oenb[95]
port 625 nsew signal input
rlabel metal2 s 90546 0 90602 800 6 la_oenb[96]
port 626 nsew signal input
rlabel metal2 s 91282 0 91338 800 6 la_oenb[97]
port 627 nsew signal input
rlabel metal2 s 91926 0 91982 800 6 la_oenb[98]
port 628 nsew signal input
rlabel metal2 s 92662 0 92718 800 6 la_oenb[99]
port 629 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 la_oenb[9]
port 630 nsew signal input
rlabel metal2 s 62026 131635 62082 132435 6 user_irq[0]
port 631 nsew signal output
rlabel metal2 s 62762 131635 62818 132435 6 user_irq[1]
port 632 nsew signal output
rlabel metal2 s 63590 131635 63646 132435 6 user_irq[2]
port 633 nsew signal output
rlabel metal4 s 4208 2128 4528 130064 6 vccd1
port 634 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 130064 6 vccd1
port 634 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 130064 6 vccd1
port 634 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 130064 6 vccd1
port 634 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 130064 6 vccd1
port 634 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 130064 6 vssd1
port 635 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 130064 6 vssd1
port 635 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 130064 6 vssd1
port 635 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 130064 6 vssd1
port 635 nsew ground bidirectional
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 636 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_rst_i
port 637 nsew signal input
rlabel metal2 s 478 0 534 800 6 wbs_ack_o
port 638 nsew signal output
rlabel metal2 s 1398 0 1454 800 6 wbs_adr_i[0]
port 639 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 wbs_adr_i[10]
port 640 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 wbs_adr_i[11]
port 641 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wbs_adr_i[12]
port 642 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 wbs_adr_i[13]
port 643 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 wbs_adr_i[14]
port 644 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_adr_i[15]
port 645 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 wbs_adr_i[16]
port 646 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 wbs_adr_i[17]
port 647 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 wbs_adr_i[18]
port 648 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 wbs_adr_i[19]
port 649 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_adr_i[1]
port 650 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 wbs_adr_i[20]
port 651 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_adr_i[21]
port 652 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_adr_i[22]
port 653 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wbs_adr_i[23]
port 654 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 wbs_adr_i[24]
port 655 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 wbs_adr_i[25]
port 656 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 wbs_adr_i[26]
port 657 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 wbs_adr_i[27]
port 658 nsew signal input
rlabel metal2 s 21546 0 21602 800 6 wbs_adr_i[28]
port 659 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 wbs_adr_i[29]
port 660 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wbs_adr_i[2]
port 661 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 wbs_adr_i[30]
port 662 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 wbs_adr_i[31]
port 663 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 wbs_adr_i[3]
port 664 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wbs_adr_i[4]
port 665 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wbs_adr_i[5]
port 666 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_adr_i[6]
port 667 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_adr_i[7]
port 668 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 wbs_adr_i[8]
port 669 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_adr_i[9]
port 670 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_cyc_i
port 671 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_dat_i[0]
port 672 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wbs_dat_i[10]
port 673 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 wbs_dat_i[11]
port 674 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 wbs_dat_i[12]
port 675 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 wbs_dat_i[13]
port 676 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 wbs_dat_i[14]
port 677 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 wbs_dat_i[15]
port 678 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 wbs_dat_i[16]
port 679 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wbs_dat_i[17]
port 680 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 wbs_dat_i[18]
port 681 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 wbs_dat_i[19]
port 682 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_i[1]
port 683 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 wbs_dat_i[20]
port 684 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 wbs_dat_i[21]
port 685 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wbs_dat_i[22]
port 686 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 wbs_dat_i[23]
port 687 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 wbs_dat_i[24]
port 688 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 wbs_dat_i[25]
port 689 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wbs_dat_i[26]
port 690 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wbs_dat_i[27]
port 691 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 wbs_dat_i[28]
port 692 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wbs_dat_i[29]
port 693 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wbs_dat_i[2]
port 694 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 wbs_dat_i[30]
port 695 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 wbs_dat_i[31]
port 696 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 wbs_dat_i[3]
port 697 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_dat_i[4]
port 698 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 wbs_dat_i[5]
port 699 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wbs_dat_i[6]
port 700 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_i[7]
port 701 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 wbs_dat_i[8]
port 702 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_dat_i[9]
port 703 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 wbs_dat_o[0]
port 704 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 wbs_dat_o[10]
port 705 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 wbs_dat_o[11]
port 706 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_o[12]
port 707 nsew signal output
rlabel metal2 s 11702 0 11758 800 6 wbs_dat_o[13]
port 708 nsew signal output
rlabel metal2 s 12438 0 12494 800 6 wbs_dat_o[14]
port 709 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 wbs_dat_o[15]
port 710 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 wbs_dat_o[16]
port 711 nsew signal output
rlabel metal2 s 14462 0 14518 800 6 wbs_dat_o[17]
port 712 nsew signal output
rlabel metal2 s 15106 0 15162 800 6 wbs_dat_o[18]
port 713 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 wbs_dat_o[19]
port 714 nsew signal output
rlabel metal2 s 2778 0 2834 800 6 wbs_dat_o[1]
port 715 nsew signal output
rlabel metal2 s 16486 0 16542 800 6 wbs_dat_o[20]
port 716 nsew signal output
rlabel metal2 s 17222 0 17278 800 6 wbs_dat_o[21]
port 717 nsew signal output
rlabel metal2 s 17866 0 17922 800 6 wbs_dat_o[22]
port 718 nsew signal output
rlabel metal2 s 18602 0 18658 800 6 wbs_dat_o[23]
port 719 nsew signal output
rlabel metal2 s 19246 0 19302 800 6 wbs_dat_o[24]
port 720 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 wbs_dat_o[25]
port 721 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_o[26]
port 722 nsew signal output
rlabel metal2 s 21362 0 21418 800 6 wbs_dat_o[27]
port 723 nsew signal output
rlabel metal2 s 22006 0 22062 800 6 wbs_dat_o[28]
port 724 nsew signal output
rlabel metal2 s 22650 0 22706 800 6 wbs_dat_o[29]
port 725 nsew signal output
rlabel metal2 s 3698 0 3754 800 6 wbs_dat_o[2]
port 726 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 wbs_dat_o[30]
port 727 nsew signal output
rlabel metal2 s 24030 0 24086 800 6 wbs_dat_o[31]
port 728 nsew signal output
rlabel metal2 s 4618 0 4674 800 6 wbs_dat_o[3]
port 729 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_o[4]
port 730 nsew signal output
rlabel metal2 s 6274 0 6330 800 6 wbs_dat_o[5]
port 731 nsew signal output
rlabel metal2 s 6918 0 6974 800 6 wbs_dat_o[6]
port 732 nsew signal output
rlabel metal2 s 7562 0 7618 800 6 wbs_dat_o[7]
port 733 nsew signal output
rlabel metal2 s 8298 0 8354 800 6 wbs_dat_o[8]
port 734 nsew signal output
rlabel metal2 s 8942 0 8998 800 6 wbs_dat_o[9]
port 735 nsew signal output
rlabel metal2 s 2134 0 2190 800 6 wbs_sel_i[0]
port 736 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_sel_i[1]
port 737 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wbs_sel_i[2]
port 738 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 wbs_sel_i[3]
port 739 nsew signal input
rlabel metal2 s 938 0 994 800 6 wbs_stb_i
port 740 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 wbs_we_i
port 741 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 130291 132435
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 43554670
string GDS_FILE /home/jure/Projekti/rvj1-caravel-soc/openlane/rvj1_caravel_soc/runs/rvj1_caravel_soc/results/signoff/rvj1_caravel_soc.magic.gds
string GDS_START 1268210
<< end >>

