VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO rvj1_caravel_soc
  CLASS BLOCK ;
  FOREIGN rvj1_caravel_soc ;
  ORIGIN 0.000 0.000 ;
  SIZE 591.480 BY 602.200 ;
  PIN dram_addr0[-1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 0.000 515.110 4.000 ;
    END
  END dram_addr0[-1]
  PIN dram_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 598.200 50.510 602.200 ;
    END
  END dram_addr0[0]
  PIN dram_clk0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 6.840 591.480 7.440 ;
    END
  END dram_clk0
  PIN dram_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 598.200 7.270 602.200 ;
    END
  END dram_csb0
  PIN dram_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END dram_din0[0]
  PIN dram_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 339.360 4.000 339.960 ;
    END
  END dram_din0[10]
  PIN dram_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 598.200 237.730 602.200 ;
    END
  END dram_din0[11]
  PIN dram_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 598.200 252.450 602.200 ;
    END
  END dram_din0[12]
  PIN dram_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 598.200 295.690 602.200 ;
    END
  END dram_din0[13]
  PIN dram_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 293.800 591.480 294.400 ;
    END
  END dram_din0[14]
  PIN dram_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.560 4.000 418.160 ;
    END
  END dram_din0[15]
  PIN dram_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 308.080 591.480 308.680 ;
    END
  END dram_din0[16]
  PIN dram_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.770 0.000 556.050 4.000 ;
    END
  END dram_din0[17]
  PIN dram_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 4.000 437.200 ;
    END
  END dram_din0[18]
  PIN dram_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.530 0.000 558.810 4.000 ;
    END
  END dram_din0[19]
  PIN dram_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.430 0.000 519.710 4.000 ;
    END
  END dram_din0[1]
  PIN dram_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 598.200 396.430 602.200 ;
    END
  END dram_din0[20]
  PIN dram_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 417.560 591.480 418.160 ;
    END
  END dram_din0[21]
  PIN dram_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.080 4.000 495.680 ;
    END
  END dram_din0[22]
  PIN dram_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 598.200 425.410 602.200 ;
    END
  END dram_din0[23]
  PIN dram_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 485.560 591.480 486.160 ;
    END
  END dram_din0[24]
  PIN dram_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 499.160 591.480 499.760 ;
    END
  END dram_din0[25]
  PIN dram_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 513.440 591.480 514.040 ;
    END
  END dram_din0[26]
  PIN dram_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.550 0.000 575.830 4.000 ;
    END
  END dram_din0[27]
  PIN dram_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.850 0.000 578.130 4.000 ;
    END
  END dram_din0[28]
  PIN dram_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.450 0.000 582.730 4.000 ;
    END
  END dram_din0[29]
  PIN dram_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 598.200 136.990 602.200 ;
    END
  END dram_din0[2]
  PIN dram_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 0.000 585.490 4.000 ;
    END
  END dram_din0[30]
  PIN dram_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 581.440 591.480 582.040 ;
    END
  END dram_din0[31]
  PIN dram_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.850 0.000 532.130 4.000 ;
    END
  END dram_din0[3]
  PIN dram_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.450 0.000 536.730 4.000 ;
    END
  END dram_din0[4]
  PIN dram_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END dram_din0[5]
  PIN dram_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 170.720 591.480 171.320 ;
    END
  END dram_din0[6]
  PIN dram_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 197.920 591.480 198.520 ;
    END
  END dram_din0[7]
  PIN dram_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 212.200 591.480 212.800 ;
    END
  END dram_din0[8]
  PIN dram_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 225.800 591.480 226.400 ;
    END
  END dram_din0[9]
  PIN dram_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 598.200 64.770 602.200 ;
    END
  END dram_dout0[0]
  PIN dram_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 598.200 194.490 602.200 ;
    END
  END dram_dout0[10]
  PIN dram_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 253.000 591.480 253.600 ;
    END
  END dram_dout0[11]
  PIN dram_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 598.200 266.710 602.200 ;
    END
  END dram_dout0[12]
  PIN dram_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 598.200 309.950 602.200 ;
    END
  END dram_dout0[13]
  PIN dram_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.800 4.000 379.400 ;
    END
  END dram_dout0[14]
  PIN dram_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.390 598.200 324.670 602.200 ;
    END
  END dram_dout0[15]
  PIN dram_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 321.680 591.480 322.280 ;
    END
  END dram_dout0[16]
  PIN dram_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.910 598.200 353.190 602.200 ;
    END
  END dram_dout0[17]
  PIN dram_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 362.480 591.480 363.080 ;
    END
  END dram_dout0[18]
  PIN dram_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.830 0.000 561.110 4.000 ;
    END
  END dram_dout0[19]
  PIN dram_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 0.000 522.470 4.000 ;
    END
  END dram_dout0[1]
  PIN dram_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 403.280 591.480 403.880 ;
    END
  END dram_dout0[20]
  PIN dram_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 431.160 591.480 431.760 ;
    END
  END dram_dout0[21]
  PIN dram_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.870 598.200 411.150 602.200 ;
    END
  END dram_dout0[22]
  PIN dram_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 598.200 439.670 602.200 ;
    END
  END dram_dout0[23]
  PIN dram_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.840 4.000 534.440 ;
    END
  END dram_dout0[24]
  PIN dram_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.490 0.000 570.770 4.000 ;
    END
  END dram_dout0[25]
  PIN dram_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.790 0.000 573.070 4.000 ;
    END
  END dram_dout0[26]
  PIN dram_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.330 598.200 526.610 602.200 ;
    END
  END dram_dout0[27]
  PIN dram_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 527.040 591.480 527.640 ;
    END
  END dram_dout0[28]
  PIN dram_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 572.600 4.000 573.200 ;
    END
  END dram_dout0[29]
  PIN dram_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END dram_dout0[2]
  PIN dram_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 554.240 591.480 554.840 ;
    END
  END dram_dout0[30]
  PIN dram_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.510 0.000 587.790 4.000 ;
    END
  END dram_dout0[31]
  PIN dram_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END dram_dout0[3]
  PIN dram_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 116.320 591.480 116.920 ;
    END
  END dram_dout0[4]
  PIN dram_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END dram_dout0[5]
  PIN dram_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END dram_dout0[6]
  PIN dram_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 0.000 539.490 4.000 ;
    END
  END dram_dout0[7]
  PIN dram_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.560 4.000 282.160 ;
    END
  END dram_dout0[8]
  PIN dram_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 239.400 591.480 240.000 ;
    END
  END dram_dout0[9]
  PIN dram_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END dram_web0
  PIN dram_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 598.200 79.030 602.200 ;
    END
  END dram_wmask0[0]
  PIN dram_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END dram_wmask0[1]
  PIN dram_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.790 0.000 527.070 4.000 ;
    END
  END dram_wmask0[2]
  PIN dram_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 88.440 591.480 89.040 ;
    END
  END dram_wmask0[3]
  PIN iram_addr0[-1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 598.200 21.530 602.200 ;
    END
  END iram_addr0[-1]
  PIN iram_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 598.200 93.750 602.200 ;
    END
  END iram_addr0[0]
  PIN iram_clk0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.130 0.000 517.410 4.000 ;
    END
  END iram_clk0
  PIN iram_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 20.440 591.480 21.040 ;
    END
  END iram_csb0
  PIN iram_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 598.200 108.010 602.200 ;
    END
  END iram_din0[0]
  PIN iram_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 598.200 209.210 602.200 ;
    END
  END iram_din0[10]
  PIN iram_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 266.600 591.480 267.200 ;
    END
  END iram_din0[11]
  PIN iram_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 0.000 544.090 4.000 ;
    END
  END iram_din0[12]
  PIN iram_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.080 4.000 359.680 ;
    END
  END iram_din0[13]
  PIN iram_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END iram_din0[14]
  PIN iram_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.170 0.000 551.450 4.000 ;
    END
  END iram_din0[15]
  PIN iram_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 0.000 553.750 4.000 ;
    END
  END iram_din0[16]
  PIN iram_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.630 598.200 367.910 602.200 ;
    END
  END iram_din0[17]
  PIN iram_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 376.080 591.480 376.680 ;
    END
  END iram_din0[18]
  PIN iram_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.130 0.000 563.410 4.000 ;
    END
  END iram_din0[19]
  PIN iram_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 61.240 591.480 61.840 ;
    END
  END iram_din0[1]
  PIN iram_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.890 0.000 566.170 4.000 ;
    END
  END iram_din0[20]
  PIN iram_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 475.360 4.000 475.960 ;
    END
  END iram_din0[21]
  PIN iram_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.800 4.000 515.400 ;
    END
  END iram_din0[22]
  PIN iram_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 598.200 454.390 602.200 ;
    END
  END iram_din0[23]
  PIN iram_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.190 0.000 568.470 4.000 ;
    END
  END iram_din0[24]
  PIN iram_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 598.200 483.370 602.200 ;
    END
  END iram_din0[25]
  PIN iram_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.350 598.200 497.630 602.200 ;
    END
  END iram_din0[26]
  PIN iram_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.590 598.200 540.870 602.200 ;
    END
  END iram_din0[27]
  PIN iram_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 598.200 569.850 602.200 ;
    END
  END iram_din0[28]
  PIN iram_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.830 598.200 584.110 602.200 ;
    END
  END iram_din0[29]
  PIN iram_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 74.840 591.480 75.440 ;
    END
  END iram_din0[2]
  PIN iram_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 592.320 4.000 592.920 ;
    END
  END iram_din0[30]
  PIN iram_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 595.040 591.480 595.640 ;
    END
  END iram_din0[31]
  PIN iram_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.150 0.000 534.430 4.000 ;
    END
  END iram_din0[3]
  PIN iram_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 129.920 591.480 130.520 ;
    END
  END iram_din0[4]
  PIN iram_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 203.360 4.000 203.960 ;
    END
  END iram_din0[5]
  PIN iram_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 184.320 591.480 184.920 ;
    END
  END iram_din0[6]
  PIN iram_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.510 0.000 541.790 4.000 ;
    END
  END iram_din0[7]
  PIN iram_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END iram_din0[8]
  PIN iram_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 598.200 165.970 602.200 ;
    END
  END iram_din0[9]
  PIN iram_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 4.000 67.960 ;
    END
  END iram_dout0[0]
  PIN iram_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 598.200 223.470 602.200 ;
    END
  END iram_dout0[10]
  PIN iram_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 280.200 591.480 280.800 ;
    END
  END iram_dout0[11]
  PIN iram_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 598.200 280.970 602.200 ;
    END
  END iram_dout0[12]
  PIN iram_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.110 0.000 546.390 4.000 ;
    END
  END iram_dout0[13]
  PIN iram_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.870 0.000 549.150 4.000 ;
    END
  END iram_dout0[14]
  PIN iram_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 598.200 338.930 602.200 ;
    END
  END iram_dout0[15]
  PIN iram_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 335.280 591.480 335.880 ;
    END
  END iram_dout0[16]
  PIN iram_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 348.880 591.480 349.480 ;
    END
  END iram_dout0[17]
  PIN iram_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 598.200 382.170 602.200 ;
    END
  END iram_dout0[18]
  PIN iram_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 389.680 591.480 390.280 ;
    END
  END iram_dout0[19]
  PIN iram_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 0.000 524.770 4.000 ;
    END
  END iram_dout0[1]
  PIN iram_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 456.320 4.000 456.920 ;
    END
  END iram_dout0[20]
  PIN iram_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 444.760 591.480 445.360 ;
    END
  END iram_dout0[21]
  PIN iram_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 458.360 591.480 458.960 ;
    END
  END iram_dout0[22]
  PIN iram_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 471.960 591.480 472.560 ;
    END
  END iram_dout0[23]
  PIN iram_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.370 598.200 468.650 602.200 ;
    END
  END iram_dout0[24]
  PIN iram_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 553.560 4.000 554.160 ;
    END
  END iram_dout0[25]
  PIN iram_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.610 598.200 511.890 602.200 ;
    END
  END iram_dout0[26]
  PIN iram_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.850 598.200 555.130 602.200 ;
    END
  END iram_dout0[27]
  PIN iram_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.150 0.000 580.430 4.000 ;
    END
  END iram_dout0[28]
  PIN iram_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 540.640 591.480 541.240 ;
    END
  END iram_dout0[29]
  PIN iram_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END iram_dout0[2]
  PIN iram_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 567.840 591.480 568.440 ;
    END
  END iram_dout0[30]
  PIN iram_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.810 0.000 590.090 4.000 ;
    END
  END iram_dout0[31]
  PIN iram_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 102.040 591.480 102.640 ;
    END
  END iram_dout0[3]
  PIN iram_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 143.520 591.480 144.120 ;
    END
  END iram_dout0[4]
  PIN iram_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 157.120 591.480 157.720 ;
    END
  END iram_dout0[5]
  PIN iram_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END iram_dout0[6]
  PIN iram_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END iram_dout0[7]
  PIN iram_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 320.320 4.000 320.920 ;
    END
  END iram_dout0[8]
  PIN iram_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 598.200 180.230 602.200 ;
    END
  END iram_dout0[9]
  PIN iram_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 34.040 591.480 34.640 ;
    END
  END iram_web0
  PIN iram_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 587.480 47.640 591.480 48.240 ;
    END
  END iram_wmask0[0]
  PIN iram_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 598.200 122.270 602.200 ;
    END
  END iram_wmask0[1]
  PIN iram_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.090 0.000 529.370 4.000 ;
    END
  END iram_wmask0[2]
  PIN iram_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 598.200 151.250 602.200 ;
    END
  END iram_wmask0[3]
  PIN jedro_1_rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END jedro_1_rstn
  PIN sel_wb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 598.200 35.790 602.200 ;
    END
  END sel_wb
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 590.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 590.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 590.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 590.480 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 590.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 590.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 590.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 590.480 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.010 0.000 1.290 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END wb_rst_i
  PIN wb_uart_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 4.000 ;
    END
  END wb_uart_ack
  PIN wb_uart_adr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END wb_uart_adr[0]
  PIN wb_uart_adr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 4.000 ;
    END
  END wb_uart_adr[10]
  PIN wb_uart_adr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 0.000 110.310 4.000 ;
    END
  END wb_uart_adr[11]
  PIN wb_uart_adr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END wb_uart_adr[12]
  PIN wb_uart_adr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END wb_uart_adr[13]
  PIN wb_uart_adr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END wb_uart_adr[14]
  PIN wb_uart_adr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 4.000 ;
    END
  END wb_uart_adr[15]
  PIN wb_uart_adr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 4.000 ;
    END
  END wb_uart_adr[16]
  PIN wb_uart_adr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 0.000 154.010 4.000 ;
    END
  END wb_uart_adr[17]
  PIN wb_uart_adr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END wb_uart_adr[18]
  PIN wb_uart_adr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 4.000 ;
    END
  END wb_uart_adr[19]
  PIN wb_uart_adr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END wb_uart_adr[1]
  PIN wb_uart_adr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END wb_uart_adr[20]
  PIN wb_uart_adr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 0.000 182.990 4.000 ;
    END
  END wb_uart_adr[21]
  PIN wb_uart_adr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END wb_uart_adr[22]
  PIN wb_uart_adr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 4.000 ;
    END
  END wb_uart_adr[23]
  PIN wb_uart_adr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 0.000 204.610 4.000 ;
    END
  END wb_uart_adr[24]
  PIN wb_uart_adr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 0.000 211.970 4.000 ;
    END
  END wb_uart_adr[25]
  PIN wb_uart_adr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END wb_uart_adr[26]
  PIN wb_uart_adr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END wb_uart_adr[27]
  PIN wb_uart_adr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 0.000 233.590 4.000 ;
    END
  END wb_uart_adr[28]
  PIN wb_uart_adr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 0.000 240.950 4.000 ;
    END
  END wb_uart_adr[29]
  PIN wb_uart_adr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END wb_uart_adr[2]
  PIN wb_uart_adr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END wb_uart_adr[30]
  PIN wb_uart_adr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 0.000 255.670 4.000 ;
    END
  END wb_uart_adr[31]
  PIN wb_uart_adr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 4.000 ;
    END
  END wb_uart_adr[3]
  PIN wb_uart_adr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END wb_uart_adr[4]
  PIN wb_uart_adr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END wb_uart_adr[5]
  PIN wb_uart_adr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END wb_uart_adr[6]
  PIN wb_uart_adr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END wb_uart_adr[7]
  PIN wb_uart_adr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 4.000 ;
    END
  END wb_uart_adr[8]
  PIN wb_uart_adr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 4.000 ;
    END
  END wb_uart_adr[9]
  PIN wb_uart_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 0.000 8.190 4.000 ;
    END
  END wb_uart_clk
  PIN wb_uart_cyc
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 0.000 10.950 4.000 ;
    END
  END wb_uart_cyc
  PIN wb_uart_dat_fromcpu[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END wb_uart_dat_fromcpu[0]
  PIN wb_uart_dat_fromcpu[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END wb_uart_dat_fromcpu[10]
  PIN wb_uart_dat_fromcpu[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END wb_uart_dat_fromcpu[11]
  PIN wb_uart_dat_fromcpu[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END wb_uart_dat_fromcpu[12]
  PIN wb_uart_dat_fromcpu[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END wb_uart_dat_fromcpu[13]
  PIN wb_uart_dat_fromcpu[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 0.000 134.230 4.000 ;
    END
  END wb_uart_dat_fromcpu[14]
  PIN wb_uart_dat_fromcpu[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 0.000 141.590 4.000 ;
    END
  END wb_uart_dat_fromcpu[15]
  PIN wb_uart_dat_fromcpu[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 0.000 148.950 4.000 ;
    END
  END wb_uart_dat_fromcpu[16]
  PIN wb_uart_dat_fromcpu[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 0.000 156.310 4.000 ;
    END
  END wb_uart_dat_fromcpu[17]
  PIN wb_uart_dat_fromcpu[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END wb_uart_dat_fromcpu[18]
  PIN wb_uart_dat_fromcpu[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END wb_uart_dat_fromcpu[19]
  PIN wb_uart_dat_fromcpu[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END wb_uart_dat_fromcpu[1]
  PIN wb_uart_dat_fromcpu[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 0.000 177.930 4.000 ;
    END
  END wb_uart_dat_fromcpu[20]
  PIN wb_uart_dat_fromcpu[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END wb_uart_dat_fromcpu[21]
  PIN wb_uart_dat_fromcpu[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END wb_uart_dat_fromcpu[22]
  PIN wb_uart_dat_fromcpu[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END wb_uart_dat_fromcpu[23]
  PIN wb_uart_dat_fromcpu[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 0.000 206.910 4.000 ;
    END
  END wb_uart_dat_fromcpu[24]
  PIN wb_uart_dat_fromcpu[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 0.000 214.270 4.000 ;
    END
  END wb_uart_dat_fromcpu[25]
  PIN wb_uart_dat_fromcpu[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 0.000 221.630 4.000 ;
    END
  END wb_uart_dat_fromcpu[26]
  PIN wb_uart_dat_fromcpu[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END wb_uart_dat_fromcpu[27]
  PIN wb_uart_dat_fromcpu[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 0.000 236.350 4.000 ;
    END
  END wb_uart_dat_fromcpu[28]
  PIN wb_uart_dat_fromcpu[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 0.000 243.710 4.000 ;
    END
  END wb_uart_dat_fromcpu[29]
  PIN wb_uart_dat_fromcpu[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END wb_uart_dat_fromcpu[2]
  PIN wb_uart_dat_fromcpu[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 0.000 250.610 4.000 ;
    END
  END wb_uart_dat_fromcpu[30]
  PIN wb_uart_dat_fromcpu[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END wb_uart_dat_fromcpu[31]
  PIN wb_uart_dat_fromcpu[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END wb_uart_dat_fromcpu[3]
  PIN wb_uart_dat_fromcpu[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END wb_uart_dat_fromcpu[4]
  PIN wb_uart_dat_fromcpu[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 4.000 ;
    END
  END wb_uart_dat_fromcpu[5]
  PIN wb_uart_dat_fromcpu[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END wb_uart_dat_fromcpu[6]
  PIN wb_uart_dat_fromcpu[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END wb_uart_dat_fromcpu[7]
  PIN wb_uart_dat_fromcpu[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 4.000 ;
    END
  END wb_uart_dat_fromcpu[8]
  PIN wb_uart_dat_fromcpu[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END wb_uart_dat_fromcpu[9]
  PIN wb_uart_dat_tocpu[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END wb_uart_dat_tocpu[0]
  PIN wb_uart_dat_tocpu[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END wb_uart_dat_tocpu[10]
  PIN wb_uart_dat_tocpu[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 4.000 ;
    END
  END wb_uart_dat_tocpu[11]
  PIN wb_uart_dat_tocpu[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 4.000 ;
    END
  END wb_uart_dat_tocpu[12]
  PIN wb_uart_dat_tocpu[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 4.000 ;
    END
  END wb_uart_dat_tocpu[13]
  PIN wb_uart_dat_tocpu[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 4.000 ;
    END
  END wb_uart_dat_tocpu[14]
  PIN wb_uart_dat_tocpu[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 4.000 ;
    END
  END wb_uart_dat_tocpu[15]
  PIN wb_uart_dat_tocpu[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END wb_uart_dat_tocpu[16]
  PIN wb_uart_dat_tocpu[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 0.000 158.610 4.000 ;
    END
  END wb_uart_dat_tocpu[17]
  PIN wb_uart_dat_tocpu[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END wb_uart_dat_tocpu[18]
  PIN wb_uart_dat_tocpu[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.330 4.000 ;
    END
  END wb_uart_dat_tocpu[19]
  PIN wb_uart_dat_tocpu[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END wb_uart_dat_tocpu[1]
  PIN wb_uart_dat_tocpu[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END wb_uart_dat_tocpu[20]
  PIN wb_uart_dat_tocpu[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 0.000 187.590 4.000 ;
    END
  END wb_uart_dat_tocpu[21]
  PIN wb_uart_dat_tocpu[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 0.000 194.950 4.000 ;
    END
  END wb_uart_dat_tocpu[22]
  PIN wb_uart_dat_tocpu[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 0.000 202.310 4.000 ;
    END
  END wb_uart_dat_tocpu[23]
  PIN wb_uart_dat_tocpu[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END wb_uart_dat_tocpu[24]
  PIN wb_uart_dat_tocpu[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 0.000 217.030 4.000 ;
    END
  END wb_uart_dat_tocpu[25]
  PIN wb_uart_dat_tocpu[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 0.000 223.930 4.000 ;
    END
  END wb_uart_dat_tocpu[26]
  PIN wb_uart_dat_tocpu[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END wb_uart_dat_tocpu[27]
  PIN wb_uart_dat_tocpu[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END wb_uart_dat_tocpu[28]
  PIN wb_uart_dat_tocpu[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 0.000 246.010 4.000 ;
    END
  END wb_uart_dat_tocpu[29]
  PIN wb_uart_dat_tocpu[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END wb_uart_dat_tocpu[2]
  PIN wb_uart_dat_tocpu[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 4.000 ;
    END
  END wb_uart_dat_tocpu[30]
  PIN wb_uart_dat_tocpu[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 0.000 260.270 4.000 ;
    END
  END wb_uart_dat_tocpu[31]
  PIN wb_uart_dat_tocpu[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END wb_uart_dat_tocpu[3]
  PIN wb_uart_dat_tocpu[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 4.000 ;
    END
  END wb_uart_dat_tocpu[4]
  PIN wb_uart_dat_tocpu[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END wb_uart_dat_tocpu[5]
  PIN wb_uart_dat_tocpu[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END wb_uart_dat_tocpu[6]
  PIN wb_uart_dat_tocpu[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END wb_uart_dat_tocpu[7]
  PIN wb_uart_dat_tocpu[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END wb_uart_dat_tocpu[8]
  PIN wb_uart_dat_tocpu[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END wb_uart_dat_tocpu[9]
  PIN wb_uart_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END wb_uart_rst
  PIN wb_uart_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 4.000 ;
    END
  END wb_uart_sel[0]
  PIN wb_uart_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 4.000 ;
    END
  END wb_uart_sel[1]
  PIN wb_uart_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END wb_uart_sel[2]
  PIN wb_uart_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 4.000 ;
    END
  END wb_uart_sel[3]
  PIN wb_uart_stb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 4.000 ;
    END
  END wb_uart_stb
  PIN wb_uart_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END wb_uart_we
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 0.000 263.030 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 0.000 272.690 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 0.000 355.030 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 0.000 362.390 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.470 0.000 369.750 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.370 0.000 376.650 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.730 0.000 384.010 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 0.000 391.370 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.450 0.000 398.730 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 0.000 412.990 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.070 0.000 420.350 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 0.000 282.350 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.430 0.000 427.710 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 0.000 435.070 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.150 0.000 442.430 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 0.000 449.790 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.410 0.000 456.690 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.130 0.000 471.410 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.490 0.000 478.770 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 0.000 486.130 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 292.010 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.110 0.000 500.390 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.470 0.000 507.750 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 0.000 301.670 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 0.000 311.330 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 0.000 318.690 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 0.000 326.050 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.130 0.000 333.410 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 0.000 340.310 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 0.000 265.330 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 0.000 274.990 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 0.000 357.330 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 0.000 364.690 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.770 0.000 372.050 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 0.000 379.410 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 0.000 393.670 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.750 0.000 401.030 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 0.000 408.390 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 0.000 415.750 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.830 0.000 423.110 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.730 0.000 430.010 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 0.000 437.370 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 0.000 444.730 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.810 0.000 452.090 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.170 0.000 459.450 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.070 0.000 466.350 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 0.000 473.710 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.790 0.000 481.070 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.150 0.000 488.430 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 0.000 495.790 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 0.000 294.310 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 0.000 510.050 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 0.000 303.970 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 0.000 313.630 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.710 0.000 320.990 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.070 0.000 328.350 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 0.000 335.710 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 0.000 343.070 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 0.000 349.970 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 0.000 360.090 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 0.000 366.990 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.070 0.000 374.350 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.430 0.000 381.710 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 0.000 389.070 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.050 0.000 403.330 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 0.000 410.690 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.770 0.000 418.050 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 0.000 432.770 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 0.000 439.670 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.750 0.000 447.030 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 0.000 461.750 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.830 0.000 469.110 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.190 0.000 476.470 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.450 0.000 490.730 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.810 0.000 498.090 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.170 0.000 505.450 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.530 0.000 512.810 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 0.000 306.730 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 0.000 316.390 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 0.000 323.290 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 0.000 330.650 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 0.000 338.010 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 0.000 345.370 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 0.000 352.730 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 0.000 289.710 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 0.000 299.370 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 0.000 309.030 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 585.580 590.325 ;
      LAYER met1 ;
        RECT 3.290 3.440 590.110 590.480 ;
      LAYER met2 ;
        RECT 1.010 597.920 6.710 598.810 ;
        RECT 7.550 597.920 20.970 598.810 ;
        RECT 21.810 597.920 35.230 598.810 ;
        RECT 36.070 597.920 49.950 598.810 ;
        RECT 50.790 597.920 64.210 598.810 ;
        RECT 65.050 597.920 78.470 598.810 ;
        RECT 79.310 597.920 93.190 598.810 ;
        RECT 94.030 597.920 107.450 598.810 ;
        RECT 108.290 597.920 121.710 598.810 ;
        RECT 122.550 597.920 136.430 598.810 ;
        RECT 137.270 597.920 150.690 598.810 ;
        RECT 151.530 597.920 165.410 598.810 ;
        RECT 166.250 597.920 179.670 598.810 ;
        RECT 180.510 597.920 193.930 598.810 ;
        RECT 194.770 597.920 208.650 598.810 ;
        RECT 209.490 597.920 222.910 598.810 ;
        RECT 223.750 597.920 237.170 598.810 ;
        RECT 238.010 597.920 251.890 598.810 ;
        RECT 252.730 597.920 266.150 598.810 ;
        RECT 266.990 597.920 280.410 598.810 ;
        RECT 281.250 597.920 295.130 598.810 ;
        RECT 295.970 597.920 309.390 598.810 ;
        RECT 310.230 597.920 324.110 598.810 ;
        RECT 324.950 597.920 338.370 598.810 ;
        RECT 339.210 597.920 352.630 598.810 ;
        RECT 353.470 597.920 367.350 598.810 ;
        RECT 368.190 597.920 381.610 598.810 ;
        RECT 382.450 597.920 395.870 598.810 ;
        RECT 396.710 597.920 410.590 598.810 ;
        RECT 411.430 597.920 424.850 598.810 ;
        RECT 425.690 597.920 439.110 598.810 ;
        RECT 439.950 597.920 453.830 598.810 ;
        RECT 454.670 597.920 468.090 598.810 ;
        RECT 468.930 597.920 482.810 598.810 ;
        RECT 483.650 597.920 497.070 598.810 ;
        RECT 497.910 597.920 511.330 598.810 ;
        RECT 512.170 597.920 526.050 598.810 ;
        RECT 526.890 597.920 540.310 598.810 ;
        RECT 541.150 597.920 554.570 598.810 ;
        RECT 555.410 597.920 569.290 598.810 ;
        RECT 570.130 597.920 583.550 598.810 ;
        RECT 584.390 597.920 590.080 598.810 ;
        RECT 1.010 4.280 590.080 597.920 ;
        RECT 1.570 3.410 3.030 4.280 ;
        RECT 3.870 3.410 5.330 4.280 ;
        RECT 6.170 3.410 7.630 4.280 ;
        RECT 8.470 3.410 10.390 4.280 ;
        RECT 11.230 3.410 12.690 4.280 ;
        RECT 13.530 3.410 14.990 4.280 ;
        RECT 15.830 3.410 17.290 4.280 ;
        RECT 18.130 3.410 20.050 4.280 ;
        RECT 20.890 3.410 22.350 4.280 ;
        RECT 23.190 3.410 24.650 4.280 ;
        RECT 25.490 3.410 26.950 4.280 ;
        RECT 27.790 3.410 29.710 4.280 ;
        RECT 30.550 3.410 32.010 4.280 ;
        RECT 32.850 3.410 34.310 4.280 ;
        RECT 35.150 3.410 37.070 4.280 ;
        RECT 37.910 3.410 39.370 4.280 ;
        RECT 40.210 3.410 41.670 4.280 ;
        RECT 42.510 3.410 43.970 4.280 ;
        RECT 44.810 3.410 46.730 4.280 ;
        RECT 47.570 3.410 49.030 4.280 ;
        RECT 49.870 3.410 51.330 4.280 ;
        RECT 52.170 3.410 53.630 4.280 ;
        RECT 54.470 3.410 56.390 4.280 ;
        RECT 57.230 3.410 58.690 4.280 ;
        RECT 59.530 3.410 60.990 4.280 ;
        RECT 61.830 3.410 63.750 4.280 ;
        RECT 64.590 3.410 66.050 4.280 ;
        RECT 66.890 3.410 68.350 4.280 ;
        RECT 69.190 3.410 70.650 4.280 ;
        RECT 71.490 3.410 73.410 4.280 ;
        RECT 74.250 3.410 75.710 4.280 ;
        RECT 76.550 3.410 78.010 4.280 ;
        RECT 78.850 3.410 80.310 4.280 ;
        RECT 81.150 3.410 83.070 4.280 ;
        RECT 83.910 3.410 85.370 4.280 ;
        RECT 86.210 3.410 87.670 4.280 ;
        RECT 88.510 3.410 90.430 4.280 ;
        RECT 91.270 3.410 92.730 4.280 ;
        RECT 93.570 3.410 95.030 4.280 ;
        RECT 95.870 3.410 97.330 4.280 ;
        RECT 98.170 3.410 100.090 4.280 ;
        RECT 100.930 3.410 102.390 4.280 ;
        RECT 103.230 3.410 104.690 4.280 ;
        RECT 105.530 3.410 106.990 4.280 ;
        RECT 107.830 3.410 109.750 4.280 ;
        RECT 110.590 3.410 112.050 4.280 ;
        RECT 112.890 3.410 114.350 4.280 ;
        RECT 115.190 3.410 116.650 4.280 ;
        RECT 117.490 3.410 119.410 4.280 ;
        RECT 120.250 3.410 121.710 4.280 ;
        RECT 122.550 3.410 124.010 4.280 ;
        RECT 124.850 3.410 126.770 4.280 ;
        RECT 127.610 3.410 129.070 4.280 ;
        RECT 129.910 3.410 131.370 4.280 ;
        RECT 132.210 3.410 133.670 4.280 ;
        RECT 134.510 3.410 136.430 4.280 ;
        RECT 137.270 3.410 138.730 4.280 ;
        RECT 139.570 3.410 141.030 4.280 ;
        RECT 141.870 3.410 143.330 4.280 ;
        RECT 144.170 3.410 146.090 4.280 ;
        RECT 146.930 3.410 148.390 4.280 ;
        RECT 149.230 3.410 150.690 4.280 ;
        RECT 151.530 3.410 153.450 4.280 ;
        RECT 154.290 3.410 155.750 4.280 ;
        RECT 156.590 3.410 158.050 4.280 ;
        RECT 158.890 3.410 160.350 4.280 ;
        RECT 161.190 3.410 163.110 4.280 ;
        RECT 163.950 3.410 165.410 4.280 ;
        RECT 166.250 3.410 167.710 4.280 ;
        RECT 168.550 3.410 170.010 4.280 ;
        RECT 170.850 3.410 172.770 4.280 ;
        RECT 173.610 3.410 175.070 4.280 ;
        RECT 175.910 3.410 177.370 4.280 ;
        RECT 178.210 3.410 180.130 4.280 ;
        RECT 180.970 3.410 182.430 4.280 ;
        RECT 183.270 3.410 184.730 4.280 ;
        RECT 185.570 3.410 187.030 4.280 ;
        RECT 187.870 3.410 189.790 4.280 ;
        RECT 190.630 3.410 192.090 4.280 ;
        RECT 192.930 3.410 194.390 4.280 ;
        RECT 195.230 3.410 196.690 4.280 ;
        RECT 197.530 3.410 199.450 4.280 ;
        RECT 200.290 3.410 201.750 4.280 ;
        RECT 202.590 3.410 204.050 4.280 ;
        RECT 204.890 3.410 206.350 4.280 ;
        RECT 207.190 3.410 209.110 4.280 ;
        RECT 209.950 3.410 211.410 4.280 ;
        RECT 212.250 3.410 213.710 4.280 ;
        RECT 214.550 3.410 216.470 4.280 ;
        RECT 217.310 3.410 218.770 4.280 ;
        RECT 219.610 3.410 221.070 4.280 ;
        RECT 221.910 3.410 223.370 4.280 ;
        RECT 224.210 3.410 226.130 4.280 ;
        RECT 226.970 3.410 228.430 4.280 ;
        RECT 229.270 3.410 230.730 4.280 ;
        RECT 231.570 3.410 233.030 4.280 ;
        RECT 233.870 3.410 235.790 4.280 ;
        RECT 236.630 3.410 238.090 4.280 ;
        RECT 238.930 3.410 240.390 4.280 ;
        RECT 241.230 3.410 243.150 4.280 ;
        RECT 243.990 3.410 245.450 4.280 ;
        RECT 246.290 3.410 247.750 4.280 ;
        RECT 248.590 3.410 250.050 4.280 ;
        RECT 250.890 3.410 252.810 4.280 ;
        RECT 253.650 3.410 255.110 4.280 ;
        RECT 255.950 3.410 257.410 4.280 ;
        RECT 258.250 3.410 259.710 4.280 ;
        RECT 260.550 3.410 262.470 4.280 ;
        RECT 263.310 3.410 264.770 4.280 ;
        RECT 265.610 3.410 267.070 4.280 ;
        RECT 267.910 3.410 269.830 4.280 ;
        RECT 270.670 3.410 272.130 4.280 ;
        RECT 272.970 3.410 274.430 4.280 ;
        RECT 275.270 3.410 276.730 4.280 ;
        RECT 277.570 3.410 279.490 4.280 ;
        RECT 280.330 3.410 281.790 4.280 ;
        RECT 282.630 3.410 284.090 4.280 ;
        RECT 284.930 3.410 286.390 4.280 ;
        RECT 287.230 3.410 289.150 4.280 ;
        RECT 289.990 3.410 291.450 4.280 ;
        RECT 292.290 3.410 293.750 4.280 ;
        RECT 294.590 3.410 296.510 4.280 ;
        RECT 297.350 3.410 298.810 4.280 ;
        RECT 299.650 3.410 301.110 4.280 ;
        RECT 301.950 3.410 303.410 4.280 ;
        RECT 304.250 3.410 306.170 4.280 ;
        RECT 307.010 3.410 308.470 4.280 ;
        RECT 309.310 3.410 310.770 4.280 ;
        RECT 311.610 3.410 313.070 4.280 ;
        RECT 313.910 3.410 315.830 4.280 ;
        RECT 316.670 3.410 318.130 4.280 ;
        RECT 318.970 3.410 320.430 4.280 ;
        RECT 321.270 3.410 322.730 4.280 ;
        RECT 323.570 3.410 325.490 4.280 ;
        RECT 326.330 3.410 327.790 4.280 ;
        RECT 328.630 3.410 330.090 4.280 ;
        RECT 330.930 3.410 332.850 4.280 ;
        RECT 333.690 3.410 335.150 4.280 ;
        RECT 335.990 3.410 337.450 4.280 ;
        RECT 338.290 3.410 339.750 4.280 ;
        RECT 340.590 3.410 342.510 4.280 ;
        RECT 343.350 3.410 344.810 4.280 ;
        RECT 345.650 3.410 347.110 4.280 ;
        RECT 347.950 3.410 349.410 4.280 ;
        RECT 350.250 3.410 352.170 4.280 ;
        RECT 353.010 3.410 354.470 4.280 ;
        RECT 355.310 3.410 356.770 4.280 ;
        RECT 357.610 3.410 359.530 4.280 ;
        RECT 360.370 3.410 361.830 4.280 ;
        RECT 362.670 3.410 364.130 4.280 ;
        RECT 364.970 3.410 366.430 4.280 ;
        RECT 367.270 3.410 369.190 4.280 ;
        RECT 370.030 3.410 371.490 4.280 ;
        RECT 372.330 3.410 373.790 4.280 ;
        RECT 374.630 3.410 376.090 4.280 ;
        RECT 376.930 3.410 378.850 4.280 ;
        RECT 379.690 3.410 381.150 4.280 ;
        RECT 381.990 3.410 383.450 4.280 ;
        RECT 384.290 3.410 386.210 4.280 ;
        RECT 387.050 3.410 388.510 4.280 ;
        RECT 389.350 3.410 390.810 4.280 ;
        RECT 391.650 3.410 393.110 4.280 ;
        RECT 393.950 3.410 395.870 4.280 ;
        RECT 396.710 3.410 398.170 4.280 ;
        RECT 399.010 3.410 400.470 4.280 ;
        RECT 401.310 3.410 402.770 4.280 ;
        RECT 403.610 3.410 405.530 4.280 ;
        RECT 406.370 3.410 407.830 4.280 ;
        RECT 408.670 3.410 410.130 4.280 ;
        RECT 410.970 3.410 412.430 4.280 ;
        RECT 413.270 3.410 415.190 4.280 ;
        RECT 416.030 3.410 417.490 4.280 ;
        RECT 418.330 3.410 419.790 4.280 ;
        RECT 420.630 3.410 422.550 4.280 ;
        RECT 423.390 3.410 424.850 4.280 ;
        RECT 425.690 3.410 427.150 4.280 ;
        RECT 427.990 3.410 429.450 4.280 ;
        RECT 430.290 3.410 432.210 4.280 ;
        RECT 433.050 3.410 434.510 4.280 ;
        RECT 435.350 3.410 436.810 4.280 ;
        RECT 437.650 3.410 439.110 4.280 ;
        RECT 439.950 3.410 441.870 4.280 ;
        RECT 442.710 3.410 444.170 4.280 ;
        RECT 445.010 3.410 446.470 4.280 ;
        RECT 447.310 3.410 449.230 4.280 ;
        RECT 450.070 3.410 451.530 4.280 ;
        RECT 452.370 3.410 453.830 4.280 ;
        RECT 454.670 3.410 456.130 4.280 ;
        RECT 456.970 3.410 458.890 4.280 ;
        RECT 459.730 3.410 461.190 4.280 ;
        RECT 462.030 3.410 463.490 4.280 ;
        RECT 464.330 3.410 465.790 4.280 ;
        RECT 466.630 3.410 468.550 4.280 ;
        RECT 469.390 3.410 470.850 4.280 ;
        RECT 471.690 3.410 473.150 4.280 ;
        RECT 473.990 3.410 475.910 4.280 ;
        RECT 476.750 3.410 478.210 4.280 ;
        RECT 479.050 3.410 480.510 4.280 ;
        RECT 481.350 3.410 482.810 4.280 ;
        RECT 483.650 3.410 485.570 4.280 ;
        RECT 486.410 3.410 487.870 4.280 ;
        RECT 488.710 3.410 490.170 4.280 ;
        RECT 491.010 3.410 492.470 4.280 ;
        RECT 493.310 3.410 495.230 4.280 ;
        RECT 496.070 3.410 497.530 4.280 ;
        RECT 498.370 3.410 499.830 4.280 ;
        RECT 500.670 3.410 502.130 4.280 ;
        RECT 502.970 3.410 504.890 4.280 ;
        RECT 505.730 3.410 507.190 4.280 ;
        RECT 508.030 3.410 509.490 4.280 ;
        RECT 510.330 3.410 512.250 4.280 ;
        RECT 513.090 3.410 514.550 4.280 ;
        RECT 515.390 3.410 516.850 4.280 ;
        RECT 517.690 3.410 519.150 4.280 ;
        RECT 519.990 3.410 521.910 4.280 ;
        RECT 522.750 3.410 524.210 4.280 ;
        RECT 525.050 3.410 526.510 4.280 ;
        RECT 527.350 3.410 528.810 4.280 ;
        RECT 529.650 3.410 531.570 4.280 ;
        RECT 532.410 3.410 533.870 4.280 ;
        RECT 534.710 3.410 536.170 4.280 ;
        RECT 537.010 3.410 538.930 4.280 ;
        RECT 539.770 3.410 541.230 4.280 ;
        RECT 542.070 3.410 543.530 4.280 ;
        RECT 544.370 3.410 545.830 4.280 ;
        RECT 546.670 3.410 548.590 4.280 ;
        RECT 549.430 3.410 550.890 4.280 ;
        RECT 551.730 3.410 553.190 4.280 ;
        RECT 554.030 3.410 555.490 4.280 ;
        RECT 556.330 3.410 558.250 4.280 ;
        RECT 559.090 3.410 560.550 4.280 ;
        RECT 561.390 3.410 562.850 4.280 ;
        RECT 563.690 3.410 565.610 4.280 ;
        RECT 566.450 3.410 567.910 4.280 ;
        RECT 568.750 3.410 570.210 4.280 ;
        RECT 571.050 3.410 572.510 4.280 ;
        RECT 573.350 3.410 575.270 4.280 ;
        RECT 576.110 3.410 577.570 4.280 ;
        RECT 578.410 3.410 579.870 4.280 ;
        RECT 580.710 3.410 582.170 4.280 ;
        RECT 583.010 3.410 584.930 4.280 ;
        RECT 585.770 3.410 587.230 4.280 ;
        RECT 588.070 3.410 589.530 4.280 ;
      LAYER met3 ;
        RECT 0.985 594.640 587.080 595.505 ;
        RECT 0.985 593.320 587.480 594.640 ;
        RECT 4.400 591.920 587.480 593.320 ;
        RECT 0.985 582.440 587.480 591.920 ;
        RECT 0.985 581.040 587.080 582.440 ;
        RECT 0.985 573.600 587.480 581.040 ;
        RECT 4.400 572.200 587.480 573.600 ;
        RECT 0.985 568.840 587.480 572.200 ;
        RECT 0.985 567.440 587.080 568.840 ;
        RECT 0.985 555.240 587.480 567.440 ;
        RECT 0.985 554.560 587.080 555.240 ;
        RECT 4.400 553.840 587.080 554.560 ;
        RECT 4.400 553.160 587.480 553.840 ;
        RECT 0.985 541.640 587.480 553.160 ;
        RECT 0.985 540.240 587.080 541.640 ;
        RECT 0.985 534.840 587.480 540.240 ;
        RECT 4.400 533.440 587.480 534.840 ;
        RECT 0.985 528.040 587.480 533.440 ;
        RECT 0.985 526.640 587.080 528.040 ;
        RECT 0.985 515.800 587.480 526.640 ;
        RECT 4.400 514.440 587.480 515.800 ;
        RECT 4.400 514.400 587.080 514.440 ;
        RECT 0.985 513.040 587.080 514.400 ;
        RECT 0.985 500.160 587.480 513.040 ;
        RECT 0.985 498.760 587.080 500.160 ;
        RECT 0.985 496.080 587.480 498.760 ;
        RECT 4.400 494.680 587.480 496.080 ;
        RECT 0.985 486.560 587.480 494.680 ;
        RECT 0.985 485.160 587.080 486.560 ;
        RECT 0.985 476.360 587.480 485.160 ;
        RECT 4.400 474.960 587.480 476.360 ;
        RECT 0.985 472.960 587.480 474.960 ;
        RECT 0.985 471.560 587.080 472.960 ;
        RECT 0.985 459.360 587.480 471.560 ;
        RECT 0.985 457.960 587.080 459.360 ;
        RECT 0.985 457.320 587.480 457.960 ;
        RECT 4.400 455.920 587.480 457.320 ;
        RECT 0.985 445.760 587.480 455.920 ;
        RECT 0.985 444.360 587.080 445.760 ;
        RECT 0.985 437.600 587.480 444.360 ;
        RECT 4.400 436.200 587.480 437.600 ;
        RECT 0.985 432.160 587.480 436.200 ;
        RECT 0.985 430.760 587.080 432.160 ;
        RECT 0.985 418.560 587.480 430.760 ;
        RECT 4.400 417.160 587.080 418.560 ;
        RECT 0.985 404.280 587.480 417.160 ;
        RECT 0.985 402.880 587.080 404.280 ;
        RECT 0.985 398.840 587.480 402.880 ;
        RECT 4.400 397.440 587.480 398.840 ;
        RECT 0.985 390.680 587.480 397.440 ;
        RECT 0.985 389.280 587.080 390.680 ;
        RECT 0.985 379.800 587.480 389.280 ;
        RECT 4.400 378.400 587.480 379.800 ;
        RECT 0.985 377.080 587.480 378.400 ;
        RECT 0.985 375.680 587.080 377.080 ;
        RECT 0.985 363.480 587.480 375.680 ;
        RECT 0.985 362.080 587.080 363.480 ;
        RECT 0.985 360.080 587.480 362.080 ;
        RECT 4.400 358.680 587.480 360.080 ;
        RECT 0.985 349.880 587.480 358.680 ;
        RECT 0.985 348.480 587.080 349.880 ;
        RECT 0.985 340.360 587.480 348.480 ;
        RECT 4.400 338.960 587.480 340.360 ;
        RECT 0.985 336.280 587.480 338.960 ;
        RECT 0.985 334.880 587.080 336.280 ;
        RECT 0.985 322.680 587.480 334.880 ;
        RECT 0.985 321.320 587.080 322.680 ;
        RECT 4.400 321.280 587.080 321.320 ;
        RECT 4.400 319.920 587.480 321.280 ;
        RECT 0.985 309.080 587.480 319.920 ;
        RECT 0.985 307.680 587.080 309.080 ;
        RECT 0.985 301.600 587.480 307.680 ;
        RECT 4.400 300.200 587.480 301.600 ;
        RECT 0.985 294.800 587.480 300.200 ;
        RECT 0.985 293.400 587.080 294.800 ;
        RECT 0.985 282.560 587.480 293.400 ;
        RECT 4.400 281.200 587.480 282.560 ;
        RECT 4.400 281.160 587.080 281.200 ;
        RECT 0.985 279.800 587.080 281.160 ;
        RECT 0.985 267.600 587.480 279.800 ;
        RECT 0.985 266.200 587.080 267.600 ;
        RECT 0.985 262.840 587.480 266.200 ;
        RECT 4.400 261.440 587.480 262.840 ;
        RECT 0.985 254.000 587.480 261.440 ;
        RECT 0.985 252.600 587.080 254.000 ;
        RECT 0.985 243.120 587.480 252.600 ;
        RECT 4.400 241.720 587.480 243.120 ;
        RECT 0.985 240.400 587.480 241.720 ;
        RECT 0.985 239.000 587.080 240.400 ;
        RECT 0.985 226.800 587.480 239.000 ;
        RECT 0.985 225.400 587.080 226.800 ;
        RECT 0.985 224.080 587.480 225.400 ;
        RECT 4.400 222.680 587.480 224.080 ;
        RECT 0.985 213.200 587.480 222.680 ;
        RECT 0.985 211.800 587.080 213.200 ;
        RECT 0.985 204.360 587.480 211.800 ;
        RECT 4.400 202.960 587.480 204.360 ;
        RECT 0.985 198.920 587.480 202.960 ;
        RECT 0.985 197.520 587.080 198.920 ;
        RECT 0.985 185.320 587.480 197.520 ;
        RECT 4.400 183.920 587.080 185.320 ;
        RECT 0.985 171.720 587.480 183.920 ;
        RECT 0.985 170.320 587.080 171.720 ;
        RECT 0.985 165.600 587.480 170.320 ;
        RECT 4.400 164.200 587.480 165.600 ;
        RECT 0.985 158.120 587.480 164.200 ;
        RECT 0.985 156.720 587.080 158.120 ;
        RECT 0.985 146.560 587.480 156.720 ;
        RECT 4.400 145.160 587.480 146.560 ;
        RECT 0.985 144.520 587.480 145.160 ;
        RECT 0.985 143.120 587.080 144.520 ;
        RECT 0.985 130.920 587.480 143.120 ;
        RECT 0.985 129.520 587.080 130.920 ;
        RECT 0.985 126.840 587.480 129.520 ;
        RECT 4.400 125.440 587.480 126.840 ;
        RECT 0.985 117.320 587.480 125.440 ;
        RECT 0.985 115.920 587.080 117.320 ;
        RECT 0.985 107.120 587.480 115.920 ;
        RECT 4.400 105.720 587.480 107.120 ;
        RECT 0.985 103.040 587.480 105.720 ;
        RECT 0.985 101.640 587.080 103.040 ;
        RECT 0.985 89.440 587.480 101.640 ;
        RECT 0.985 88.080 587.080 89.440 ;
        RECT 4.400 88.040 587.080 88.080 ;
        RECT 4.400 86.680 587.480 88.040 ;
        RECT 0.985 75.840 587.480 86.680 ;
        RECT 0.985 74.440 587.080 75.840 ;
        RECT 0.985 68.360 587.480 74.440 ;
        RECT 4.400 66.960 587.480 68.360 ;
        RECT 0.985 62.240 587.480 66.960 ;
        RECT 0.985 60.840 587.080 62.240 ;
        RECT 0.985 49.320 587.480 60.840 ;
        RECT 4.400 48.640 587.480 49.320 ;
        RECT 4.400 47.920 587.080 48.640 ;
        RECT 0.985 47.240 587.080 47.920 ;
        RECT 0.985 35.040 587.480 47.240 ;
        RECT 0.985 33.640 587.080 35.040 ;
        RECT 0.985 29.600 587.480 33.640 ;
        RECT 4.400 28.200 587.480 29.600 ;
        RECT 0.985 21.440 587.480 28.200 ;
        RECT 0.985 20.040 587.080 21.440 ;
        RECT 0.985 10.560 587.480 20.040 ;
        RECT 4.400 9.160 587.480 10.560 ;
        RECT 0.985 7.840 587.480 9.160 ;
        RECT 0.985 6.975 587.080 7.840 ;
      LAYER met4 ;
        RECT 3.055 590.880 569.185 591.425 ;
        RECT 3.055 10.240 20.640 590.880 ;
        RECT 23.040 10.240 97.440 590.880 ;
        RECT 99.840 10.240 174.240 590.880 ;
        RECT 176.640 10.240 251.040 590.880 ;
        RECT 253.440 10.240 327.840 590.880 ;
        RECT 330.240 10.240 404.640 590.880 ;
        RECT 407.040 10.240 481.440 590.880 ;
        RECT 483.840 10.240 558.240 590.880 ;
        RECT 560.640 10.240 569.185 590.880 ;
        RECT 3.055 9.695 569.185 10.240 ;
  END
END rvj1_caravel_soc
END LIBRARY

