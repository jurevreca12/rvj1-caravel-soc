magic
tech sky130A
magscale 1 2
timestamp 1653944755
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 219342 700408 219348 700460
rect 219400 700448 219406 700460
rect 267642 700448 267648 700460
rect 219400 700420 267648 700448
rect 219400 700408 219406 700420
rect 267642 700408 267648 700420
rect 267700 700408 267706 700460
rect 137830 700340 137836 700392
rect 137888 700380 137894 700392
rect 138658 700380 138664 700392
rect 137888 700352 138664 700380
rect 137888 700340 137894 700352
rect 138658 700340 138664 700352
rect 138716 700340 138722 700392
rect 217962 700340 217968 700392
rect 218020 700380 218026 700392
rect 283834 700380 283840 700392
rect 218020 700352 283840 700380
rect 218020 700340 218026 700352
rect 283834 700340 283840 700352
rect 283892 700340 283898 700392
rect 348786 700340 348792 700392
rect 348844 700380 348850 700392
rect 358814 700380 358820 700392
rect 348844 700352 358820 700380
rect 348844 700340 348850 700352
rect 358814 700340 358820 700352
rect 358872 700340 358878 700392
rect 24302 700272 24308 700324
rect 24360 700312 24366 700324
rect 215938 700312 215944 700324
rect 24360 700284 215944 700312
rect 24360 700272 24366 700284
rect 215938 700272 215944 700284
rect 215996 700272 216002 700324
rect 217870 700272 217876 700324
rect 217928 700312 217934 700324
rect 300118 700312 300124 700324
rect 217928 700284 300124 700312
rect 217928 700272 217934 700284
rect 300118 700272 300124 700284
rect 300176 700272 300182 700324
rect 332502 700272 332508 700324
rect 332560 700312 332566 700324
rect 357434 700312 357440 700324
rect 332560 700284 357440 700312
rect 332560 700272 332566 700284
rect 357434 700272 357440 700284
rect 357492 700272 357498 700324
rect 359458 700272 359464 700324
rect 359516 700312 359522 700324
rect 429838 700312 429844 700324
rect 359516 700284 429844 700312
rect 359516 700272 359522 700284
rect 429838 700272 429844 700284
rect 429896 700272 429902 700324
rect 442258 700272 442264 700324
rect 442316 700312 442322 700324
rect 559650 700312 559656 700324
rect 442316 700284 559656 700312
rect 442316 700272 442322 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 105446 699728 105452 699780
rect 105504 699768 105510 699780
rect 108298 699768 108304 699780
rect 105504 699740 108304 699768
rect 105504 699728 105510 699740
rect 108298 699728 108304 699740
rect 108356 699728 108362 699780
rect 8110 699660 8116 699712
rect 8168 699700 8174 699712
rect 10318 699700 10324 699712
rect 8168 699672 10324 699700
rect 8168 699660 8174 699672
rect 10318 699660 10324 699672
rect 10376 699660 10382 699712
rect 396718 699660 396724 699712
rect 396776 699700 396782 699712
rect 397454 699700 397460 699712
rect 396776 699672 397460 699700
rect 396776 699660 396782 699672
rect 397454 699660 397460 699672
rect 397512 699660 397518 699712
rect 391198 696940 391204 696992
rect 391256 696980 391262 696992
rect 580166 696980 580172 696992
rect 391256 696952 580172 696980
rect 391256 696940 391262 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 21358 683176 21364 683188
rect 3476 683148 21364 683176
rect 3476 683136 3482 683148
rect 21358 683136 21364 683148
rect 21416 683136 21422 683188
rect 378778 683136 378784 683188
rect 378836 683176 378842 683188
rect 580166 683176 580172 683188
rect 378836 683148 580172 683176
rect 378836 683136 378842 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 214558 670732 214564 670744
rect 3568 670704 214564 670732
rect 3568 670692 3574 670704
rect 214558 670692 214564 670704
rect 214616 670692 214622 670744
rect 377398 670692 377404 670744
rect 377456 670732 377462 670744
rect 580166 670732 580172 670744
rect 377456 670704 580172 670732
rect 377456 670692 377462 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 28258 656928 28264 656940
rect 3476 656900 28264 656928
rect 3476 656888 3482 656900
rect 28258 656888 28264 656900
rect 28316 656888 28322 656940
rect 373258 643084 373264 643136
rect 373316 643124 373322 643136
rect 580166 643124 580172 643136
rect 373316 643096 580172 643124
rect 373316 643084 373322 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 2774 632068 2780 632120
rect 2832 632108 2838 632120
rect 4798 632108 4804 632120
rect 2832 632080 4804 632108
rect 2832 632068 2838 632080
rect 4798 632068 4804 632080
rect 4856 632068 4862 632120
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 211798 618304 211804 618316
rect 3200 618276 211804 618304
rect 3200 618264 3206 618276
rect 211798 618264 211804 618276
rect 211856 618264 211862 618316
rect 363598 616836 363604 616888
rect 363656 616876 363662 616888
rect 580166 616876 580172 616888
rect 363656 616848 580172 616876
rect 363656 616836 363662 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3418 606024 3424 606076
rect 3476 606064 3482 606076
rect 7558 606064 7564 606076
rect 3476 606036 7564 606064
rect 3476 606024 3482 606036
rect 7558 606024 7564 606036
rect 7616 606024 7622 606076
rect 374638 590656 374644 590708
rect 374696 590696 374702 590708
rect 580166 590696 580172 590708
rect 374696 590668 580172 590696
rect 374696 590656 374702 590668
rect 580166 590656 580172 590668
rect 580224 590656 580230 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 57238 579680 57244 579692
rect 3384 579652 57244 579680
rect 3384 579640 3390 579652
rect 57238 579640 57244 579652
rect 57296 579640 57302 579692
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 210418 565876 210424 565888
rect 3476 565848 210424 565876
rect 3476 565836 3482 565848
rect 210418 565836 210424 565848
rect 210476 565836 210482 565888
rect 217778 565088 217784 565140
rect 217836 565128 217842 565140
rect 234614 565128 234620 565140
rect 217836 565100 234620 565128
rect 217836 565088 217842 565100
rect 234614 565088 234620 565100
rect 234672 565088 234678 565140
rect 360838 563048 360844 563100
rect 360896 563088 360902 563100
rect 579890 563088 579896 563100
rect 360896 563060 579896 563088
rect 360896 563048 360902 563060
rect 579890 563048 579896 563060
rect 579948 563048 579954 563100
rect 3418 553664 3424 553716
rect 3476 553704 3482 553716
rect 8938 553704 8944 553716
rect 3476 553676 8944 553704
rect 3476 553664 3482 553676
rect 8938 553664 8944 553676
rect 8996 553664 9002 553716
rect 369118 536800 369124 536852
rect 369176 536840 369182 536852
rect 580166 536840 580172 536852
rect 369176 536812 580172 536840
rect 369176 536800 369182 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 3418 527144 3424 527196
rect 3476 527184 3482 527196
rect 35158 527184 35164 527196
rect 3476 527156 35164 527184
rect 3476 527144 3482 527156
rect 35158 527144 35164 527156
rect 35216 527144 35222 527196
rect 371878 524424 371884 524476
rect 371936 524464 371942 524476
rect 580166 524464 580172 524476
rect 371936 524436 580172 524464
rect 371936 524424 371942 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3418 514768 3424 514820
rect 3476 514808 3482 514820
rect 207658 514808 207664 514820
rect 3476 514780 207664 514808
rect 3476 514768 3482 514780
rect 207658 514768 207664 514780
rect 207716 514768 207722 514820
rect 358078 510620 358084 510672
rect 358136 510660 358142 510672
rect 580166 510660 580172 510672
rect 358136 510632 580172 510660
rect 358136 510620 358142 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 13078 501004 13084 501016
rect 3108 500976 13084 501004
rect 3108 500964 3114 500976
rect 13078 500964 13084 500976
rect 13136 500964 13142 501016
rect 367738 484372 367744 484424
rect 367796 484412 367802 484424
rect 580166 484412 580172 484424
rect 367796 484384 580172 484412
rect 367796 484372 367802 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 217870 478592 217876 478644
rect 217928 478632 217934 478644
rect 269942 478632 269948 478644
rect 217928 478604 269948 478632
rect 217928 478592 217934 478604
rect 269942 478592 269948 478604
rect 270000 478592 270006 478644
rect 217962 478524 217968 478576
rect 218020 478564 218026 478576
rect 271230 478564 271236 478576
rect 218020 478536 271236 478564
rect 218020 478524 218026 478536
rect 271230 478524 271236 478536
rect 271288 478524 271294 478576
rect 268654 478456 268660 478508
rect 268712 478496 268718 478508
rect 357434 478496 357440 478508
rect 268712 478468 357440 478496
rect 268712 478456 268718 478468
rect 357434 478456 357440 478468
rect 357492 478456 357498 478508
rect 269298 478388 269304 478440
rect 269356 478428 269362 478440
rect 358814 478428 358820 478440
rect 269356 478400 358820 478428
rect 269356 478388 269362 478400
rect 358814 478388 358820 478400
rect 358872 478388 358878 478440
rect 217410 478320 217416 478372
rect 217468 478360 217474 478372
rect 308582 478360 308588 478372
rect 217468 478332 308588 478360
rect 217468 478320 217474 478332
rect 308582 478320 308588 478332
rect 308640 478320 308646 478372
rect 218974 478252 218980 478304
rect 219032 478292 219038 478304
rect 314470 478292 314476 478304
rect 219032 478264 314476 478292
rect 219032 478252 219038 478264
rect 314470 478252 314476 478264
rect 314528 478252 314534 478304
rect 256878 478184 256884 478236
rect 256936 478224 256942 478236
rect 374638 478224 374644 478236
rect 256936 478196 374644 478224
rect 256936 478184 256942 478196
rect 374638 478184 374644 478196
rect 374696 478184 374702 478236
rect 7558 478116 7564 478168
rect 7616 478156 7622 478168
rect 282362 478156 282368 478168
rect 7616 478128 282368 478156
rect 7616 478116 7622 478128
rect 282362 478116 282368 478128
rect 282420 478116 282426 478168
rect 241422 476824 241428 476876
rect 241480 476864 241486 476876
rect 241480 476836 248414 476864
rect 241480 476824 241486 476836
rect 238478 476756 238484 476808
rect 238536 476796 238542 476808
rect 248386 476796 248414 476836
rect 316402 476796 316408 476808
rect 238536 476768 243584 476796
rect 248386 476768 316408 476796
rect 238536 476756 238542 476768
rect 237282 476688 237288 476740
rect 237340 476728 237346 476740
rect 239398 476728 239404 476740
rect 237340 476700 239404 476728
rect 237340 476688 237346 476700
rect 239398 476688 239404 476700
rect 239456 476688 239462 476740
rect 243556 476728 243584 476768
rect 316402 476756 316408 476768
rect 316460 476756 316466 476808
rect 311250 476728 311256 476740
rect 243556 476700 311256 476728
rect 311250 476688 311256 476700
rect 311308 476688 311314 476740
rect 242802 476620 242808 476672
rect 242860 476660 242866 476672
rect 319070 476660 319076 476672
rect 242860 476632 319076 476660
rect 242860 476620 242866 476632
rect 319070 476620 319076 476632
rect 319128 476620 319134 476672
rect 271782 476552 271788 476604
rect 271840 476592 271846 476604
rect 330202 476592 330208 476604
rect 271840 476564 330208 476592
rect 271840 476552 271846 476564
rect 330202 476552 330208 476564
rect 330260 476552 330266 476604
rect 266262 476484 266268 476536
rect 266320 476524 266326 476536
rect 326890 476524 326896 476536
rect 266320 476496 326896 476524
rect 266320 476484 266326 476496
rect 326890 476484 326896 476496
rect 326948 476484 326954 476536
rect 256602 476416 256608 476468
rect 256660 476456 256666 476468
rect 318426 476456 318432 476468
rect 256660 476428 318432 476456
rect 256660 476416 256666 476428
rect 318426 476416 318432 476428
rect 318484 476416 318490 476468
rect 318702 476416 318708 476468
rect 318760 476456 318766 476468
rect 335998 476456 336004 476468
rect 318760 476428 336004 476456
rect 318760 476416 318766 476428
rect 335998 476416 336004 476428
rect 336056 476416 336062 476468
rect 262122 476348 262128 476400
rect 262180 476388 262186 476400
rect 323026 476388 323032 476400
rect 262180 476360 323032 476388
rect 262180 476348 262186 476360
rect 323026 476348 323032 476360
rect 323084 476348 323090 476400
rect 326982 476348 326988 476400
rect 327040 476388 327046 476400
rect 338758 476388 338764 476400
rect 327040 476360 338764 476388
rect 327040 476348 327046 476360
rect 338758 476348 338764 476360
rect 338816 476348 338822 476400
rect 309042 476280 309048 476332
rect 309100 476320 309106 476332
rect 329098 476320 329104 476332
rect 309100 476292 329104 476320
rect 309100 476280 309106 476292
rect 329098 476280 329104 476292
rect 329156 476280 329162 476332
rect 311802 476212 311808 476264
rect 311860 476252 311866 476264
rect 331858 476252 331864 476264
rect 311860 476224 331864 476252
rect 311860 476212 311866 476224
rect 331858 476212 331864 476224
rect 331916 476212 331922 476264
rect 315942 476144 315948 476196
rect 316000 476184 316006 476196
rect 334618 476184 334624 476196
rect 316000 476156 334624 476184
rect 316000 476144 316006 476156
rect 334618 476144 334624 476156
rect 334676 476144 334682 476196
rect 240042 476076 240048 476128
rect 240100 476116 240106 476128
rect 313826 476116 313832 476128
rect 240100 476088 313832 476116
rect 240100 476076 240106 476088
rect 313826 476076 313832 476088
rect 313884 476076 313890 476128
rect 314562 476076 314568 476128
rect 314620 476116 314626 476128
rect 333238 476116 333244 476128
rect 314620 476088 333244 476116
rect 314620 476076 314626 476088
rect 333238 476076 333244 476088
rect 333296 476076 333302 476128
rect 274542 475464 274548 475516
rect 274600 475504 274606 475516
rect 331490 475504 331496 475516
rect 274600 475476 331496 475504
rect 274600 475464 274606 475476
rect 331490 475464 331496 475476
rect 331548 475464 331554 475516
rect 219066 475396 219072 475448
rect 219124 475436 219130 475448
rect 321646 475436 321652 475448
rect 219124 475408 321652 475436
rect 219124 475396 219130 475408
rect 321646 475396 321652 475408
rect 321704 475396 321710 475448
rect 324222 475396 324228 475448
rect 324280 475436 324286 475448
rect 352558 475436 352564 475448
rect 324280 475408 352564 475436
rect 324280 475396 324286 475408
rect 352558 475396 352564 475408
rect 352616 475396 352622 475448
rect 255590 475328 255596 475380
rect 255648 475368 255654 475380
rect 371878 475368 371884 475380
rect 255648 475340 371884 475368
rect 255648 475328 255654 475340
rect 371878 475328 371884 475340
rect 371936 475328 371942 475380
rect 3418 474716 3424 474768
rect 3476 474756 3482 474768
rect 287606 474756 287612 474768
rect 3476 474728 287612 474756
rect 3476 474716 3482 474728
rect 287606 474716 287612 474728
rect 287664 474716 287670 474768
rect 253750 474172 253756 474224
rect 253808 474212 253814 474224
rect 329558 474212 329564 474224
rect 253808 474184 329564 474212
rect 253808 474172 253814 474184
rect 329558 474172 329564 474184
rect 329616 474172 329622 474224
rect 217502 474104 217508 474156
rect 217560 474144 217566 474156
rect 323670 474144 323676 474156
rect 217560 474116 323676 474144
rect 217560 474104 217566 474116
rect 323670 474104 323676 474116
rect 323728 474104 323734 474156
rect 254854 474036 254860 474088
rect 254912 474076 254918 474088
rect 369118 474076 369124 474088
rect 254912 474048 369124 474076
rect 254912 474036 254918 474048
rect 369118 474036 369124 474048
rect 369176 474036 369182 474088
rect 8938 473968 8944 474020
rect 8996 474008 9002 474020
rect 284386 474008 284392 474020
rect 8996 473980 284392 474008
rect 8996 473968 9002 473980
rect 284386 473968 284392 473980
rect 284444 473968 284450 474020
rect 321462 473968 321468 474020
rect 321520 474008 321526 474020
rect 356422 474008 356428 474020
rect 321520 473980 356428 474008
rect 321520 473968 321526 473980
rect 356422 473968 356428 473980
rect 356480 473968 356486 474020
rect 259270 472812 259276 472864
rect 259328 472852 259334 472864
rect 294598 472852 294604 472864
rect 259328 472824 294604 472852
rect 259328 472812 259334 472824
rect 294598 472812 294604 472824
rect 294656 472812 294662 472864
rect 219158 472744 219164 472796
rect 219216 472784 219222 472796
rect 319714 472784 319720 472796
rect 219216 472756 319720 472784
rect 219216 472744 219222 472756
rect 319714 472744 319720 472756
rect 319772 472744 319778 472796
rect 252922 472676 252928 472728
rect 252980 472716 252986 472728
rect 367738 472716 367744 472728
rect 252980 472688 367744 472716
rect 252980 472676 252986 472688
rect 367738 472676 367744 472688
rect 367796 472676 367802 472728
rect 153194 472608 153200 472660
rect 153252 472648 153258 472660
rect 275186 472648 275192 472660
rect 153252 472620 275192 472648
rect 153252 472608 153258 472620
rect 275186 472608 275192 472620
rect 275244 472608 275250 472660
rect 275922 472608 275928 472660
rect 275980 472648 275986 472660
rect 354398 472648 354404 472660
rect 275980 472620 354404 472648
rect 275980 472608 275986 472620
rect 354398 472608 354404 472620
rect 354456 472608 354462 472660
rect 264790 471384 264796 471436
rect 264848 471424 264854 471436
rect 295978 471424 295984 471436
rect 264848 471396 295984 471424
rect 264848 471384 264854 471396
rect 295978 471384 295984 471396
rect 296036 471384 296042 471436
rect 217594 471316 217600 471368
rect 217652 471356 217658 471368
rect 327534 471356 327540 471368
rect 217652 471328 327540 471356
rect 217652 471316 217658 471328
rect 327534 471316 327540 471328
rect 327592 471316 327598 471368
rect 13078 471248 13084 471300
rect 13136 471288 13142 471300
rect 286318 471288 286324 471300
rect 13136 471260 286324 471288
rect 13136 471248 13142 471260
rect 286318 471248 286324 471260
rect 286376 471248 286382 471300
rect 286502 471248 286508 471300
rect 286560 471288 286566 471300
rect 338022 471288 338028 471300
rect 286560 471260 338028 471288
rect 286560 471248 286566 471260
rect 338022 471248 338028 471260
rect 338080 471248 338086 471300
rect 253198 470568 253204 470620
rect 253256 470608 253262 470620
rect 580166 470608 580172 470620
rect 253256 470580 580172 470608
rect 253256 470568 253262 470580
rect 580166 470568 580172 470580
rect 580224 470568 580230 470620
rect 253842 470024 253848 470076
rect 253900 470064 253906 470076
rect 315758 470064 315764 470076
rect 253900 470036 315764 470064
rect 253900 470024 253906 470036
rect 315758 470024 315764 470036
rect 315816 470024 315822 470076
rect 255222 469956 255228 470008
rect 255280 469996 255286 470008
rect 330846 469996 330852 470008
rect 255280 469968 330852 469996
rect 255280 469956 255286 469968
rect 330846 469956 330852 469968
rect 330904 469956 330910 470008
rect 261478 469888 261484 469940
rect 261536 469928 261542 469940
rect 378778 469928 378784 469940
rect 261536 469900 378784 469928
rect 261536 469888 261542 469900
rect 378778 469888 378784 469900
rect 378836 469888 378842 469940
rect 35158 469820 35164 469872
rect 35216 469860 35222 469872
rect 285674 469860 285680 469872
rect 35216 469832 285680 469860
rect 35216 469820 35222 469832
rect 285674 469820 285680 469832
rect 285732 469820 285738 469872
rect 288342 469820 288348 469872
rect 288400 469860 288406 469872
rect 339402 469860 339408 469872
rect 288400 469832 339408 469860
rect 288400 469820 288406 469832
rect 339402 469820 339408 469832
rect 339460 469820 339466 469872
rect 248230 468664 248236 468716
rect 248288 468704 248294 468716
rect 320358 468704 320364 468716
rect 248288 468676 320364 468704
rect 248288 468664 248294 468676
rect 320358 468664 320364 468676
rect 320416 468664 320422 468716
rect 219250 468596 219256 468648
rect 219308 468636 219314 468648
rect 317138 468636 317144 468648
rect 219308 468608 317144 468636
rect 219308 468596 219314 468608
rect 317138 468596 317144 468608
rect 317196 468596 317202 468648
rect 264698 468528 264704 468580
rect 264756 468568 264762 468580
rect 462314 468568 462320 468580
rect 264756 468540 462320 468568
rect 264756 468528 264762 468540
rect 462314 468528 462320 468540
rect 462372 468528 462378 468580
rect 57238 468460 57244 468512
rect 57296 468500 57302 468512
rect 283742 468500 283748 468512
rect 57296 468472 283748 468500
rect 57296 468460 57302 468472
rect 283742 468460 283748 468472
rect 283800 468460 283806 468512
rect 296622 468460 296628 468512
rect 296680 468500 296686 468512
rect 343266 468500 343272 468512
rect 296680 468472 343272 468500
rect 296680 468460 296686 468472
rect 343266 468460 343272 468472
rect 343324 468460 343330 468512
rect 252370 467304 252376 467356
rect 252428 467344 252434 467356
rect 326246 467344 326252 467356
rect 252428 467316 326252 467344
rect 252428 467304 252434 467316
rect 326246 467304 326252 467316
rect 326304 467304 326310 467356
rect 217686 467236 217692 467288
rect 217744 467276 217750 467288
rect 325602 467276 325608 467288
rect 217744 467248 325608 467276
rect 217744 467236 217750 467248
rect 325602 467236 325608 467248
rect 325660 467236 325666 467288
rect 262766 467168 262772 467220
rect 262824 467208 262830 467220
rect 527174 467208 527180 467220
rect 262824 467180 527180 467208
rect 262824 467168 262830 467180
rect 527174 467168 527180 467180
rect 527232 467168 527238 467220
rect 4798 467100 4804 467152
rect 4856 467140 4862 467152
rect 281718 467140 281724 467152
rect 4856 467112 281724 467140
rect 4856 467100 4862 467112
rect 281718 467100 281724 467112
rect 281776 467100 281782 467152
rect 306282 467100 306288 467152
rect 306340 467140 306346 467152
rect 348510 467140 348516 467152
rect 306340 467112 348516 467140
rect 306340 467100 306346 467112
rect 348510 467100 348516 467112
rect 348568 467100 348574 467152
rect 268930 465944 268936 465996
rect 268988 465984 268994 465996
rect 291838 465984 291844 465996
rect 268988 465956 291844 465984
rect 268988 465944 268994 465956
rect 291838 465944 291844 465956
rect 291896 465944 291902 465996
rect 277210 465876 277216 465928
rect 277268 465916 277274 465928
rect 355686 465916 355692 465928
rect 277268 465888 355692 465916
rect 277268 465876 277274 465888
rect 355686 465876 355692 465888
rect 355744 465876 355750 465928
rect 218882 465808 218888 465860
rect 218940 465848 218946 465860
rect 307294 465848 307300 465860
rect 218940 465820 307300 465848
rect 218940 465808 218946 465820
rect 307294 465808 307300 465820
rect 307352 465808 307358 465860
rect 258810 465740 258816 465792
rect 258868 465780 258874 465792
rect 373258 465780 373264 465792
rect 258868 465752 373264 465780
rect 258868 465740 258874 465752
rect 373258 465740 373264 465752
rect 373316 465740 373322 465792
rect 21358 465672 21364 465724
rect 21416 465712 21422 465724
rect 279786 465712 279792 465724
rect 21416 465684 279792 465712
rect 21416 465672 21422 465684
rect 279786 465672 279792 465684
rect 279844 465672 279850 465724
rect 299382 465672 299388 465724
rect 299440 465712 299446 465724
rect 344554 465712 344560 465724
rect 299440 465684 344560 465712
rect 299440 465672 299446 465684
rect 344554 465672 344560 465684
rect 344612 465672 344618 465724
rect 246942 464448 246948 464500
rect 247000 464488 247006 464500
rect 317782 464488 317788 464500
rect 247000 464460 317788 464488
rect 247000 464448 247006 464460
rect 317782 464448 317788 464460
rect 317840 464448 317846 464500
rect 218054 464380 218060 464432
rect 218112 464420 218118 464432
rect 273254 464420 273260 464432
rect 218112 464392 273260 464420
rect 218112 464380 218118 464392
rect 273254 464380 273260 464392
rect 273312 464380 273318 464432
rect 274450 464380 274456 464432
rect 274508 464420 274514 464432
rect 351822 464420 351828 464432
rect 274508 464392 351828 464420
rect 274508 464380 274514 464392
rect 351822 464380 351828 464392
rect 351880 464380 351886 464432
rect 266722 464312 266728 464364
rect 266780 464352 266786 464364
rect 396718 464352 396724 464364
rect 266780 464324 396724 464352
rect 266780 464312 266786 464324
rect 396718 464312 396724 464324
rect 396776 464312 396782 464364
rect 293862 463156 293868 463208
rect 293920 463196 293926 463208
rect 341978 463196 341984 463208
rect 293920 463168 341984 463196
rect 293920 463156 293926 463168
rect 341978 463156 341984 463168
rect 342036 463156 342042 463208
rect 244182 463088 244188 463140
rect 244240 463128 244246 463140
rect 309870 463128 309876 463140
rect 244240 463100 309876 463128
rect 244240 463088 244246 463100
rect 309870 463088 309876 463100
rect 309928 463088 309934 463140
rect 249702 463020 249708 463072
rect 249760 463060 249766 463072
rect 322290 463060 322296 463072
rect 249760 463032 322296 463060
rect 249760 463020 249766 463032
rect 322290 463020 322296 463032
rect 322348 463020 322354 463072
rect 260834 462952 260840 463004
rect 260892 462992 260898 463004
rect 391198 462992 391204 463004
rect 260892 462964 391204 462992
rect 260892 462952 260898 462964
rect 391198 462952 391204 462964
rect 391256 462952 391262 463004
rect 3234 462340 3240 462392
rect 3292 462380 3298 462392
rect 288986 462380 288992 462392
rect 3292 462352 288992 462380
rect 3292 462340 3298 462352
rect 288986 462340 288992 462352
rect 289044 462340 289050 462392
rect 210418 461796 210424 461848
rect 210476 461836 210482 461848
rect 285030 461836 285036 461848
rect 210476 461808 285036 461836
rect 210476 461796 210482 461808
rect 285030 461796 285036 461808
rect 285088 461796 285094 461848
rect 262030 461728 262036 461780
rect 262088 461768 262094 461780
rect 338666 461768 338672 461780
rect 262088 461740 338672 461768
rect 262088 461728 262094 461740
rect 338666 461728 338672 461740
rect 338724 461728 338730 461780
rect 268010 461660 268016 461712
rect 268068 461700 268074 461712
rect 364334 461700 364340 461712
rect 268068 461672 364340 461700
rect 268068 461660 268074 461672
rect 364334 461660 364340 461672
rect 364392 461660 364398 461712
rect 71774 461592 71780 461644
rect 71832 461632 71838 461644
rect 276474 461632 276480 461644
rect 71832 461604 276480 461632
rect 71832 461592 71838 461604
rect 276474 461592 276480 461604
rect 276532 461592 276538 461644
rect 291102 461592 291108 461644
rect 291160 461632 291166 461644
rect 340690 461632 340696 461644
rect 291160 461604 340696 461632
rect 291160 461592 291166 461604
rect 340690 461592 340696 461604
rect 340748 461592 340754 461644
rect 250990 460368 250996 460420
rect 251048 460408 251054 460420
rect 313182 460408 313188 460420
rect 251048 460380 313188 460408
rect 251048 460368 251054 460380
rect 313182 460368 313188 460380
rect 313240 460368 313246 460420
rect 239398 460300 239404 460352
rect 239456 460340 239462 460352
rect 309226 460340 309232 460352
rect 239456 460312 309232 460340
rect 239456 460300 239462 460312
rect 309226 460300 309232 460312
rect 309284 460300 309290 460352
rect 265986 460232 265992 460284
rect 266044 460272 266050 460284
rect 359458 460272 359464 460284
rect 266044 460244 359464 460272
rect 266044 460232 266050 460244
rect 359458 460232 359464 460244
rect 359516 460232 359522 460284
rect 10318 460164 10324 460216
rect 10376 460204 10382 460216
rect 278498 460204 278504 460216
rect 10376 460176 278504 460204
rect 10376 460164 10382 460176
rect 278498 460164 278504 460176
rect 278556 460164 278562 460216
rect 278590 460164 278596 460216
rect 278648 460204 278654 460216
rect 357066 460204 357072 460216
rect 278648 460176 357072 460204
rect 278648 460164 278654 460176
rect 357066 460164 357072 460176
rect 357124 460164 357130 460216
rect 214558 459008 214564 459060
rect 214616 459048 214622 459060
rect 281074 459048 281080 459060
rect 214616 459020 281080 459048
rect 214616 459008 214622 459020
rect 281074 459008 281080 459020
rect 281132 459008 281138 459060
rect 259362 458940 259368 458992
rect 259420 458980 259426 458992
rect 334802 458980 334808 458992
rect 259420 458952 334808 458980
rect 259420 458940 259426 458952
rect 334802 458940 334808 458952
rect 334860 458940 334866 458992
rect 138658 458872 138664 458924
rect 138716 458912 138722 458924
rect 274542 458912 274548 458924
rect 138716 458884 274548 458912
rect 138716 458872 138722 458884
rect 274542 458872 274548 458884
rect 274600 458872 274606 458924
rect 281442 458872 281448 458924
rect 281500 458912 281506 458924
rect 335446 458912 335452 458924
rect 281500 458884 335452 458912
rect 281500 458872 281506 458884
rect 335446 458872 335452 458884
rect 335504 458872 335510 458924
rect 264054 458804 264060 458856
rect 264112 458844 264118 458856
rect 494054 458844 494060 458856
rect 264112 458816 494060 458844
rect 264112 458804 264118 458816
rect 494054 458804 494060 458816
rect 494112 458804 494118 458856
rect 251082 457580 251088 457632
rect 251140 457620 251146 457632
rect 324314 457620 324320 457632
rect 251140 457592 324320 457620
rect 251140 457580 251146 457592
rect 324314 457580 324320 457592
rect 324372 457580 324378 457632
rect 256510 457512 256516 457564
rect 256568 457552 256574 457564
rect 332134 457552 332140 457564
rect 256568 457524 332140 457552
rect 256568 457512 256574 457524
rect 332134 457512 332140 457524
rect 332192 457512 332198 457564
rect 28258 457444 28264 457496
rect 28316 457484 28322 457496
rect 280430 457484 280436 457496
rect 28316 457456 280436 457484
rect 28316 457444 28322 457456
rect 280430 457444 280436 457456
rect 280488 457444 280494 457496
rect 252278 456764 252284 456816
rect 252336 456804 252342 456816
rect 580166 456804 580172 456816
rect 252336 456776 580172 456804
rect 252336 456764 252342 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 215938 456220 215944 456272
rect 215996 456260 216002 456272
rect 279142 456260 279148 456272
rect 215996 456232 279148 456260
rect 215996 456220 216002 456232
rect 279142 456220 279148 456232
rect 279200 456220 279206 456272
rect 201494 456152 201500 456204
rect 201552 456192 201558 456204
rect 272610 456192 272616 456204
rect 201552 456164 272616 456192
rect 201552 456152 201558 456164
rect 272610 456152 272616 456164
rect 272668 456152 272674 456204
rect 278682 456152 278688 456204
rect 278740 456192 278746 456204
rect 334158 456192 334164 456204
rect 278740 456164 334164 456192
rect 278740 456152 278746 456164
rect 334158 456152 334164 456164
rect 334216 456152 334222 456204
rect 260650 456084 260656 456136
rect 260708 456124 260714 456136
rect 336090 456124 336096 456136
rect 260708 456096 336096 456124
rect 260708 456084 260714 456096
rect 336090 456084 336096 456096
rect 336148 456084 336154 456136
rect 262122 456016 262128 456068
rect 262180 456056 262186 456068
rect 442258 456056 442264 456068
rect 262180 456028 442264 456056
rect 262180 456016 262186 456028
rect 442258 456016 442264 456028
rect 442316 456016 442322 456068
rect 237190 454792 237196 454844
rect 237248 454832 237254 454844
rect 311894 454832 311900 454844
rect 237248 454804 311900 454832
rect 237248 454792 237254 454804
rect 311894 454792 311900 454804
rect 311952 454792 311958 454844
rect 260098 454724 260104 454776
rect 260156 454764 260162 454776
rect 377398 454764 377404 454776
rect 260156 454736 377404 454764
rect 260156 454724 260162 454736
rect 377398 454724 377404 454736
rect 377456 454724 377462 454776
rect 40034 454656 40040 454708
rect 40092 454696 40098 454708
rect 277854 454696 277860 454708
rect 40092 454668 277860 454696
rect 40092 454656 40098 454668
rect 277854 454656 277860 454668
rect 277912 454656 277918 454708
rect 280062 454656 280068 454708
rect 280120 454696 280126 454708
rect 358354 454696 358360 454708
rect 280120 454668 358360 454696
rect 280120 454656 280126 454668
rect 358354 454656 358360 454668
rect 358412 454656 358418 454708
rect 248322 453568 248328 453620
rect 248380 453608 248386 453620
rect 310514 453608 310520 453620
rect 248380 453580 310520 453608
rect 248380 453568 248386 453580
rect 310514 453568 310520 453580
rect 310572 453568 310578 453620
rect 211798 453500 211804 453552
rect 211856 453540 211862 453552
rect 283006 453540 283012 453552
rect 211856 453512 283012 453540
rect 211856 453500 211862 453512
rect 283006 453500 283012 453512
rect 283064 453500 283070 453552
rect 271690 453432 271696 453484
rect 271748 453472 271754 453484
rect 349154 453472 349160 453484
rect 271748 453444 349160 453472
rect 271748 453432 271754 453444
rect 349154 453432 349160 453444
rect 349212 453432 349218 453484
rect 169754 453364 169760 453416
rect 169812 453404 169818 453416
rect 273898 453404 273904 453416
rect 169812 453376 273904 453404
rect 169812 453364 169818 453376
rect 273898 453364 273904 453376
rect 273956 453364 273962 453416
rect 302142 453364 302148 453416
rect 302200 453404 302206 453416
rect 345934 453404 345940 453416
rect 302200 453376 345940 453404
rect 302200 453364 302206 453376
rect 345934 453364 345940 453376
rect 345992 453364 345998 453416
rect 258166 453296 258172 453348
rect 258224 453336 258230 453348
rect 363598 453336 363604 453348
rect 258224 453308 363604 453336
rect 258224 453296 258230 453308
rect 363598 453296 363604 453308
rect 363656 453296 363662 453348
rect 273162 452072 273168 452124
rect 273220 452112 273226 452124
rect 350534 452112 350540 452124
rect 273220 452084 350540 452112
rect 273220 452072 273226 452084
rect 350534 452072 350540 452084
rect 350592 452072 350598 452124
rect 207658 452004 207664 452056
rect 207716 452044 207722 452056
rect 286962 452044 286968 452056
rect 207716 452016 286968 452044
rect 207716 452004 207722 452016
rect 286962 452004 286968 452016
rect 287020 452004 287026 452056
rect 256234 451936 256240 451988
rect 256292 451976 256298 451988
rect 360838 451976 360844 451988
rect 256292 451948 360844 451976
rect 256292 451936 256298 451948
rect 360838 451936 360844 451948
rect 360896 451936 360902 451988
rect 108298 451868 108304 451920
rect 108356 451908 108362 451920
rect 275830 451908 275836 451920
rect 108356 451880 275836 451908
rect 108356 451868 108362 451880
rect 275830 451868 275836 451880
rect 275888 451868 275894 451920
rect 284202 451868 284208 451920
rect 284260 451908 284266 451920
rect 336734 451908 336740 451920
rect 284260 451880 336740 451908
rect 284260 451868 284266 451880
rect 336734 451868 336740 451880
rect 336792 451868 336798 451920
rect 260742 450644 260748 450696
rect 260800 450684 260806 450696
rect 337378 450684 337384 450696
rect 260800 450656 337384 450684
rect 260800 450644 260806 450656
rect 337378 450644 337384 450656
rect 337436 450644 337442 450696
rect 254210 450576 254216 450628
rect 254268 450616 254274 450628
rect 358078 450616 358084 450628
rect 254268 450588 358084 450616
rect 254268 450576 254274 450588
rect 358078 450576 358084 450588
rect 358136 450576 358142 450628
rect 88334 450508 88340 450560
rect 88392 450548 88398 450560
rect 277118 450548 277124 450560
rect 88392 450520 277124 450548
rect 88392 450508 88398 450520
rect 277118 450508 277124 450520
rect 277176 450508 277182 450560
rect 277302 450508 277308 450560
rect 277360 450548 277366 450560
rect 332778 450548 332784 450560
rect 277360 450520 332784 450548
rect 277360 450508 277366 450520
rect 332778 450508 332784 450520
rect 332836 450508 332842 450560
rect 245562 449692 245568 449744
rect 245620 449732 245626 449744
rect 312538 449732 312544 449744
rect 245620 449704 312544 449732
rect 245620 449692 245626 449704
rect 312538 449692 312544 449704
rect 312596 449692 312602 449744
rect 245470 449624 245476 449676
rect 245528 449664 245534 449676
rect 315114 449664 315120 449676
rect 245528 449636 315120 449664
rect 245528 449624 245534 449636
rect 315114 449624 315120 449636
rect 315172 449624 315178 449676
rect 266170 449556 266176 449608
rect 266228 449596 266234 449608
rect 342622 449596 342628 449608
rect 266228 449568 342628 449596
rect 266228 449556 266234 449568
rect 342622 449556 342628 449568
rect 342680 449556 342686 449608
rect 264882 449488 264888 449540
rect 264940 449528 264946 449540
rect 341334 449528 341340 449540
rect 264940 449500 341340 449528
rect 264940 449488 264946 449500
rect 341334 449488 341340 449500
rect 341392 449488 341398 449540
rect 267642 449420 267648 449472
rect 267700 449460 267706 449472
rect 343910 449460 343916 449472
rect 267700 449432 343916 449460
rect 267700 449420 267706 449432
rect 343910 449420 343916 449432
rect 343968 449420 343974 449472
rect 263502 449352 263508 449404
rect 263560 449392 263566 449404
rect 340046 449392 340052 449404
rect 263560 449364 340052 449392
rect 263560 449352 263566 449364
rect 340046 449352 340052 449364
rect 340104 449352 340110 449404
rect 269022 449284 269028 449336
rect 269080 449324 269086 449336
rect 346578 449324 346584 449336
rect 269080 449296 346584 449324
rect 269080 449284 269086 449296
rect 346578 449284 346584 449296
rect 346636 449284 346642 449336
rect 270402 449216 270408 449268
rect 270460 449256 270466 449268
rect 347866 449256 347872 449268
rect 270460 449228 347872 449256
rect 270460 449216 270466 449228
rect 347866 449216 347872 449228
rect 347924 449216 347930 449268
rect 267550 449148 267556 449200
rect 267608 449188 267614 449200
rect 345290 449188 345296 449200
rect 267608 449160 345296 449188
rect 267608 449148 267614 449160
rect 345290 449148 345296 449160
rect 345348 449148 345354 449200
rect 257982 447992 257988 448044
rect 258040 448032 258046 448044
rect 333422 448032 333428 448044
rect 258040 448004 333428 448032
rect 258040 447992 258046 448004
rect 333422 447992 333428 448004
rect 333480 447992 333486 448044
rect 252462 447924 252468 447976
rect 252520 447964 252526 447976
rect 328270 447964 328276 447976
rect 252520 447936 328276 447964
rect 252520 447924 252526 447936
rect 328270 447924 328276 447936
rect 328328 447924 328334 447976
rect 274358 447856 274364 447908
rect 274416 447896 274422 447908
rect 353110 447896 353116 447908
rect 274416 447868 353116 447896
rect 274416 447856 274422 447868
rect 353110 447856 353116 447868
rect 353168 447856 353174 447908
rect 217318 447788 217324 447840
rect 217376 447828 217382 447840
rect 307938 447828 307944 447840
rect 217376 447800 307944 447828
rect 217376 447788 217382 447800
rect 307938 447788 307944 447800
rect 307996 447788 308002 447840
rect 267366 446700 267372 446752
rect 267424 446740 267430 446752
rect 412634 446740 412640 446752
rect 267424 446712 412640 446740
rect 267424 446700 267430 446712
rect 412634 446700 412640 446712
rect 412692 446700 412698 446752
rect 265342 446632 265348 446684
rect 265400 446672 265406 446684
rect 477494 446672 477500 446684
rect 265400 446644 477500 446672
rect 265400 446632 265406 446644
rect 477494 446632 477500 446644
rect 477552 446632 477558 446684
rect 263410 446564 263416 446616
rect 263468 446604 263474 446616
rect 542354 446604 542360 446616
rect 263468 446576 542360 446604
rect 263468 446564 263474 446576
rect 542354 446564 542360 446576
rect 542412 446564 542418 446616
rect 4154 446496 4160 446548
rect 4212 446536 4218 446548
rect 288250 446536 288256 446548
rect 4212 446508 288256 446536
rect 4212 446496 4218 446508
rect 288250 446496 288256 446508
rect 288308 446496 288314 446548
rect 259454 446428 259460 446480
rect 259512 446468 259518 446480
rect 580258 446468 580264 446480
rect 259512 446440 580264 446468
rect 259512 446428 259518 446440
rect 580258 446428 580264 446440
rect 580316 446428 580322 446480
rect 257522 446360 257528 446412
rect 257580 446400 257586 446412
rect 580350 446400 580356 446412
rect 257580 446372 580356 446400
rect 257580 446360 257586 446372
rect 580350 446360 580356 446372
rect 580408 446360 580414 446412
rect 206278 446020 206284 446072
rect 206336 446060 206342 446072
rect 300118 446060 300124 446072
rect 206336 446032 300124 446060
rect 206336 446020 206342 446032
rect 300118 446020 300124 446032
rect 300176 446020 300182 446072
rect 203610 445952 203616 446004
rect 203668 445992 203674 446004
rect 298094 445992 298100 446004
rect 203668 445964 298100 445992
rect 203668 445952 203674 445964
rect 298094 445952 298100 445964
rect 298152 445952 298158 446004
rect 192478 445884 192484 445936
rect 192536 445924 192542 445936
rect 302694 445924 302700 445936
rect 192536 445896 302700 445924
rect 192536 445884 192542 445896
rect 302694 445884 302700 445896
rect 302752 445884 302758 445936
rect 235902 445816 235908 445868
rect 235960 445856 235966 445868
rect 373258 445856 373264 445868
rect 235960 445828 373264 445856
rect 235960 445816 235966 445828
rect 373258 445816 373264 445828
rect 373316 445816 373322 445868
rect 8938 445748 8944 445800
rect 8996 445788 9002 445800
rect 296806 445788 296812 445800
rect 8996 445760 296812 445788
rect 8996 445748 9002 445760
rect 296806 445748 296812 445760
rect 296864 445748 296870 445800
rect 231118 444864 231124 444916
rect 231176 444904 231182 444916
rect 290274 444904 290280 444916
rect 231176 444876 290280 444904
rect 231176 444864 231182 444876
rect 290274 444864 290280 444876
rect 290332 444864 290338 444916
rect 225598 444796 225604 444848
rect 225656 444836 225662 444848
rect 295518 444836 295524 444848
rect 225656 444808 295524 444836
rect 225656 444796 225662 444808
rect 295518 444796 295524 444808
rect 295576 444796 295582 444848
rect 199378 444728 199384 444780
rect 199436 444768 199442 444780
rect 303982 444768 303988 444780
rect 199436 444740 303988 444768
rect 199436 444728 199442 444740
rect 303982 444728 303988 444740
rect 304040 444728 304046 444780
rect 249702 444660 249708 444712
rect 249760 444700 249766 444712
rect 378778 444700 378784 444712
rect 249760 444672 378784 444700
rect 249760 444660 249766 444672
rect 378778 444660 378784 444672
rect 378836 444660 378842 444712
rect 100018 444592 100024 444644
rect 100076 444632 100082 444644
rect 291562 444632 291568 444644
rect 100076 444604 291568 444632
rect 100076 444592 100082 444604
rect 291562 444592 291568 444604
rect 291620 444592 291626 444644
rect 98638 444524 98644 444576
rect 98696 444564 98702 444576
rect 293494 444564 293500 444576
rect 98696 444536 293500 444564
rect 98696 444524 98702 444536
rect 293494 444524 293500 444536
rect 293552 444524 293558 444576
rect 7558 444456 7564 444508
rect 7616 444496 7622 444508
rect 289630 444496 289636 444508
rect 7616 444468 289636 444496
rect 7616 444456 7622 444468
rect 289630 444456 289636 444468
rect 289688 444456 289694 444508
rect 244458 444388 244464 444440
rect 244516 444428 244522 444440
rect 578878 444428 578884 444440
rect 244516 444400 578884 444428
rect 244516 444388 244522 444400
rect 578878 444388 578884 444400
rect 578936 444388 578942 444440
rect 245746 444116 245752 444168
rect 245804 444156 245810 444168
rect 362218 444156 362224 444168
rect 245804 444128 362224 444156
rect 245804 444116 245810 444128
rect 362218 444116 362224 444128
rect 362276 444116 362282 444168
rect 335998 444048 336004 444100
rect 336056 444088 336062 444100
rect 355042 444088 355048 444100
rect 336056 444060 355048 444088
rect 336056 444048 336062 444060
rect 355042 444048 355048 444060
rect 355100 444048 355106 444100
rect 334618 443980 334624 444032
rect 334676 444020 334682 444032
rect 353754 444020 353760 444032
rect 334676 443992 353760 444020
rect 334676 443980 334682 443992
rect 353754 443980 353760 443992
rect 353812 443980 353818 444032
rect 252554 443912 252560 443964
rect 252612 443952 252618 443964
rect 301406 443952 301412 443964
rect 252612 443924 301412 443952
rect 252612 443912 252618 443924
rect 301406 443912 301412 443924
rect 301464 443912 301470 443964
rect 331858 443912 331864 443964
rect 331916 443952 331922 443964
rect 351178 443952 351184 443964
rect 331916 443924 351184 443952
rect 331916 443912 331922 443924
rect 351178 443912 351184 443924
rect 351236 443912 351242 443964
rect 239214 443844 239220 443896
rect 239272 443884 239278 443896
rect 282914 443884 282920 443896
rect 239272 443856 282920 443884
rect 239272 443844 239278 443856
rect 282914 443844 282920 443856
rect 282972 443844 282978 443896
rect 294598 443844 294604 443896
rect 294656 443884 294662 443896
rect 321002 443884 321008 443896
rect 294656 443856 321008 443884
rect 294656 443844 294662 443856
rect 321002 443844 321008 443856
rect 321060 443844 321066 443896
rect 333238 443844 333244 443896
rect 333296 443884 333302 443896
rect 352466 443884 352472 443896
rect 333296 443856 352472 443884
rect 333296 443844 333302 443856
rect 352466 443844 352472 443856
rect 352524 443844 352530 443896
rect 94498 443776 94504 443828
rect 94556 443816 94562 443828
rect 294874 443816 294880 443828
rect 94556 443788 294880 443816
rect 94556 443776 94562 443788
rect 294874 443776 294880 443788
rect 294932 443776 294938 443828
rect 295978 443776 295984 443828
rect 296036 443816 296042 443828
rect 324958 443816 324964 443828
rect 296036 443788 324964 443816
rect 296036 443776 296042 443788
rect 324958 443776 324964 443788
rect 325016 443776 325022 443828
rect 338758 443776 338764 443828
rect 338816 443816 338822 443828
rect 358998 443816 359004 443828
rect 338816 443788 359004 443816
rect 338816 443776 338822 443788
rect 358998 443776 359004 443788
rect 359056 443776 359062 443828
rect 219342 443708 219348 443760
rect 219400 443748 219406 443760
rect 270586 443748 270592 443760
rect 219400 443720 270592 443748
rect 219400 443708 219406 443720
rect 270586 443708 270592 443720
rect 270644 443708 270650 443760
rect 291838 443708 291844 443760
rect 291896 443748 291902 443760
rect 328914 443748 328920 443760
rect 291896 443720 328920 443748
rect 291896 443708 291902 443720
rect 328914 443708 328920 443720
rect 328972 443708 328978 443760
rect 329098 443708 329104 443760
rect 329156 443748 329162 443760
rect 349798 443748 349804 443760
rect 329156 443720 349804 443748
rect 329156 443708 329162 443720
rect 349798 443708 349804 443720
rect 349856 443708 349862 443760
rect 217778 443640 217784 443692
rect 217836 443680 217842 443692
rect 271966 443680 271972 443692
rect 217836 443652 271972 443680
rect 217836 443640 217842 443652
rect 271966 443640 271972 443652
rect 272024 443640 272030 443692
rect 303522 443640 303528 443692
rect 303580 443680 303586 443692
rect 347222 443680 347228 443692
rect 303580 443652 347228 443680
rect 303580 443640 303586 443652
rect 347222 443640 347228 443652
rect 347280 443640 347286 443692
rect 352558 443640 352564 443692
rect 352616 443680 352622 443692
rect 357710 443680 357716 443692
rect 352616 443652 357716 443680
rect 352616 443640 352622 443652
rect 357710 443640 357716 443652
rect 357768 443640 357774 443692
rect 246390 443572 246396 443624
rect 246448 443612 246454 443624
rect 277394 443612 277400 443624
rect 246448 443584 277400 443612
rect 246448 443572 246454 443584
rect 277394 443572 277400 443584
rect 277452 443572 277458 443624
rect 241146 443504 241152 443556
rect 241204 443544 241210 443556
rect 274726 443544 274732 443556
rect 241204 443516 274732 443544
rect 241204 443504 241210 443516
rect 274726 443504 274732 443516
rect 274784 443504 274790 443556
rect 245102 443436 245108 443488
rect 245160 443476 245166 443488
rect 288342 443476 288348 443488
rect 245160 443448 288348 443476
rect 245160 443436 245166 443448
rect 288342 443436 288348 443448
rect 288400 443436 288406 443488
rect 248322 443368 248328 443420
rect 248380 443408 248386 443420
rect 276106 443408 276112 443420
rect 248380 443380 276112 443408
rect 248380 443368 248386 443380
rect 276106 443368 276112 443380
rect 276164 443368 276170 443420
rect 279510 443368 279516 443420
rect 279568 443408 279574 443420
rect 296162 443408 296168 443420
rect 279568 443380 296168 443408
rect 279568 443368 279574 443380
rect 296162 443368 296168 443380
rect 296220 443368 296226 443420
rect 229738 443300 229744 443352
rect 229796 443340 229802 443352
rect 253198 443340 253204 443352
rect 229796 443312 253204 443340
rect 229796 443300 229802 443312
rect 253198 443300 253204 443312
rect 253256 443340 253262 443352
rect 253566 443340 253572 443352
rect 253256 443312 253572 443340
rect 253256 443300 253262 443312
rect 253566 443300 253572 443312
rect 253624 443300 253630 443352
rect 224218 443232 224224 443284
rect 224276 443272 224282 443284
rect 292850 443272 292856 443284
rect 224276 443244 292856 443272
rect 224276 443232 224282 443244
rect 292850 443232 292856 443244
rect 292908 443232 292914 443284
rect 196710 443164 196716 443216
rect 196768 443204 196774 443216
rect 298738 443204 298744 443216
rect 196768 443176 298744 443204
rect 196768 443164 196774 443176
rect 298738 443164 298744 443176
rect 298796 443164 298802 443216
rect 359642 443164 359648 443216
rect 359700 443204 359706 443216
rect 388438 443204 388444 443216
rect 359700 443176 388444 443204
rect 359700 443164 359706 443176
rect 388438 443164 388444 443176
rect 388496 443164 388502 443216
rect 140774 443096 140780 443148
rect 140832 443136 140838 443148
rect 250346 443136 250352 443148
rect 140832 443108 250352 443136
rect 140832 443096 140838 443108
rect 250346 443096 250352 443108
rect 250404 443136 250410 443148
rect 362494 443136 362500 443148
rect 250404 443108 362500 443136
rect 250404 443096 250410 443108
rect 362494 443096 362500 443108
rect 362552 443096 362558 443148
rect 233970 443028 233976 443080
rect 234028 443068 234034 443080
rect 246942 443068 246948 443080
rect 234028 443040 246948 443068
rect 234028 443028 234034 443040
rect 246942 443028 246948 443040
rect 247000 443028 247006 443080
rect 269022 443028 269028 443080
rect 269080 443068 269086 443080
rect 292206 443068 292212 443080
rect 269080 443040 292212 443068
rect 269080 443028 269086 443040
rect 292206 443028 292212 443040
rect 292264 443028 292270 443080
rect 360286 443028 360292 443080
rect 360344 443068 360350 443080
rect 581086 443068 581092 443080
rect 360344 443040 581092 443068
rect 360344 443028 360350 443040
rect 581086 443028 581092 443040
rect 581144 443028 581150 443080
rect 250990 442960 250996 443012
rect 251048 443000 251054 443012
rect 268562 443000 268568 443012
rect 251048 442972 268568 443000
rect 251048 442960 251054 442972
rect 268562 442960 268568 442972
rect 268620 442960 268626 443012
rect 274634 442960 274640 443012
rect 274692 443000 274698 443012
rect 294138 443000 294144 443012
rect 274692 442972 294144 443000
rect 274692 442960 274698 442972
rect 294138 442960 294144 442972
rect 294196 442960 294202 443012
rect 360930 442960 360936 443012
rect 360988 443000 360994 443012
rect 582374 443000 582380 443012
rect 360988 442972 582380 443000
rect 360988 442960 360994 442972
rect 582374 442960 582380 442972
rect 582432 442960 582438 443012
rect 231210 442484 231216 442536
rect 231268 442524 231274 442536
rect 290918 442524 290924 442536
rect 231268 442496 290924 442524
rect 231268 442484 231274 442496
rect 290918 442484 290924 442496
rect 290976 442484 290982 442536
rect 3602 442416 3608 442468
rect 3660 442456 3666 442468
rect 274634 442456 274640 442468
rect 3660 442428 274640 442456
rect 3660 442416 3666 442428
rect 274634 442416 274640 442428
rect 274692 442416 274698 442468
rect 288342 442416 288348 442468
rect 288400 442456 288406 442468
rect 580810 442456 580816 442468
rect 288400 442428 580816 442456
rect 288400 442416 288406 442428
rect 580810 442416 580816 442428
rect 580868 442416 580874 442468
rect 3510 442348 3516 442400
rect 3568 442388 3574 442400
rect 279510 442388 279516 442400
rect 3568 442360 279516 442388
rect 3568 442348 3574 442360
rect 279510 442348 279516 442360
rect 279568 442348 279574 442400
rect 282914 442348 282920 442400
rect 282972 442388 282978 442400
rect 580626 442388 580632 442400
rect 282972 442360 580632 442388
rect 282972 442348 282978 442360
rect 580626 442348 580632 442360
rect 580684 442348 580690 442400
rect 269022 442320 269028 442332
rect 253906 442292 269028 442320
rect 3694 442212 3700 442264
rect 3752 442252 3758 442264
rect 253906 442252 253934 442292
rect 269022 442280 269028 442292
rect 269080 442280 269086 442332
rect 274726 442280 274732 442332
rect 274784 442320 274790 442332
rect 580718 442320 580724 442332
rect 274784 442292 580724 442320
rect 274784 442280 274790 442292
rect 580718 442280 580724 442292
rect 580776 442280 580782 442332
rect 3752 442224 253934 442252
rect 3752 442212 3758 442224
rect 268562 442212 268568 442264
rect 268620 442252 268626 442264
rect 580074 442252 580080 442264
rect 268620 442224 580080 442252
rect 268620 442212 268626 442224
rect 580074 442212 580080 442224
rect 580132 442212 580138 442264
rect 200758 442144 200764 442196
rect 200816 442184 200822 442196
rect 302050 442184 302056 442196
rect 200816 442156 302056 442184
rect 200816 442144 200822 442156
rect 302050 442144 302056 442156
rect 302108 442144 302114 442196
rect 197998 442076 198004 442128
rect 198056 442116 198062 442128
rect 300762 442116 300768 442128
rect 198056 442088 300768 442116
rect 198056 442076 198062 442088
rect 300762 442076 300768 442088
rect 300820 442076 300826 442128
rect 248966 442008 248972 442060
rect 249024 442048 249030 442060
rect 362402 442048 362408 442060
rect 249024 442020 362408 442048
rect 249024 442008 249030 442020
rect 362402 442008 362408 442020
rect 362460 442008 362466 442060
rect 247034 441940 247040 441992
rect 247092 441980 247098 441992
rect 362310 441980 362316 441992
rect 247092 441952 362316 441980
rect 247092 441940 247098 441952
rect 362310 441940 362316 441952
rect 362368 441940 362374 441992
rect 241790 441872 241796 441924
rect 241848 441912 241854 441924
rect 374730 441912 374736 441924
rect 241848 441884 374736 441912
rect 241848 441872 241854 441884
rect 374730 441872 374736 441884
rect 374788 441872 374794 441924
rect 64138 441804 64144 441856
rect 64196 441844 64202 441856
rect 306650 441844 306656 441856
rect 64196 441816 306656 441844
rect 64196 441804 64202 441816
rect 306650 441804 306656 441816
rect 306708 441804 306714 441856
rect 242434 441736 242440 441788
rect 242492 441776 242498 441788
rect 577590 441776 577596 441788
rect 242492 441748 577596 441776
rect 242492 441736 242498 441748
rect 577590 441736 577596 441748
rect 577648 441736 577654 441788
rect 237190 441668 237196 441720
rect 237248 441708 237254 441720
rect 580442 441708 580448 441720
rect 237248 441680 580448 441708
rect 237248 441668 237254 441680
rect 580442 441668 580448 441680
rect 580500 441668 580506 441720
rect 233326 441600 233332 441652
rect 233384 441640 233390 441652
rect 577498 441640 577504 441652
rect 233384 441612 577504 441640
rect 233384 441600 233390 441612
rect 577498 441600 577504 441612
rect 577556 441600 577562 441652
rect 289998 441396 290004 441448
rect 290056 441436 290062 441448
rect 294598 441436 294604 441448
rect 290056 441408 294604 441436
rect 290056 441396 290062 441408
rect 294598 441396 294604 441408
rect 294656 441396 294662 441448
rect 289786 441340 302234 441368
rect 252554 441164 252560 441176
rect 234586 441136 252560 441164
rect 3418 440852 3424 440904
rect 3476 440892 3482 440904
rect 234586 440892 234614 441136
rect 252554 441124 252560 441136
rect 252612 441124 252618 441176
rect 289786 441096 289814 441340
rect 293586 441300 293592 441312
rect 290936 441272 293592 441300
rect 290734 441124 290740 441176
rect 290792 441124 290798 441176
rect 3476 440864 234614 440892
rect 240106 441068 256694 441096
rect 3476 440852 3482 440864
rect 207658 440580 207664 440632
rect 207716 440620 207722 440632
rect 240106 440620 240134 441068
rect 240778 440988 240784 441040
rect 240836 440988 240842 441040
rect 247954 440988 247960 441040
rect 248012 440988 248018 441040
rect 252002 440988 252008 441040
rect 252060 440988 252066 441040
rect 207716 440592 240134 440620
rect 207716 440580 207722 440592
rect 240796 440416 240824 440988
rect 247972 440484 248000 440988
rect 252020 440552 252048 440988
rect 256666 440824 256694 441068
rect 287026 441068 289814 441096
rect 276106 440988 276112 441040
rect 276164 440988 276170 441040
rect 277394 440988 277400 441040
rect 277452 440988 277458 441040
rect 276124 440892 276152 440988
rect 277412 440960 277440 440988
rect 287026 440960 287054 441068
rect 289814 441028 289820 441040
rect 277412 440932 287054 440960
rect 289786 440988 289820 441028
rect 289872 440988 289878 441040
rect 289998 440988 290004 441040
rect 290056 440988 290062 441040
rect 289786 440892 289814 440988
rect 259426 440864 260834 440892
rect 276124 440864 289814 440892
rect 259426 440824 259454 440864
rect 256666 440796 259454 440824
rect 260806 440688 260834 440864
rect 290016 440688 290044 440988
rect 260806 440660 263594 440688
rect 263566 440620 263594 440660
rect 289786 440660 290044 440688
rect 289786 440620 289814 440660
rect 263566 440592 289814 440620
rect 290752 440552 290780 441124
rect 252020 440524 290780 440552
rect 290936 440484 290964 441272
rect 293586 441260 293592 441272
rect 293644 441260 293650 441312
rect 293402 441232 293408 441244
rect 291304 441204 293408 441232
rect 291304 440960 291332 441204
rect 293402 441192 293408 441204
rect 293460 441192 293466 441244
rect 294598 441192 294604 441244
rect 294656 441232 294662 441244
rect 294656 441204 300854 441232
rect 294656 441192 294662 441204
rect 292224 441068 299474 441096
rect 291304 440932 291424 440960
rect 291396 440552 291424 440932
rect 292224 440620 292252 441068
rect 293402 440988 293408 441040
rect 293460 440988 293466 441040
rect 293586 441028 293592 441040
rect 293512 441000 293592 441028
rect 292224 440592 292344 440620
rect 247972 440456 290964 440484
rect 291304 440524 291424 440552
rect 291304 440416 291332 440524
rect 240796 440388 291332 440416
rect 25498 440308 25504 440360
rect 25556 440348 25562 440360
rect 292316 440348 292344 440592
rect 293420 440416 293448 440988
rect 293512 440824 293540 441000
rect 293586 440988 293592 441000
rect 293644 440988 293650 441040
rect 293678 440988 293684 441040
rect 293736 440988 293742 441040
rect 293770 440988 293776 441040
rect 293828 440988 293834 441040
rect 293512 440796 293632 440824
rect 293604 440484 293632 440796
rect 293696 440552 293724 440988
rect 293788 440824 293816 440988
rect 299446 440960 299474 441068
rect 300826 441028 300854 441204
rect 302206 441096 302234 441340
rect 302206 441068 311894 441096
rect 303062 441028 303068 441040
rect 300826 441000 303068 441028
rect 303062 440988 303068 441000
rect 303120 440988 303126 441040
rect 304350 440988 304356 441040
rect 304408 440988 304414 441040
rect 299446 440932 302234 440960
rect 302206 440892 302234 440932
rect 304368 440892 304396 440988
rect 311866 440960 311894 441068
rect 580902 440960 580908 440972
rect 311866 440932 580908 440960
rect 580902 440920 580908 440932
rect 580960 440920 580966 440972
rect 580166 440892 580172 440904
rect 302206 440864 304396 440892
rect 309106 440864 580172 440892
rect 293788 440796 300854 440824
rect 300826 440620 300854 440796
rect 309106 440756 309134 440864
rect 580166 440852 580172 440864
rect 580224 440852 580230 440904
rect 307726 440728 309134 440756
rect 307726 440620 307754 440728
rect 300826 440592 307754 440620
rect 363598 440552 363604 440564
rect 293696 440524 363604 440552
rect 363598 440512 363604 440524
rect 363656 440512 363662 440564
rect 377398 440484 377404 440496
rect 293604 440456 377404 440484
rect 377398 440444 377404 440456
rect 377456 440444 377462 440496
rect 371970 440416 371976 440428
rect 293420 440388 300854 440416
rect 25556 440320 292344 440348
rect 300826 440348 300854 440388
rect 302206 440388 371976 440416
rect 302206 440348 302234 440388
rect 371970 440376 371976 440388
rect 372028 440376 372034 440428
rect 300826 440320 302234 440348
rect 25556 440308 25562 440320
rect 3326 423580 3332 423632
rect 3384 423620 3390 423632
rect 7558 423620 7564 423632
rect 3384 423592 7564 423620
rect 3384 423580 3390 423592
rect 7558 423580 7564 423592
rect 7616 423580 7622 423632
rect 363598 419432 363604 419484
rect 363656 419472 363662 419484
rect 579982 419472 579988 419484
rect 363656 419444 579988 419472
rect 363656 419432 363662 419444
rect 579982 419432 579988 419444
rect 580040 419432 580046 419484
rect 2958 411204 2964 411256
rect 3016 411244 3022 411256
rect 231210 411244 231216 411256
rect 3016 411216 231216 411244
rect 3016 411204 3022 411216
rect 231210 411204 231216 411216
rect 231268 411204 231274 411256
rect 362494 405628 362500 405680
rect 362552 405668 362558 405680
rect 579798 405668 579804 405680
rect 362552 405640 579804 405668
rect 362552 405628 362558 405640
rect 579798 405628 579804 405640
rect 579856 405628 579862 405680
rect 3050 398760 3056 398812
rect 3108 398800 3114 398812
rect 231118 398800 231124 398812
rect 3108 398772 231124 398800
rect 3108 398760 3114 398772
rect 231118 398760 231124 398772
rect 231176 398760 231182 398812
rect 362402 379448 362408 379500
rect 362460 379488 362466 379500
rect 580074 379488 580080 379500
rect 362460 379460 580080 379488
rect 362460 379448 362466 379460
rect 580074 379448 580080 379460
rect 580132 379448 580138 379500
rect 3786 378768 3792 378820
rect 3844 378808 3850 378820
rect 224218 378808 224224 378820
rect 3844 378780 224224 378808
rect 3844 378768 3850 378780
rect 224218 378768 224224 378780
rect 224276 378768 224282 378820
rect 97810 377408 97816 377460
rect 97868 377448 97874 377460
rect 229738 377448 229744 377460
rect 97868 377420 229744 377448
rect 97868 377408 97874 377420
rect 229738 377408 229744 377420
rect 229796 377408 229802 377460
rect 154758 374824 154764 374876
rect 154816 374864 154822 374876
rect 173158 374864 173164 374876
rect 154816 374836 173164 374864
rect 154816 374824 154822 374836
rect 173158 374824 173164 374836
rect 173216 374824 173222 374876
rect 110966 374756 110972 374808
rect 111024 374796 111030 374808
rect 228358 374796 228364 374808
rect 111024 374768 228364 374796
rect 111024 374756 111030 374768
rect 228358 374756 228364 374768
rect 228416 374756 228422 374808
rect 100662 374688 100668 374740
rect 100720 374728 100726 374740
rect 229830 374728 229836 374740
rect 100720 374700 229836 374728
rect 100720 374688 100726 374700
rect 229830 374688 229836 374700
rect 229888 374688 229894 374740
rect 126422 374620 126428 374672
rect 126480 374660 126486 374672
rect 170582 374660 170588 374672
rect 126480 374632 170588 374660
rect 126480 374620 126486 374632
rect 170582 374620 170588 374632
rect 170640 374620 170646 374672
rect 121270 374552 121276 374604
rect 121328 374592 121334 374604
rect 170950 374592 170956 374604
rect 121328 374564 170956 374592
rect 121328 374552 121334 374564
rect 170950 374552 170956 374564
rect 171008 374552 171014 374604
rect 165522 374484 165528 374536
rect 165580 374524 165586 374536
rect 227070 374524 227076 374536
rect 165580 374496 227076 374524
rect 165580 374484 165586 374496
rect 227070 374484 227076 374496
rect 227128 374484 227134 374536
rect 105814 374416 105820 374468
rect 105872 374456 105878 374468
rect 171778 374456 171784 374468
rect 105872 374428 171784 374456
rect 105872 374416 105878 374428
rect 171778 374416 171784 374428
rect 171836 374416 171842 374468
rect 157334 374348 157340 374400
rect 157392 374388 157398 374400
rect 228542 374388 228548 374400
rect 157392 374360 228548 374388
rect 157392 374348 157398 374360
rect 228542 374348 228548 374360
rect 228600 374348 228606 374400
rect 108390 374280 108396 374332
rect 108448 374320 108454 374332
rect 180058 374320 180064 374332
rect 108448 374292 180064 374320
rect 108448 374280 108454 374292
rect 180058 374280 180064 374292
rect 180116 374280 180122 374332
rect 152182 374212 152188 374264
rect 152240 374252 152246 374264
rect 231210 374252 231216 374264
rect 152240 374224 231216 374252
rect 152240 374212 152246 374224
rect 231210 374212 231216 374224
rect 231268 374212 231274 374264
rect 147030 374144 147036 374196
rect 147088 374184 147094 374196
rect 229738 374184 229744 374196
rect 147088 374156 229744 374184
rect 147088 374144 147094 374156
rect 229738 374144 229744 374156
rect 229796 374144 229802 374196
rect 139302 374008 139308 374060
rect 139360 374048 139366 374060
rect 155862 374048 155868 374060
rect 139360 374020 155868 374048
rect 139360 374008 139366 374020
rect 155862 374008 155868 374020
rect 155920 374008 155926 374060
rect 162486 374008 162492 374060
rect 162544 374048 162550 374060
rect 170398 374048 170404 374060
rect 162544 374020 170404 374048
rect 162544 374008 162550 374020
rect 170398 374008 170404 374020
rect 170456 374008 170462 374060
rect 32398 373124 32404 373176
rect 32456 373164 32462 373176
rect 165062 373164 165068 373176
rect 32456 373136 165068 373164
rect 32456 373124 32462 373136
rect 165062 373124 165068 373136
rect 165120 373164 165126 373176
rect 165522 373164 165528 373176
rect 165120 373136 165528 373164
rect 165120 373124 165126 373136
rect 165522 373124 165528 373136
rect 165580 373124 165586 373176
rect 123846 373056 123852 373108
rect 123904 373096 123910 373108
rect 174538 373096 174544 373108
rect 123904 373068 174544 373096
rect 123904 373056 123910 373068
rect 174538 373056 174544 373068
rect 174596 373056 174602 373108
rect 118694 372988 118700 373040
rect 118752 373028 118758 373040
rect 173250 373028 173256 373040
rect 118752 373000 173256 373028
rect 118752 372988 118758 373000
rect 173250 372988 173256 373000
rect 173308 372988 173314 373040
rect 103238 372920 103244 372972
rect 103296 372960 103302 372972
rect 173434 372960 173440 372972
rect 103296 372932 173440 372960
rect 103296 372920 103302 372932
rect 173434 372920 173440 372932
rect 173492 372920 173498 372972
rect 134150 372852 134156 372904
rect 134208 372892 134214 372904
rect 226978 372892 226984 372904
rect 134208 372864 226984 372892
rect 134208 372852 134214 372864
rect 226978 372852 226984 372864
rect 227036 372852 227042 372904
rect 131574 372784 131580 372836
rect 131632 372824 131638 372836
rect 231118 372824 231124 372836
rect 131632 372796 231124 372824
rect 131632 372784 131638 372796
rect 231118 372784 231124 372796
rect 231176 372784 231182 372836
rect 128998 372716 129004 372768
rect 129056 372756 129062 372768
rect 228450 372756 228456 372768
rect 129056 372728 228456 372756
rect 129056 372716 129062 372728
rect 228450 372716 228456 372728
rect 228508 372716 228514 372768
rect 113542 372648 113548 372700
rect 113600 372688 113606 372700
rect 229922 372688 229928 372700
rect 113600 372660 229928 372688
rect 113600 372648 113606 372660
rect 229922 372648 229928 372660
rect 229980 372648 229986 372700
rect 149606 372580 149612 372632
rect 149664 372620 149670 372632
rect 170490 372620 170496 372632
rect 149664 372592 170496 372620
rect 149664 372580 149670 372592
rect 170490 372580 170496 372592
rect 170548 372580 170554 372632
rect 3142 372512 3148 372564
rect 3200 372552 3206 372564
rect 100018 372552 100024 372564
rect 3200 372524 100024 372552
rect 3200 372512 3206 372524
rect 100018 372512 100024 372524
rect 100076 372512 100082 372564
rect 124766 371832 124772 371884
rect 124824 371872 124830 371884
rect 124824 371844 125824 371872
rect 124824 371832 124830 371844
rect 125686 371804 125692 371816
rect 118666 371776 125692 371804
rect 116394 371628 116400 371680
rect 116452 371668 116458 371680
rect 118666 371668 118694 371776
rect 125686 371764 125692 371776
rect 125744 371764 125750 371816
rect 125796 371804 125824 371844
rect 128262 371832 128268 371884
rect 128320 371872 128326 371884
rect 128320 371844 135254 371872
rect 128320 371832 128326 371844
rect 125796 371776 129734 371804
rect 128262 371736 128268 371748
rect 116452 371640 118694 371668
rect 123496 371708 128268 371736
rect 116452 371628 116458 371640
rect 97718 371560 97724 371612
rect 97776 371600 97782 371612
rect 123496 371600 123524 371708
rect 128262 371696 128268 371708
rect 128320 371696 128326 371748
rect 124876 371640 128400 371668
rect 97776 371572 123524 371600
rect 97776 371560 97782 371572
rect 124674 371560 124680 371612
rect 124732 371560 124738 371612
rect 124766 371560 124772 371612
rect 124824 371560 124830 371612
rect 97626 371492 97632 371544
rect 97684 371532 97690 371544
rect 124692 371532 124720 371560
rect 97684 371504 124720 371532
rect 97684 371492 97690 371504
rect 99834 371424 99840 371476
rect 99892 371464 99898 371476
rect 124784 371464 124812 371560
rect 99892 371436 124812 371464
rect 99892 371424 99898 371436
rect 97902 371356 97908 371408
rect 97960 371396 97966 371408
rect 97960 371368 118694 371396
rect 97960 371356 97966 371368
rect 118666 371260 118694 371368
rect 124876 371260 124904 371640
rect 125686 371560 125692 371612
rect 125744 371600 125750 371612
rect 125744 371572 125824 371600
rect 125744 371560 125750 371572
rect 118666 371232 124904 371260
rect 125796 371260 125824 371572
rect 128372 371464 128400 371640
rect 129706 371600 129734 371776
rect 135226 371736 135254 371844
rect 137002 371832 137008 371884
rect 137060 371872 137066 371884
rect 138474 371872 138480 371884
rect 137060 371844 138480 371872
rect 137060 371832 137066 371844
rect 138474 371832 138480 371844
rect 138532 371832 138538 371884
rect 138014 371764 138020 371816
rect 138072 371804 138078 371816
rect 143994 371804 144000 371816
rect 138072 371776 144000 371804
rect 138072 371764 138078 371776
rect 143994 371764 144000 371776
rect 144052 371764 144058 371816
rect 135226 371708 143764 371736
rect 143736 371668 143764 371708
rect 144012 371708 144224 371736
rect 144012 371668 144040 371708
rect 138400 371640 139394 371668
rect 143736 371640 144040 371668
rect 144196 371668 144224 371708
rect 167914 371696 167920 371748
rect 167972 371736 167978 371748
rect 170766 371736 170772 371748
rect 167972 371708 170772 371736
rect 167972 371696 167978 371708
rect 170766 371696 170772 371708
rect 170824 371696 170830 371748
rect 144196 371640 144408 371668
rect 129706 371572 132494 371600
rect 129844 371504 131068 371532
rect 128372 371436 129734 371464
rect 129706 371396 129734 371436
rect 129844 371396 129872 371504
rect 129706 371368 129872 371396
rect 131040 371328 131068 371504
rect 132466 371396 132494 371572
rect 135208 371560 135214 371612
rect 135266 371600 135272 371612
rect 137922 371600 137928 371612
rect 135266 371572 137928 371600
rect 135266 371560 135272 371572
rect 137922 371560 137928 371572
rect 137980 371560 137986 371612
rect 138014 371560 138020 371612
rect 138072 371560 138078 371612
rect 138032 371532 138060 371560
rect 136928 371504 138060 371532
rect 136928 371464 136956 371504
rect 135226 371436 136956 371464
rect 135226 371396 135254 371436
rect 138400 371396 138428 371640
rect 138474 371560 138480 371612
rect 138532 371560 138538 371612
rect 132466 371368 135254 371396
rect 137986 371368 138428 371396
rect 138492 371396 138520 371560
rect 139366 371464 139394 371640
rect 143994 371560 144000 371612
rect 144052 371560 144058 371612
rect 144178 371560 144184 371612
rect 144236 371560 144242 371612
rect 144380 371600 144408 371640
rect 144730 371628 144736 371680
rect 144788 371668 144794 371680
rect 174630 371668 174636 371680
rect 144788 371640 174636 371668
rect 144788 371628 144794 371640
rect 174630 371628 174636 371640
rect 174688 371628 174694 371680
rect 228634 371600 228640 371612
rect 144380 371572 228640 371600
rect 228634 371560 228640 371572
rect 228692 371560 228698 371612
rect 144012 371464 144040 371560
rect 144196 371532 144224 371560
rect 230014 371532 230020 371544
rect 144196 371504 230020 371532
rect 230014 371492 230020 371504
rect 230072 371492 230078 371544
rect 231302 371464 231308 371476
rect 139366 371436 139716 371464
rect 144012 371436 231308 371464
rect 138492 371368 138704 371396
rect 137986 371328 138014 371368
rect 131040 371300 138014 371328
rect 125796 371234 128308 371260
rect 138676 371234 138704 371368
rect 139688 371328 139716 371436
rect 231302 371424 231308 371436
rect 231360 371424 231366 371476
rect 231486 371396 231492 371408
rect 141528 371368 143534 371396
rect 141528 371328 141556 371368
rect 139688 371300 141556 371328
rect 125796 371232 128400 371234
rect 128280 371206 128400 371232
rect 128372 371124 128400 371206
rect 138492 371206 138704 371234
rect 131086 371164 132494 371192
rect 131086 371124 131114 371164
rect 128372 371096 131114 371124
rect 132466 371124 132494 371164
rect 133846 371164 135254 371192
rect 133846 371124 133874 371164
rect 132466 371096 133874 371124
rect 135226 371124 135254 371164
rect 135226 371096 136634 371124
rect 136606 370920 136634 371096
rect 138492 370988 138520 371206
rect 143506 371056 143534 371368
rect 144196 371368 231492 371396
rect 144196 371056 144224 371368
rect 231486 371356 231492 371368
rect 231544 371356 231550 371408
rect 231394 371328 231400 371340
rect 143506 371028 144224 371056
rect 144564 371300 231400 371328
rect 144564 370988 144592 371300
rect 231394 371288 231400 371300
rect 231452 371288 231458 371340
rect 231578 371260 231584 371272
rect 138492 370960 144592 370988
rect 144886 371232 231584 371260
rect 144886 370920 144914 371232
rect 231578 371220 231584 371232
rect 231636 371220 231642 371272
rect 136606 370892 144914 370920
rect 172330 368500 172336 368552
rect 172388 368540 172394 368552
rect 232222 368540 232228 368552
rect 172388 368512 232228 368540
rect 172388 368500 172394 368512
rect 232222 368500 232228 368512
rect 232280 368500 232286 368552
rect 169938 367888 169944 367940
rect 169996 367928 170002 367940
rect 170674 367928 170680 367940
rect 169996 367900 170680 367928
rect 169996 367888 170002 367900
rect 170674 367888 170680 367900
rect 170732 367888 170738 367940
rect 172422 365712 172428 365764
rect 172480 365752 172486 365764
rect 231670 365752 231676 365764
rect 172480 365724 231676 365752
rect 172480 365712 172486 365724
rect 231670 365712 231676 365724
rect 231728 365712 231734 365764
rect 378778 365644 378784 365696
rect 378836 365684 378842 365696
rect 580074 365684 580080 365696
rect 378836 365656 580080 365684
rect 378836 365644 378842 365656
rect 580074 365644 580080 365656
rect 580132 365644 580138 365696
rect 172330 362924 172336 362976
rect 172388 362964 172394 362976
rect 230106 362964 230112 362976
rect 172388 362936 230112 362964
rect 172388 362924 172394 362936
rect 230106 362924 230112 362936
rect 230164 362924 230170 362976
rect 171686 357416 171692 357468
rect 171744 357456 171750 357468
rect 228726 357456 228732 357468
rect 171744 357428 228732 357456
rect 171744 357416 171750 357428
rect 228726 357416 228732 357428
rect 228784 357416 228790 357468
rect 172422 351908 172428 351960
rect 172480 351948 172486 351960
rect 224218 351948 224224 351960
rect 172480 351920 224224 351948
rect 172480 351908 172486 351920
rect 224218 351908 224224 351920
rect 224276 351908 224282 351960
rect 172422 346400 172428 346452
rect 172480 346440 172486 346452
rect 220078 346440 220084 346452
rect 172480 346412 220084 346440
rect 172480 346400 172486 346412
rect 220078 346400 220084 346412
rect 220136 346400 220142 346452
rect 171134 345040 171140 345092
rect 171192 345080 171198 345092
rect 178678 345080 178684 345092
rect 171192 345052 178684 345080
rect 171192 345040 171198 345052
rect 178678 345040 178684 345052
rect 178736 345040 178742 345092
rect 172422 336744 172428 336796
rect 172480 336784 172486 336796
rect 225690 336784 225696 336796
rect 172480 336756 225696 336784
rect 172480 336744 172486 336756
rect 225690 336744 225696 336756
rect 225748 336744 225754 336796
rect 172422 333956 172428 334008
rect 172480 333996 172486 334008
rect 225782 333996 225788 334008
rect 172480 333968 225788 333996
rect 172480 333956 172486 333968
rect 225782 333956 225788 333968
rect 225840 333956 225846 334008
rect 172422 331236 172428 331288
rect 172480 331276 172486 331288
rect 230198 331276 230204 331288
rect 172480 331248 230204 331276
rect 172480 331236 172486 331248
rect 230198 331236 230204 331248
rect 230256 331236 230262 331288
rect 172422 325660 172428 325712
rect 172480 325700 172486 325712
rect 232222 325700 232228 325712
rect 172480 325672 232228 325700
rect 172480 325660 172486 325672
rect 232222 325660 232228 325672
rect 232280 325660 232286 325712
rect 362310 325592 362316 325644
rect 362368 325632 362374 325644
rect 580166 325632 580172 325644
rect 362368 325604 580172 325632
rect 362368 325592 362374 325604
rect 580166 325592 580172 325604
rect 580224 325592 580230 325644
rect 171318 322940 171324 322992
rect 171376 322980 171382 322992
rect 231762 322980 231768 322992
rect 171376 322952 231768 322980
rect 171376 322940 171382 322952
rect 231762 322940 231768 322952
rect 231820 322940 231826 322992
rect 171502 320152 171508 320204
rect 171560 320192 171566 320204
rect 231026 320192 231032 320204
rect 171560 320164 231032 320192
rect 171560 320152 171566 320164
rect 231026 320152 231032 320164
rect 231084 320152 231090 320204
rect 2958 320084 2964 320136
rect 3016 320124 3022 320136
rect 98638 320124 98644 320136
rect 3016 320096 98644 320124
rect 3016 320084 3022 320096
rect 98638 320084 98644 320096
rect 98696 320084 98702 320136
rect 171502 317432 171508 317484
rect 171560 317472 171566 317484
rect 231854 317472 231860 317484
rect 171560 317444 231860 317472
rect 171560 317432 171566 317444
rect 231854 317432 231860 317444
rect 231912 317432 231918 317484
rect 172422 314644 172428 314696
rect 172480 314684 172486 314696
rect 230382 314684 230388 314696
rect 172480 314656 230388 314684
rect 172480 314644 172486 314656
rect 230382 314644 230388 314656
rect 230440 314644 230446 314696
rect 377398 313216 377404 313268
rect 377456 313256 377462 313268
rect 580166 313256 580172 313268
rect 377456 313228 580172 313256
rect 377456 313216 377462 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 172422 311856 172428 311908
rect 172480 311896 172486 311908
rect 232038 311896 232044 311908
rect 172480 311868 232044 311896
rect 172480 311856 172486 311868
rect 232038 311856 232044 311868
rect 232096 311856 232102 311908
rect 172330 311380 172336 311432
rect 172388 311420 172394 311432
rect 230842 311420 230848 311432
rect 172388 311392 230848 311420
rect 172388 311380 172394 311392
rect 230842 311380 230848 311392
rect 230900 311380 230906 311432
rect 171870 311244 171876 311296
rect 171928 311284 171934 311296
rect 232222 311284 232228 311296
rect 171928 311256 232228 311284
rect 171928 311244 171934 311256
rect 232222 311244 232228 311256
rect 232280 311244 232286 311296
rect 172238 311176 172244 311228
rect 172296 311216 172302 311228
rect 230934 311216 230940 311228
rect 172296 311188 230940 311216
rect 172296 311176 172302 311188
rect 230934 311176 230940 311188
rect 230992 311176 230998 311228
rect 178678 311108 178684 311160
rect 178736 311148 178742 311160
rect 232222 311148 232228 311160
rect 178736 311120 232228 311148
rect 178736 311108 178742 311120
rect 232222 311108 232228 311120
rect 232280 311108 232286 311160
rect 230382 310700 230388 310752
rect 230440 310740 230446 310752
rect 230440 310712 232544 310740
rect 230440 310700 230446 310712
rect 172146 310564 172152 310616
rect 172204 310604 172210 310616
rect 230750 310604 230756 310616
rect 172204 310576 230756 310604
rect 172204 310564 172210 310576
rect 230750 310564 230756 310576
rect 230808 310564 230814 310616
rect 227070 310496 227076 310548
rect 227128 310536 227134 310548
rect 232516 310536 232544 310712
rect 235442 310536 235448 310548
rect 227128 310508 232268 310536
rect 232516 310508 235448 310536
rect 227128 310496 227134 310508
rect 232240 310468 232268 310508
rect 235442 310496 235448 310508
rect 235500 310496 235506 310548
rect 255406 310496 255412 310548
rect 255464 310536 255470 310548
rect 255590 310536 255596 310548
rect 255464 310508 255596 310536
rect 255464 310496 255470 310508
rect 255590 310496 255596 310508
rect 255648 310496 255654 310548
rect 273530 310496 273536 310548
rect 273588 310536 273594 310548
rect 273714 310536 273720 310548
rect 273588 310508 273720 310536
rect 273588 310496 273594 310508
rect 273714 310496 273720 310508
rect 273772 310496 273778 310548
rect 315022 310496 315028 310548
rect 315080 310536 315086 310548
rect 315390 310536 315396 310548
rect 315080 310508 315396 310536
rect 315080 310496 315086 310508
rect 315390 310496 315396 310508
rect 315448 310496 315454 310548
rect 232590 310468 232596 310480
rect 232240 310440 232596 310468
rect 232590 310428 232596 310440
rect 232648 310428 232654 310480
rect 231946 310360 231952 310412
rect 232004 310400 232010 310412
rect 232004 310372 238754 310400
rect 232004 310360 232010 310372
rect 230106 310292 230112 310344
rect 230164 310332 230170 310344
rect 233234 310332 233240 310344
rect 230164 310304 233240 310332
rect 230164 310292 230170 310304
rect 233234 310292 233240 310304
rect 233292 310292 233298 310344
rect 238726 310332 238754 310372
rect 244458 310332 244464 310344
rect 238726 310304 244464 310332
rect 244458 310292 244464 310304
rect 244516 310292 244522 310344
rect 230934 310224 230940 310276
rect 230992 310264 230998 310276
rect 231946 310264 231952 310276
rect 230992 310236 231952 310264
rect 230992 310224 230998 310236
rect 231946 310224 231952 310236
rect 232004 310224 232010 310276
rect 232038 310224 232044 310276
rect 232096 310264 232102 310276
rect 236270 310264 236276 310276
rect 232096 310236 236276 310264
rect 232096 310224 232102 310236
rect 236270 310224 236276 310236
rect 236328 310224 236334 310276
rect 231854 310156 231860 310208
rect 231912 310196 231918 310208
rect 241790 310196 241796 310208
rect 231912 310168 241796 310196
rect 231912 310156 231918 310168
rect 241790 310156 241796 310168
rect 241848 310156 241854 310208
rect 230842 310088 230848 310140
rect 230900 310128 230906 310140
rect 232038 310128 232044 310140
rect 230900 310100 232044 310128
rect 230900 310088 230906 310100
rect 232038 310088 232044 310100
rect 232096 310088 232102 310140
rect 171962 310020 171968 310072
rect 172020 310060 172026 310072
rect 237466 310060 237472 310072
rect 172020 310032 237472 310060
rect 172020 310020 172026 310032
rect 237466 310020 237472 310032
rect 237524 310020 237530 310072
rect 225690 309952 225696 310004
rect 225748 309992 225754 310004
rect 238938 309992 238944 310004
rect 225748 309964 238944 309992
rect 225748 309952 225754 309964
rect 238938 309952 238944 309964
rect 238996 309952 239002 310004
rect 286962 309952 286968 310004
rect 287020 309992 287026 310004
rect 287606 309992 287612 310004
rect 287020 309964 287612 309992
rect 287020 309952 287026 309964
rect 287606 309952 287612 309964
rect 287664 309952 287670 310004
rect 231762 309884 231768 309936
rect 231820 309924 231826 309936
rect 239490 309924 239496 309936
rect 231820 309896 239496 309924
rect 231820 309884 231826 309896
rect 239490 309884 239496 309896
rect 239548 309884 239554 309936
rect 230198 309748 230204 309800
rect 230256 309788 230262 309800
rect 241698 309788 241704 309800
rect 230256 309760 241704 309788
rect 230256 309748 230262 309760
rect 241698 309748 241704 309760
rect 241756 309748 241762 309800
rect 228726 309544 228732 309596
rect 228784 309584 228790 309596
rect 242986 309584 242992 309596
rect 228784 309556 242992 309584
rect 228784 309544 228790 309556
rect 242986 309544 242992 309556
rect 243044 309544 243050 309596
rect 232130 309476 232136 309528
rect 232188 309516 232194 309528
rect 249058 309516 249064 309528
rect 232188 309488 249064 309516
rect 232188 309476 232194 309488
rect 249058 309476 249064 309488
rect 249116 309476 249122 309528
rect 231670 309408 231676 309460
rect 231728 309448 231734 309460
rect 247494 309448 247500 309460
rect 231728 309420 247500 309448
rect 231728 309408 231734 309420
rect 247494 309408 247500 309420
rect 247552 309408 247558 309460
rect 241790 309340 241796 309392
rect 241848 309380 241854 309392
rect 249610 309380 249616 309392
rect 241848 309352 249616 309380
rect 241848 309340 241854 309352
rect 249610 309340 249616 309352
rect 249668 309340 249674 309392
rect 231026 309272 231032 309324
rect 231084 309312 231090 309324
rect 249794 309312 249800 309324
rect 231084 309284 249800 309312
rect 231084 309272 231090 309284
rect 249794 309272 249800 309284
rect 249852 309272 249858 309324
rect 170674 309204 170680 309256
rect 170732 309244 170738 309256
rect 234154 309244 234160 309256
rect 170732 309216 234160 309244
rect 170732 309204 170738 309216
rect 234154 309204 234160 309216
rect 234212 309204 234218 309256
rect 172238 309136 172244 309188
rect 172296 309176 172302 309188
rect 235902 309176 235908 309188
rect 172296 309148 235908 309176
rect 172296 309136 172302 309148
rect 235902 309136 235908 309148
rect 235960 309136 235966 309188
rect 237466 309136 237472 309188
rect 237524 309176 237530 309188
rect 237524 309148 238754 309176
rect 237524 309136 237530 309148
rect 238726 309120 238754 309148
rect 230014 309068 230020 309120
rect 230072 309108 230078 309120
rect 233602 309108 233608 309120
rect 230072 309080 233608 309108
rect 230072 309068 230078 309080
rect 233602 309068 233608 309080
rect 233660 309068 233666 309120
rect 234062 309068 234068 309120
rect 234120 309108 234126 309120
rect 238570 309108 238576 309120
rect 234120 309080 238576 309108
rect 234120 309068 234126 309080
rect 238570 309068 238576 309080
rect 238628 309068 238634 309120
rect 238726 309080 238760 309120
rect 238754 309068 238760 309080
rect 238812 309068 238818 309120
rect 347682 309068 347688 309120
rect 347740 309108 347746 309120
rect 347740 309080 351500 309108
rect 347740 309068 347746 309080
rect 229922 309000 229928 309052
rect 229980 309040 229986 309052
rect 235350 309040 235356 309052
rect 229980 309012 235356 309040
rect 229980 309000 229986 309012
rect 235350 309000 235356 309012
rect 235408 309000 235414 309052
rect 239766 309000 239772 309052
rect 239824 309040 239830 309052
rect 246758 309040 246764 309052
rect 239824 309012 246764 309040
rect 239824 309000 239830 309012
rect 246758 309000 246764 309012
rect 246816 309000 246822 309052
rect 326154 309000 326160 309052
rect 326212 309040 326218 309052
rect 340138 309040 340144 309052
rect 326212 309012 340144 309040
rect 326212 309000 326218 309012
rect 340138 309000 340144 309012
rect 340196 309000 340202 309052
rect 348970 309000 348976 309052
rect 349028 309040 349034 309052
rect 350902 309040 350908 309052
rect 349028 309012 350908 309040
rect 349028 309000 349034 309012
rect 350902 309000 350908 309012
rect 350960 309000 350966 309052
rect 231394 308932 231400 308984
rect 231452 308972 231458 308984
rect 237006 308972 237012 308984
rect 231452 308944 237012 308972
rect 231452 308932 231458 308944
rect 237006 308932 237012 308944
rect 237064 308932 237070 308984
rect 237098 308932 237104 308984
rect 237156 308972 237162 308984
rect 247126 308972 247132 308984
rect 237156 308944 247132 308972
rect 237156 308932 237162 308944
rect 247126 308932 247132 308944
rect 247184 308932 247190 308984
rect 310330 308932 310336 308984
rect 310388 308972 310394 308984
rect 310388 308944 311894 308972
rect 310388 308932 310394 308944
rect 230750 308864 230756 308916
rect 230808 308904 230814 308916
rect 252830 308904 252836 308916
rect 230808 308876 252836 308904
rect 230808 308864 230814 308876
rect 252830 308864 252836 308876
rect 252888 308864 252894 308916
rect 226978 308796 226984 308848
rect 227036 308836 227042 308848
rect 243354 308836 243360 308848
rect 227036 308808 243360 308836
rect 227036 308796 227042 308808
rect 243354 308796 243360 308808
rect 243412 308796 243418 308848
rect 251082 308796 251088 308848
rect 251140 308836 251146 308848
rect 257798 308836 257804 308848
rect 251140 308808 257804 308836
rect 251140 308796 251146 308808
rect 257798 308796 257804 308808
rect 257856 308796 257862 308848
rect 259546 308836 259552 308848
rect 257908 308808 259552 308836
rect 228450 308728 228456 308780
rect 228508 308768 228514 308780
rect 242158 308768 242164 308780
rect 228508 308740 242164 308768
rect 228508 308728 228514 308740
rect 242158 308728 242164 308740
rect 242216 308728 242222 308780
rect 247954 308728 247960 308780
rect 248012 308768 248018 308780
rect 254394 308768 254400 308780
rect 248012 308740 254400 308768
rect 248012 308728 248018 308740
rect 254394 308728 254400 308740
rect 254452 308728 254458 308780
rect 231118 308660 231124 308712
rect 231176 308700 231182 308712
rect 237098 308700 237104 308712
rect 231176 308672 237104 308700
rect 231176 308660 231182 308672
rect 237098 308660 237104 308672
rect 237156 308660 237162 308712
rect 237282 308660 237288 308712
rect 237340 308700 237346 308712
rect 241606 308700 241612 308712
rect 237340 308672 241612 308700
rect 237340 308660 237346 308672
rect 241606 308660 241612 308672
rect 241664 308660 241670 308712
rect 246298 308660 246304 308712
rect 246356 308700 246362 308712
rect 255958 308700 255964 308712
rect 246356 308672 255964 308700
rect 246356 308660 246362 308672
rect 255958 308660 255964 308672
rect 256016 308660 256022 308712
rect 170490 308592 170496 308644
rect 170548 308632 170554 308644
rect 239766 308632 239772 308644
rect 170548 308604 239772 308632
rect 170548 308592 170554 308604
rect 239766 308592 239772 308604
rect 239824 308592 239830 308644
rect 242342 308632 242348 308644
rect 239968 308604 242348 308632
rect 174538 308524 174544 308576
rect 174596 308564 174602 308576
rect 239968 308564 239996 308604
rect 242342 308592 242348 308604
rect 242400 308592 242406 308644
rect 250898 308592 250904 308644
rect 250956 308632 250962 308644
rect 257908 308632 257936 308808
rect 259546 308796 259552 308808
rect 259604 308796 259610 308848
rect 311866 308836 311894 308944
rect 333974 308932 333980 308984
rect 334032 308972 334038 308984
rect 334250 308972 334256 308984
rect 334032 308944 334256 308972
rect 334032 308932 334038 308944
rect 334250 308932 334256 308944
rect 334308 308932 334314 308984
rect 336734 308932 336740 308984
rect 336792 308972 336798 308984
rect 337378 308972 337384 308984
rect 336792 308944 337384 308972
rect 336792 308932 336798 308944
rect 337378 308932 337384 308944
rect 337436 308932 337442 308984
rect 350626 308932 350632 308984
rect 350684 308972 350690 308984
rect 351362 308972 351368 308984
rect 350684 308944 351368 308972
rect 350684 308932 350690 308944
rect 351362 308932 351368 308944
rect 351420 308932 351426 308984
rect 351472 308972 351500 309080
rect 354214 309068 354220 309120
rect 354272 309108 354278 309120
rect 367554 309108 367560 309120
rect 354272 309080 367560 309108
rect 354272 309068 354278 309080
rect 367554 309068 367560 309080
rect 367612 309068 367618 309120
rect 354582 309000 354588 309052
rect 354640 309040 354646 309052
rect 367830 309040 367836 309052
rect 354640 309012 367836 309040
rect 354640 309000 354646 309012
rect 367830 309000 367836 309012
rect 367888 309000 367894 309052
rect 366174 308972 366180 308984
rect 351472 308944 366180 308972
rect 366174 308932 366180 308944
rect 366232 308932 366238 308984
rect 312170 308864 312176 308916
rect 312228 308904 312234 308916
rect 355226 308904 355232 308916
rect 312228 308876 355232 308904
rect 312228 308864 312234 308876
rect 355226 308864 355232 308876
rect 355284 308864 355290 308916
rect 355318 308864 355324 308916
rect 355376 308904 355382 308916
rect 367370 308904 367376 308916
rect 355376 308876 367376 308904
rect 355376 308864 355382 308876
rect 367370 308864 367376 308876
rect 367428 308864 367434 308916
rect 356882 308836 356888 308848
rect 311866 308808 356888 308836
rect 356882 308796 356888 308808
rect 356940 308796 356946 308848
rect 358814 308796 358820 308848
rect 358872 308836 358878 308848
rect 359182 308836 359188 308848
rect 358872 308808 359188 308836
rect 358872 308796 358878 308808
rect 359182 308796 359188 308808
rect 359240 308796 359246 308848
rect 258166 308728 258172 308780
rect 258224 308768 258230 308780
rect 258810 308768 258816 308780
rect 258224 308740 258816 308768
rect 258224 308728 258230 308740
rect 258810 308728 258816 308740
rect 258868 308728 258874 308780
rect 267090 308728 267096 308780
rect 267148 308768 267154 308780
rect 281258 308768 281264 308780
rect 267148 308740 281264 308768
rect 267148 308728 267154 308740
rect 281258 308728 281264 308740
rect 281316 308728 281322 308780
rect 303798 308728 303804 308780
rect 303856 308768 303862 308780
rect 355594 308768 355600 308780
rect 303856 308740 355600 308768
rect 303856 308728 303862 308740
rect 355594 308728 355600 308740
rect 355652 308728 355658 308780
rect 356054 308728 356060 308780
rect 356112 308768 356118 308780
rect 363506 308768 363512 308780
rect 356112 308740 363512 308768
rect 356112 308728 356118 308740
rect 363506 308728 363512 308740
rect 363564 308728 363570 308780
rect 267182 308700 267188 308712
rect 250956 308604 257936 308632
rect 258736 308672 267188 308700
rect 250956 308592 250962 308604
rect 241974 308564 241980 308576
rect 174596 308536 239996 308564
rect 240060 308536 241980 308564
rect 174596 308524 174602 308536
rect 232406 308456 232412 308508
rect 232464 308496 232470 308508
rect 237282 308496 237288 308508
rect 232464 308468 237288 308496
rect 232464 308456 232470 308468
rect 237282 308456 237288 308468
rect 237340 308456 237346 308508
rect 237926 308456 237932 308508
rect 237984 308496 237990 308508
rect 240060 308496 240088 308536
rect 241974 308524 241980 308536
rect 242032 308524 242038 308576
rect 242802 308524 242808 308576
rect 242860 308564 242866 308576
rect 252462 308564 252468 308576
rect 242860 308536 252468 308564
rect 242860 308524 242866 308536
rect 252462 308524 252468 308536
rect 252520 308524 252526 308576
rect 253198 308524 253204 308576
rect 253256 308564 253262 308576
rect 258736 308564 258764 308672
rect 267182 308660 267188 308672
rect 267240 308660 267246 308712
rect 287238 308660 287244 308712
rect 287296 308700 287302 308712
rect 287514 308700 287520 308712
rect 287296 308672 287520 308700
rect 287296 308660 287302 308672
rect 287514 308660 287520 308672
rect 287572 308660 287578 308712
rect 302694 308660 302700 308712
rect 302752 308700 302758 308712
rect 355410 308700 355416 308712
rect 302752 308672 355416 308700
rect 302752 308660 302758 308672
rect 355410 308660 355416 308672
rect 355468 308660 355474 308712
rect 356514 308660 356520 308712
rect 356572 308700 356578 308712
rect 367278 308700 367284 308712
rect 356572 308672 367284 308700
rect 356572 308660 356578 308672
rect 367278 308660 367284 308672
rect 367336 308660 367342 308712
rect 260558 308592 260564 308644
rect 260616 308632 260622 308644
rect 268746 308632 268752 308644
rect 260616 308604 268752 308632
rect 260616 308592 260622 308604
rect 268746 308592 268752 308604
rect 268804 308592 268810 308644
rect 287146 308592 287152 308644
rect 287204 308632 287210 308644
rect 287204 308604 287376 308632
rect 287204 308592 287210 308604
rect 253256 308536 258764 308564
rect 253256 308524 253262 308536
rect 258810 308524 258816 308576
rect 258868 308564 258874 308576
rect 271598 308564 271604 308576
rect 258868 308536 271604 308564
rect 258868 308524 258874 308536
rect 271598 308524 271604 308536
rect 271656 308524 271662 308576
rect 237984 308468 240088 308496
rect 237984 308456 237990 308468
rect 240134 308456 240140 308508
rect 240192 308496 240198 308508
rect 241054 308496 241060 308508
rect 240192 308468 241060 308496
rect 240192 308456 240198 308468
rect 241054 308456 241060 308468
rect 241112 308456 241118 308508
rect 271138 308456 271144 308508
rect 271196 308496 271202 308508
rect 273438 308496 273444 308508
rect 271196 308468 273444 308496
rect 271196 308456 271202 308468
rect 273438 308456 273444 308468
rect 273496 308456 273502 308508
rect 236178 308388 236184 308440
rect 236236 308428 236242 308440
rect 236822 308428 236828 308440
rect 236236 308400 236828 308428
rect 236236 308388 236242 308400
rect 236822 308388 236828 308400
rect 236880 308388 236886 308440
rect 238846 308388 238852 308440
rect 238904 308428 238910 308440
rect 239306 308428 239312 308440
rect 238904 308400 239312 308428
rect 238904 308388 238910 308400
rect 239306 308388 239312 308400
rect 239364 308388 239370 308440
rect 240226 308388 240232 308440
rect 240284 308428 240290 308440
rect 240686 308428 240692 308440
rect 240284 308400 240692 308428
rect 240284 308388 240290 308400
rect 240686 308388 240692 308400
rect 240744 308388 240750 308440
rect 242986 308388 242992 308440
rect 243044 308428 243050 308440
rect 243538 308428 243544 308440
rect 243044 308400 243544 308428
rect 243044 308388 243050 308400
rect 243538 308388 243544 308400
rect 243596 308388 243602 308440
rect 272702 308428 272708 308440
rect 253906 308400 272708 308428
rect 174630 308320 174636 308372
rect 174688 308360 174694 308372
rect 238202 308360 238208 308372
rect 174688 308332 238208 308360
rect 174688 308320 174694 308332
rect 238202 308320 238208 308332
rect 238260 308320 238266 308372
rect 238938 308320 238944 308372
rect 238996 308360 239002 308372
rect 239858 308360 239864 308372
rect 238996 308332 239864 308360
rect 238996 308320 239002 308332
rect 239858 308320 239864 308332
rect 239916 308320 239922 308372
rect 240318 308320 240324 308372
rect 240376 308360 240382 308372
rect 240870 308360 240876 308372
rect 240376 308332 240876 308360
rect 240376 308320 240382 308332
rect 240870 308320 240876 308332
rect 240928 308320 240934 308372
rect 246390 308360 246396 308372
rect 242544 308332 246396 308360
rect 236086 308252 236092 308304
rect 236144 308292 236150 308304
rect 236362 308292 236368 308304
rect 236144 308264 236368 308292
rect 236144 308252 236150 308264
rect 236362 308252 236368 308264
rect 236420 308252 236426 308304
rect 237558 308252 237564 308304
rect 237616 308292 237622 308304
rect 237834 308292 237840 308304
rect 237616 308264 237840 308292
rect 237616 308252 237622 308264
rect 237834 308252 237840 308264
rect 237892 308252 237898 308304
rect 242544 308292 242572 308332
rect 246390 308320 246396 308332
rect 246448 308320 246454 308372
rect 237944 308264 242572 308292
rect 231578 308184 231584 308236
rect 231636 308224 231642 308236
rect 237944 308224 237972 308264
rect 243170 308252 243176 308304
rect 243228 308292 243234 308304
rect 244090 308292 244096 308304
rect 243228 308264 244096 308292
rect 243228 308252 243234 308264
rect 244090 308252 244096 308264
rect 244148 308252 244154 308304
rect 231636 308196 237972 308224
rect 231636 308184 231642 308196
rect 236086 308116 236092 308168
rect 236144 308156 236150 308168
rect 236638 308156 236644 308168
rect 236144 308128 236644 308156
rect 236144 308116 236150 308128
rect 236638 308116 236644 308128
rect 236696 308116 236702 308168
rect 232038 308048 232044 308100
rect 232096 308088 232102 308100
rect 237926 308088 237932 308100
rect 232096 308060 237932 308088
rect 232096 308048 232102 308060
rect 237926 308048 237932 308060
rect 237984 308048 237990 308100
rect 231946 307980 231952 308032
rect 232004 308020 232010 308032
rect 245838 308020 245844 308032
rect 232004 307992 245844 308020
rect 232004 307980 232010 307992
rect 245838 307980 245844 307992
rect 245896 307980 245902 308032
rect 251082 307952 251088 307964
rect 250456 307924 251088 307952
rect 250456 307896 250484 307924
rect 251082 307912 251088 307924
rect 251140 307912 251146 307964
rect 252186 307912 252192 307964
rect 252244 307952 252250 307964
rect 253906 307952 253934 308400
rect 272702 308388 272708 308400
rect 272760 308388 272766 308440
rect 284294 308388 284300 308440
rect 284352 308428 284358 308440
rect 285122 308428 285128 308440
rect 284352 308400 285128 308428
rect 284352 308388 284358 308400
rect 285122 308388 285128 308400
rect 285180 308388 285186 308440
rect 286134 308388 286140 308440
rect 286192 308428 286198 308440
rect 286410 308428 286416 308440
rect 286192 308400 286416 308428
rect 286192 308388 286198 308400
rect 286410 308388 286416 308400
rect 286468 308388 286474 308440
rect 287348 308304 287376 308604
rect 288526 308592 288532 308644
rect 288584 308592 288590 308644
rect 302326 308592 302332 308644
rect 302384 308632 302390 308644
rect 355686 308632 355692 308644
rect 302384 308604 355692 308632
rect 302384 308592 302390 308604
rect 355686 308592 355692 308604
rect 355744 308592 355750 308644
rect 356974 308592 356980 308644
rect 357032 308632 357038 308644
rect 369946 308632 369952 308644
rect 357032 308604 369952 308632
rect 357032 308592 357038 308604
rect 369946 308592 369952 308604
rect 370004 308592 370010 308644
rect 287790 308496 287796 308508
rect 287440 308468 287796 308496
rect 287440 308304 287468 308468
rect 287790 308456 287796 308468
rect 287848 308456 287854 308508
rect 287974 308456 287980 308508
rect 288032 308456 288038 308508
rect 287330 308252 287336 308304
rect 287388 308252 287394 308304
rect 287422 308252 287428 308304
rect 287480 308252 287486 308304
rect 287238 308184 287244 308236
rect 287296 308224 287302 308236
rect 287992 308224 288020 308456
rect 288544 308372 288572 308592
rect 301682 308524 301688 308576
rect 301740 308564 301746 308576
rect 355042 308564 355048 308576
rect 301740 308536 355048 308564
rect 301740 308524 301746 308536
rect 355042 308524 355048 308536
rect 355100 308524 355106 308576
rect 357250 308524 357256 308576
rect 357308 308564 357314 308576
rect 370498 308564 370504 308576
rect 357308 308536 370504 308564
rect 357308 308524 357314 308536
rect 370498 308524 370504 308536
rect 370556 308524 370562 308576
rect 289814 308456 289820 308508
rect 289872 308496 289878 308508
rect 290274 308496 290280 308508
rect 289872 308468 290280 308496
rect 289872 308456 289878 308468
rect 290274 308456 290280 308468
rect 290332 308456 290338 308508
rect 291286 308456 291292 308508
rect 291344 308496 291350 308508
rect 291654 308496 291660 308508
rect 291344 308468 291660 308496
rect 291344 308456 291350 308468
rect 291654 308456 291660 308468
rect 291712 308456 291718 308508
rect 300762 308456 300768 308508
rect 300820 308496 300826 308508
rect 356790 308496 356796 308508
rect 300820 308468 356796 308496
rect 300820 308456 300826 308468
rect 356790 308456 356796 308468
rect 356848 308456 356854 308508
rect 288802 308388 288808 308440
rect 288860 308428 288866 308440
rect 289722 308428 289728 308440
rect 288860 308400 289728 308428
rect 288860 308388 288866 308400
rect 289722 308388 289728 308400
rect 289780 308388 289786 308440
rect 291470 308388 291476 308440
rect 291528 308428 291534 308440
rect 292390 308428 292396 308440
rect 291528 308400 292396 308428
rect 291528 308388 291534 308400
rect 292390 308388 292396 308400
rect 292448 308388 292454 308440
rect 299658 308388 299664 308440
rect 299716 308428 299722 308440
rect 354674 308428 354680 308440
rect 299716 308400 354680 308428
rect 299716 308388 299722 308400
rect 354674 308388 354680 308400
rect 354732 308388 354738 308440
rect 354858 308388 354864 308440
rect 354916 308428 354922 308440
rect 355870 308428 355876 308440
rect 354916 308400 355876 308428
rect 354916 308388 354922 308400
rect 355870 308388 355876 308400
rect 355928 308388 355934 308440
rect 359274 308388 359280 308440
rect 359332 308428 359338 308440
rect 359918 308428 359924 308440
rect 359332 308400 359924 308428
rect 359332 308388 359338 308400
rect 359918 308388 359924 308400
rect 359976 308388 359982 308440
rect 288526 308320 288532 308372
rect 288584 308320 288590 308372
rect 291654 308320 291660 308372
rect 291712 308360 291718 308372
rect 292206 308360 292212 308372
rect 291712 308332 292212 308360
rect 291712 308320 291718 308332
rect 292206 308320 292212 308332
rect 292264 308320 292270 308372
rect 331214 308320 331220 308372
rect 331272 308360 331278 308372
rect 332226 308360 332232 308372
rect 331272 308332 332232 308360
rect 331272 308320 331278 308332
rect 332226 308320 332232 308332
rect 332284 308320 332290 308372
rect 333054 308320 333060 308372
rect 333112 308360 333118 308372
rect 333606 308360 333612 308372
rect 333112 308332 333612 308360
rect 333112 308320 333118 308332
rect 333606 308320 333612 308332
rect 333664 308320 333670 308372
rect 334434 308320 334440 308372
rect 334492 308360 334498 308372
rect 334894 308360 334900 308372
rect 334492 308332 334900 308360
rect 334492 308320 334498 308332
rect 334894 308320 334900 308332
rect 334952 308320 334958 308372
rect 335814 308320 335820 308372
rect 335872 308360 335878 308372
rect 336458 308360 336464 308372
rect 335872 308332 336464 308360
rect 335872 308320 335878 308332
rect 336458 308320 336464 308332
rect 336516 308320 336522 308372
rect 338482 308320 338488 308372
rect 338540 308360 338546 308372
rect 339310 308360 339316 308372
rect 338540 308332 339316 308360
rect 338540 308320 338546 308332
rect 339310 308320 339316 308332
rect 339368 308320 339374 308372
rect 352098 308320 352104 308372
rect 352156 308360 352162 308372
rect 352466 308360 352472 308372
rect 352156 308332 352472 308360
rect 352156 308320 352162 308332
rect 352466 308320 352472 308332
rect 352524 308320 352530 308372
rect 353386 308320 353392 308372
rect 353444 308360 353450 308372
rect 354030 308360 354036 308372
rect 353444 308332 354036 308360
rect 353444 308320 353450 308332
rect 354030 308320 354036 308332
rect 354088 308320 354094 308372
rect 367646 308360 367652 308372
rect 354508 308332 367652 308360
rect 288618 308252 288624 308304
rect 288676 308292 288682 308304
rect 289078 308292 289084 308304
rect 288676 308264 289084 308292
rect 288676 308252 288682 308264
rect 289078 308252 289084 308264
rect 289136 308252 289142 308304
rect 290274 308252 290280 308304
rect 290332 308292 290338 308304
rect 291010 308292 291016 308304
rect 290332 308264 291016 308292
rect 290332 308252 290338 308264
rect 291010 308252 291016 308264
rect 291068 308252 291074 308304
rect 291194 308252 291200 308304
rect 291252 308292 291258 308304
rect 291746 308292 291752 308304
rect 291252 308264 291752 308292
rect 291252 308252 291258 308264
rect 291746 308252 291752 308264
rect 291804 308252 291810 308304
rect 331306 308252 331312 308304
rect 331364 308292 331370 308304
rect 331766 308292 331772 308304
rect 331364 308264 331772 308292
rect 331364 308252 331370 308264
rect 331766 308252 331772 308264
rect 331824 308252 331830 308304
rect 332686 308252 332692 308304
rect 332744 308292 332750 308304
rect 333422 308292 333428 308304
rect 332744 308264 333428 308292
rect 332744 308252 332750 308264
rect 333422 308252 333428 308264
rect 333480 308252 333486 308304
rect 334526 308252 334532 308304
rect 334584 308292 334590 308304
rect 335078 308292 335084 308304
rect 334584 308264 335084 308292
rect 334584 308252 334590 308264
rect 335078 308252 335084 308264
rect 335136 308252 335142 308304
rect 335538 308252 335544 308304
rect 335596 308292 335602 308304
rect 336274 308292 336280 308304
rect 335596 308264 336280 308292
rect 335596 308252 335602 308264
rect 336274 308252 336280 308264
rect 336332 308252 336338 308304
rect 336826 308252 336832 308304
rect 336884 308292 336890 308304
rect 337102 308292 337108 308304
rect 336884 308264 337108 308292
rect 336884 308252 336890 308264
rect 337102 308252 337108 308264
rect 337160 308252 337166 308304
rect 338206 308252 338212 308304
rect 338264 308292 338270 308304
rect 338666 308292 338672 308304
rect 338264 308264 338672 308292
rect 338264 308252 338270 308264
rect 338666 308252 338672 308264
rect 338724 308252 338730 308304
rect 339862 308252 339868 308304
rect 339920 308292 339926 308304
rect 340230 308292 340236 308304
rect 339920 308264 340236 308292
rect 339920 308252 339926 308264
rect 340230 308252 340236 308264
rect 340288 308252 340294 308304
rect 350534 308252 350540 308304
rect 350592 308292 350598 308304
rect 350994 308292 351000 308304
rect 350592 308264 351000 308292
rect 350592 308252 350598 308264
rect 350994 308252 351000 308264
rect 351052 308252 351058 308304
rect 351178 308252 351184 308304
rect 351236 308292 351242 308304
rect 352006 308292 352012 308304
rect 351236 308264 352012 308292
rect 351236 308252 351242 308264
rect 352006 308252 352012 308264
rect 352064 308252 352070 308304
rect 352190 308252 352196 308304
rect 352248 308292 352254 308304
rect 352650 308292 352656 308304
rect 352248 308264 352656 308292
rect 352248 308252 352254 308264
rect 352650 308252 352656 308264
rect 352708 308252 352714 308304
rect 353294 308252 353300 308304
rect 353352 308292 353358 308304
rect 354398 308292 354404 308304
rect 353352 308264 354404 308292
rect 353352 308252 353358 308264
rect 354398 308252 354404 308264
rect 354456 308252 354462 308304
rect 287296 308196 288020 308224
rect 287296 308184 287302 308196
rect 288710 308184 288716 308236
rect 288768 308224 288774 308236
rect 289538 308224 289544 308236
rect 288768 308196 289544 308224
rect 288768 308184 288774 308196
rect 289538 308184 289544 308196
rect 289596 308184 289602 308236
rect 332594 308184 332600 308236
rect 332652 308224 332658 308236
rect 333790 308224 333796 308236
rect 332652 308196 333796 308224
rect 332652 308184 332658 308196
rect 333790 308184 333796 308196
rect 333848 308184 333854 308236
rect 334066 308184 334072 308236
rect 334124 308224 334130 308236
rect 334710 308224 334716 308236
rect 334124 308196 334716 308224
rect 334124 308184 334130 308196
rect 334710 308184 334716 308196
rect 334768 308184 334774 308236
rect 335354 308184 335360 308236
rect 335412 308224 335418 308236
rect 336090 308224 336096 308236
rect 335412 308196 336096 308224
rect 335412 308184 335418 308196
rect 336090 308184 336096 308196
rect 336148 308184 336154 308236
rect 338114 308184 338120 308236
rect 338172 308224 338178 308236
rect 338942 308224 338948 308236
rect 338172 308196 338948 308224
rect 338172 308184 338178 308196
rect 338942 308184 338948 308196
rect 339000 308184 339006 308236
rect 339678 308184 339684 308236
rect 339736 308224 339742 308236
rect 340046 308224 340052 308236
rect 339736 308196 340052 308224
rect 339736 308184 339742 308196
rect 340046 308184 340052 308196
rect 340104 308184 340110 308236
rect 350902 308184 350908 308236
rect 350960 308224 350966 308236
rect 351730 308224 351736 308236
rect 350960 308196 351736 308224
rect 350960 308184 350966 308196
rect 351730 308184 351736 308196
rect 351788 308184 351794 308236
rect 352834 308224 352840 308236
rect 352024 308196 352840 308224
rect 352024 308168 352052 308196
rect 352834 308184 352840 308196
rect 352892 308184 352898 308236
rect 353018 308184 353024 308236
rect 353076 308184 353082 308236
rect 353846 308184 353852 308236
rect 353904 308224 353910 308236
rect 354508 308224 354536 308332
rect 367646 308320 367652 308332
rect 367704 308320 367710 308372
rect 365070 308292 365076 308304
rect 353904 308196 354536 308224
rect 354646 308264 365076 308292
rect 353904 308184 353910 308196
rect 284662 308116 284668 308168
rect 284720 308156 284726 308168
rect 285490 308156 285496 308168
rect 284720 308128 285496 308156
rect 284720 308116 284726 308128
rect 285490 308116 285496 308128
rect 285548 308116 285554 308168
rect 285858 308116 285864 308168
rect 285916 308156 285922 308168
rect 286042 308156 286048 308168
rect 285916 308128 286048 308156
rect 285916 308116 285922 308128
rect 286042 308116 286048 308128
rect 286100 308116 286106 308168
rect 291194 308116 291200 308168
rect 291252 308156 291258 308168
rect 292022 308156 292028 308168
rect 291252 308128 292028 308156
rect 291252 308116 291258 308128
rect 292022 308116 292028 308128
rect 292080 308116 292086 308168
rect 331306 308116 331312 308168
rect 331364 308156 331370 308168
rect 332042 308156 332048 308168
rect 331364 308128 332048 308156
rect 331364 308116 331370 308128
rect 332042 308116 332048 308128
rect 332100 308116 332106 308168
rect 332502 308116 332508 308168
rect 332560 308156 332566 308168
rect 332870 308156 332876 308168
rect 332560 308128 332876 308156
rect 332560 308116 332566 308128
rect 332870 308116 332876 308128
rect 332928 308116 332934 308168
rect 334158 308116 334164 308168
rect 334216 308156 334222 308168
rect 335262 308156 335268 308168
rect 334216 308128 335268 308156
rect 334216 308116 334222 308128
rect 335262 308116 335268 308128
rect 335320 308116 335326 308168
rect 335446 308116 335452 308168
rect 335504 308156 335510 308168
rect 336642 308156 336648 308168
rect 335504 308128 336648 308156
rect 335504 308116 335510 308128
rect 336642 308116 336648 308128
rect 336700 308116 336706 308168
rect 336918 308116 336924 308168
rect 336976 308156 336982 308168
rect 337286 308156 337292 308168
rect 336976 308128 337292 308156
rect 336976 308116 336982 308128
rect 337286 308116 337292 308128
rect 337344 308116 337350 308168
rect 338206 308116 338212 308168
rect 338264 308156 338270 308168
rect 339126 308156 339132 308168
rect 338264 308128 339132 308156
rect 338264 308116 338270 308128
rect 339126 308116 339132 308128
rect 339184 308116 339190 308168
rect 352006 308116 352012 308168
rect 352064 308116 352070 308168
rect 353036 308156 353064 308184
rect 354646 308156 354674 308264
rect 365070 308252 365076 308264
rect 365128 308252 365134 308304
rect 357342 308184 357348 308236
rect 357400 308224 357406 308236
rect 357802 308224 357808 308236
rect 357400 308196 357808 308224
rect 357400 308184 357406 308196
rect 357802 308184 357808 308196
rect 357860 308184 357866 308236
rect 359090 308184 359096 308236
rect 359148 308224 359154 308236
rect 359734 308224 359740 308236
rect 359148 308196 359740 308224
rect 359148 308184 359154 308196
rect 359734 308184 359740 308196
rect 359792 308184 359798 308236
rect 353036 308128 354674 308156
rect 355778 308116 355784 308168
rect 355836 308156 355842 308168
rect 355836 308128 359136 308156
rect 355836 308116 355842 308128
rect 284754 308048 284760 308100
rect 284812 308088 284818 308100
rect 285306 308088 285312 308100
rect 284812 308060 285312 308088
rect 284812 308048 284818 308060
rect 285306 308048 285312 308060
rect 285364 308048 285370 308100
rect 354674 308048 354680 308100
rect 354732 308088 354738 308100
rect 356974 308088 356980 308100
rect 354732 308060 356980 308088
rect 354732 308048 354738 308060
rect 356974 308048 356980 308060
rect 357032 308048 357038 308100
rect 357618 308048 357624 308100
rect 357676 308088 357682 308100
rect 357986 308088 357992 308100
rect 357676 308060 357992 308088
rect 357676 308048 357682 308060
rect 357986 308048 357992 308060
rect 358044 308048 358050 308100
rect 359108 308088 359136 308128
rect 359182 308116 359188 308168
rect 359240 308156 359246 308168
rect 360102 308156 360108 308168
rect 359240 308128 360108 308156
rect 359240 308116 359246 308128
rect 360102 308116 360108 308128
rect 360160 308116 360166 308168
rect 366358 308088 366364 308100
rect 359108 308060 366364 308088
rect 366358 308048 366364 308060
rect 366416 308048 366422 308100
rect 351914 307980 351920 308032
rect 351972 308020 351978 308032
rect 352558 308020 352564 308032
rect 351972 307992 352564 308020
rect 351972 307980 351978 307992
rect 352558 307980 352564 307992
rect 352616 307980 352622 308032
rect 353478 307980 353484 308032
rect 353536 308020 353542 308032
rect 364886 308020 364892 308032
rect 353536 307992 364892 308020
rect 353536 307980 353542 307992
rect 364886 307980 364892 307992
rect 364944 307980 364950 308032
rect 252244 307924 253934 307952
rect 252244 307912 252250 307924
rect 256234 307912 256240 307964
rect 256292 307952 256298 307964
rect 262398 307952 262404 307964
rect 256292 307924 262404 307952
rect 256292 307912 256298 307924
rect 262398 307912 262404 307924
rect 262456 307912 262462 307964
rect 356698 307912 356704 307964
rect 356756 307952 356762 307964
rect 359550 307952 359556 307964
rect 356756 307924 359556 307952
rect 356756 307912 356762 307924
rect 359550 307912 359556 307924
rect 359608 307912 359614 307964
rect 250438 307844 250444 307896
rect 250496 307844 250502 307896
rect 250530 307844 250536 307896
rect 250588 307884 250594 307896
rect 250898 307884 250904 307896
rect 250588 307856 250904 307884
rect 250588 307844 250594 307856
rect 250898 307844 250904 307856
rect 250956 307844 250962 307896
rect 252002 307844 252008 307896
rect 252060 307884 252066 307896
rect 258810 307884 258816 307896
rect 252060 307856 258816 307884
rect 252060 307844 252066 307856
rect 258810 307844 258816 307856
rect 258868 307844 258874 307896
rect 261754 307844 261760 307896
rect 261812 307884 261818 307896
rect 269850 307884 269856 307896
rect 261812 307856 269856 307884
rect 261812 307844 261818 307856
rect 269850 307844 269856 307856
rect 269908 307844 269914 307896
rect 282914 307844 282920 307896
rect 282972 307884 282978 307896
rect 283282 307884 283288 307896
rect 282972 307856 283288 307884
rect 282972 307844 282978 307856
rect 283282 307844 283288 307856
rect 283340 307844 283346 307896
rect 283374 307844 283380 307896
rect 283432 307884 283438 307896
rect 284018 307884 284024 307896
rect 283432 307856 284024 307884
rect 283432 307844 283438 307856
rect 284018 307844 284024 307856
rect 284076 307844 284082 307896
rect 285674 307844 285680 307896
rect 285732 307884 285738 307896
rect 285950 307884 285956 307896
rect 285732 307856 285956 307884
rect 285732 307844 285738 307856
rect 285950 307844 285956 307856
rect 286008 307844 286014 307896
rect 289814 307844 289820 307896
rect 289872 307884 289878 307896
rect 290642 307884 290648 307896
rect 289872 307856 290648 307884
rect 289872 307844 289878 307856
rect 290642 307844 290648 307856
rect 290700 307844 290706 307896
rect 336918 307844 336924 307896
rect 336976 307884 336982 307896
rect 337746 307884 337752 307896
rect 336976 307856 337752 307884
rect 336976 307844 336982 307856
rect 337746 307844 337752 307856
rect 337804 307844 337810 307896
rect 354950 307844 354956 307896
rect 355008 307884 355014 307896
rect 367462 307884 367468 307896
rect 355008 307856 367468 307884
rect 355008 307844 355014 307856
rect 367462 307844 367468 307856
rect 367520 307844 367526 307896
rect 247770 307776 247776 307828
rect 247828 307816 247834 307828
rect 248506 307816 248512 307828
rect 247828 307788 248512 307816
rect 247828 307776 247834 307788
rect 248506 307776 248512 307788
rect 248564 307776 248570 307828
rect 250622 307776 250628 307828
rect 250680 307816 250686 307828
rect 251358 307816 251364 307828
rect 250680 307788 251364 307816
rect 250680 307776 250686 307788
rect 251358 307776 251364 307788
rect 251416 307776 251422 307828
rect 257706 307776 257712 307828
rect 257764 307816 257770 307828
rect 258994 307816 259000 307828
rect 257764 307788 259000 307816
rect 257764 307776 257770 307788
rect 258994 307776 259000 307788
rect 259052 307776 259058 307828
rect 264422 307776 264428 307828
rect 264480 307816 264486 307828
rect 266998 307816 267004 307828
rect 264480 307788 267004 307816
rect 264480 307776 264486 307788
rect 266998 307776 267004 307788
rect 267056 307776 267062 307828
rect 284386 307776 284392 307828
rect 284444 307816 284450 307828
rect 284846 307816 284852 307828
rect 284444 307788 284852 307816
rect 284444 307776 284450 307788
rect 284846 307776 284852 307788
rect 284904 307776 284910 307828
rect 285858 307776 285864 307828
rect 285916 307816 285922 307828
rect 286870 307816 286876 307828
rect 285916 307788 286876 307816
rect 285916 307776 285922 307788
rect 286870 307776 286876 307788
rect 286928 307776 286934 307828
rect 317322 307776 317328 307828
rect 317380 307816 317386 307828
rect 318058 307816 318064 307828
rect 317380 307788 318064 307816
rect 317380 307776 317386 307788
rect 318058 307776 318064 307788
rect 318116 307776 318122 307828
rect 336826 307776 336832 307828
rect 336884 307816 336890 307828
rect 337930 307816 337936 307828
rect 336884 307788 337936 307816
rect 336884 307776 336890 307788
rect 337930 307776 337936 307788
rect 337988 307776 337994 307828
rect 348418 307776 348424 307828
rect 348476 307816 348482 307828
rect 350350 307816 350356 307828
rect 348476 307788 350356 307816
rect 348476 307776 348482 307788
rect 350350 307776 350356 307788
rect 350408 307776 350414 307828
rect 228358 307708 228364 307760
rect 228416 307748 228422 307760
rect 246574 307748 246580 307760
rect 228416 307720 246580 307748
rect 228416 307708 228422 307720
rect 246574 307708 246580 307720
rect 246632 307708 246638 307760
rect 282914 307708 282920 307760
rect 282972 307748 282978 307760
rect 283742 307748 283748 307760
rect 282972 307720 283748 307748
rect 282972 307708 282978 307720
rect 283742 307708 283748 307720
rect 283800 307708 283806 307760
rect 285674 307708 285680 307760
rect 285732 307748 285738 307760
rect 286502 307748 286508 307760
rect 285732 307720 286508 307748
rect 285732 307708 285738 307720
rect 286502 307708 286508 307720
rect 286560 307708 286566 307760
rect 354950 307708 354956 307760
rect 355008 307748 355014 307760
rect 355134 307748 355140 307760
rect 355008 307720 355140 307748
rect 355008 307708 355014 307720
rect 355134 307708 355140 307720
rect 355192 307708 355198 307760
rect 171410 307640 171416 307692
rect 171468 307680 171474 307692
rect 246942 307680 246948 307692
rect 171468 307652 246948 307680
rect 171468 307640 171474 307652
rect 246942 307640 246948 307652
rect 247000 307640 247006 307692
rect 331582 307640 331588 307692
rect 331640 307680 331646 307692
rect 332410 307680 332416 307692
rect 331640 307652 332416 307680
rect 331640 307640 331646 307652
rect 332410 307640 332416 307652
rect 332468 307640 332474 307692
rect 171778 307572 171784 307624
rect 171836 307612 171842 307624
rect 244274 307612 244280 307624
rect 171836 307584 244280 307612
rect 171836 307572 171842 307584
rect 244274 307572 244280 307584
rect 244332 307572 244338 307624
rect 354766 307572 354772 307624
rect 354824 307612 354830 307624
rect 355502 307612 355508 307624
rect 354824 307584 355508 307612
rect 354824 307572 354830 307584
rect 355502 307572 355508 307584
rect 355560 307572 355566 307624
rect 229738 307504 229744 307556
rect 229796 307544 229802 307556
rect 250254 307544 250260 307556
rect 229796 307516 250260 307544
rect 229796 307504 229802 307516
rect 250254 307504 250260 307516
rect 250312 307504 250318 307556
rect 180058 307436 180064 307488
rect 180116 307476 180122 307488
rect 244826 307476 244832 307488
rect 180116 307448 244832 307476
rect 180116 307436 180122 307448
rect 244826 307436 244832 307448
rect 244884 307436 244890 307488
rect 220078 307368 220084 307420
rect 220136 307408 220142 307420
rect 242526 307408 242532 307420
rect 220136 307380 242532 307408
rect 220136 307368 220142 307380
rect 242526 307368 242532 307380
rect 242584 307368 242590 307420
rect 229830 307300 229836 307352
rect 229888 307340 229894 307352
rect 252278 307340 252284 307352
rect 229888 307312 252284 307340
rect 229888 307300 229894 307312
rect 252278 307300 252284 307312
rect 252336 307300 252342 307352
rect 332962 307300 332968 307352
rect 333020 307340 333026 307352
rect 333238 307340 333244 307352
rect 333020 307312 333244 307340
rect 333020 307300 333026 307312
rect 333238 307300 333244 307312
rect 333296 307300 333302 307352
rect 224218 307232 224224 307284
rect 224276 307272 224282 307284
rect 243722 307272 243728 307284
rect 224276 307244 243728 307272
rect 224276 307232 224282 307244
rect 243722 307232 243728 307244
rect 243780 307232 243786 307284
rect 339586 307232 339592 307284
rect 339644 307272 339650 307284
rect 340598 307272 340604 307284
rect 339644 307244 340604 307272
rect 339644 307232 339650 307244
rect 340598 307232 340604 307244
rect 340656 307232 340662 307284
rect 170398 307164 170404 307216
rect 170456 307204 170462 307216
rect 249978 307204 249984 307216
rect 170456 307176 249984 307204
rect 170456 307164 170462 307176
rect 249978 307164 249984 307176
rect 250036 307164 250042 307216
rect 314102 307164 314108 307216
rect 314160 307204 314166 307216
rect 378778 307204 378784 307216
rect 314160 307176 378784 307204
rect 314160 307164 314166 307176
rect 378778 307164 378784 307176
rect 378836 307164 378842 307216
rect 170582 307096 170588 307148
rect 170640 307136 170646 307148
rect 238386 307136 238392 307148
rect 170640 307108 238392 307136
rect 170640 307096 170646 307108
rect 238386 307096 238392 307108
rect 238444 307096 238450 307148
rect 243078 307096 243084 307148
rect 243136 307136 243142 307148
rect 243906 307136 243912 307148
rect 243136 307108 243912 307136
rect 243136 307096 243142 307108
rect 243906 307096 243912 307108
rect 243964 307096 243970 307148
rect 284938 307136 284944 307148
rect 273226 307108 284944 307136
rect 200114 307028 200120 307080
rect 200172 307068 200178 307080
rect 273226 307068 273254 307108
rect 284938 307096 284944 307108
rect 284996 307096 285002 307148
rect 317782 307096 317788 307148
rect 317840 307136 317846 307148
rect 402974 307136 402980 307148
rect 317840 307108 402980 307136
rect 317840 307096 317846 307108
rect 402974 307096 402980 307108
rect 403032 307096 403038 307148
rect 200172 307040 273254 307068
rect 200172 307028 200178 307040
rect 283098 307028 283104 307080
rect 283156 307068 283162 307080
rect 283926 307068 283932 307080
rect 283156 307040 283932 307068
rect 283156 307028 283162 307040
rect 283926 307028 283932 307040
rect 283984 307028 283990 307080
rect 340414 307028 340420 307080
rect 340472 307068 340478 307080
rect 543734 307068 543740 307080
rect 340472 307040 543740 307068
rect 340472 307028 340478 307040
rect 543734 307028 543740 307040
rect 543792 307028 543798 307080
rect 173158 306960 173164 307012
rect 173216 307000 173222 307012
rect 239674 307000 239680 307012
rect 173216 306972 239680 307000
rect 173216 306960 173222 306972
rect 239674 306960 239680 306972
rect 239732 306960 239738 307012
rect 253014 307000 253020 307012
rect 252848 306972 253020 307000
rect 252848 306808 252876 306972
rect 253014 306960 253020 306972
rect 253072 306960 253078 307012
rect 281718 306960 281724 307012
rect 281776 307000 281782 307012
rect 281994 307000 282000 307012
rect 281776 306972 282000 307000
rect 281776 306960 281782 306972
rect 281994 306960 282000 306972
rect 282052 306960 282058 307012
rect 297174 306960 297180 307012
rect 297232 306960 297238 307012
rect 321830 306960 321836 307012
rect 321888 307000 321894 307012
rect 322106 307000 322112 307012
rect 321888 306972 322112 307000
rect 321888 306960 321894 306972
rect 322106 306960 322112 306972
rect 322164 306960 322170 307012
rect 252830 306756 252836 306808
rect 252888 306756 252894 306808
rect 297082 306756 297088 306808
rect 297140 306796 297146 306808
rect 297192 306796 297220 306960
rect 330110 306824 330116 306876
rect 330168 306824 330174 306876
rect 356054 306824 356060 306876
rect 356112 306864 356118 306876
rect 357066 306864 357072 306876
rect 356112 306836 357072 306864
rect 356112 306824 356118 306836
rect 357066 306824 357072 306836
rect 357124 306824 357130 306876
rect 357526 306824 357532 306876
rect 357584 306864 357590 306876
rect 358354 306864 358360 306876
rect 357584 306836 358360 306864
rect 357584 306824 357590 306836
rect 358354 306824 358360 306836
rect 358412 306824 358418 306876
rect 297140 306768 297220 306796
rect 297140 306756 297146 306768
rect 267918 306688 267924 306740
rect 267976 306688 267982 306740
rect 295610 306688 295616 306740
rect 295668 306688 295674 306740
rect 300854 306688 300860 306740
rect 300912 306728 300918 306740
rect 301130 306728 301136 306740
rect 300912 306700 301136 306728
rect 300912 306688 300918 306700
rect 301130 306688 301136 306700
rect 301188 306688 301194 306740
rect 252738 306484 252744 306536
rect 252796 306524 252802 306536
rect 253106 306524 253112 306536
rect 252796 306496 253112 306524
rect 252796 306484 252802 306496
rect 253106 306484 253112 306496
rect 253164 306484 253170 306536
rect 256602 306484 256608 306536
rect 256660 306524 256666 306536
rect 257246 306524 257252 306536
rect 256660 306496 257252 306524
rect 256660 306484 256666 306496
rect 257246 306484 257252 306496
rect 257304 306484 257310 306536
rect 267936 306468 267964 306688
rect 295628 306468 295656 306688
rect 330128 306672 330156 306824
rect 342714 306688 342720 306740
rect 342772 306688 342778 306740
rect 360654 306688 360660 306740
rect 360712 306688 360718 306740
rect 328638 306620 328644 306672
rect 328696 306660 328702 306672
rect 328914 306660 328920 306672
rect 328696 306632 328920 306660
rect 328696 306620 328702 306632
rect 328914 306620 328920 306632
rect 328972 306620 328978 306672
rect 330110 306620 330116 306672
rect 330168 306620 330174 306672
rect 309318 306552 309324 306604
rect 309376 306552 309382 306604
rect 316218 306552 316224 306604
rect 316276 306592 316282 306604
rect 316862 306592 316868 306604
rect 316276 306564 316868 306592
rect 316276 306552 316282 306564
rect 316862 306552 316868 306564
rect 316920 306552 316926 306604
rect 317690 306552 317696 306604
rect 317748 306592 317754 306604
rect 318242 306592 318248 306604
rect 317748 306564 318248 306592
rect 317748 306552 317754 306564
rect 318242 306552 318248 306564
rect 318300 306552 318306 306604
rect 323302 306592 323308 306604
rect 322952 306564 323308 306592
rect 252646 306416 252652 306468
rect 252704 306456 252710 306468
rect 253474 306456 253480 306468
rect 252704 306428 253480 306456
rect 252704 306416 252710 306428
rect 253474 306416 253480 306428
rect 253532 306416 253538 306468
rect 256786 306416 256792 306468
rect 256844 306456 256850 306468
rect 257430 306456 257436 306468
rect 256844 306428 257436 306456
rect 256844 306416 256850 306428
rect 257430 306416 257436 306428
rect 257488 306416 257494 306468
rect 267918 306416 267924 306468
rect 267976 306416 267982 306468
rect 269206 306416 269212 306468
rect 269264 306456 269270 306468
rect 269666 306456 269672 306468
rect 269264 306428 269672 306456
rect 269264 306416 269270 306428
rect 269666 306416 269672 306428
rect 269724 306416 269730 306468
rect 270678 306416 270684 306468
rect 270736 306456 270742 306468
rect 270954 306456 270960 306468
rect 270736 306428 270960 306456
rect 270736 306416 270742 306428
rect 270954 306416 270960 306428
rect 271012 306416 271018 306468
rect 277394 306416 277400 306468
rect 277452 306456 277458 306468
rect 277854 306456 277860 306468
rect 277452 306428 277860 306456
rect 277452 306416 277458 306428
rect 277854 306416 277860 306428
rect 277912 306416 277918 306468
rect 278774 306416 278780 306468
rect 278832 306456 278838 306468
rect 279786 306456 279792 306468
rect 278832 306428 279792 306456
rect 278832 306416 278838 306428
rect 279786 306416 279792 306428
rect 279844 306416 279850 306468
rect 280338 306416 280344 306468
rect 280396 306456 280402 306468
rect 280798 306456 280804 306468
rect 280396 306428 280804 306456
rect 280396 306416 280402 306428
rect 280798 306416 280804 306428
rect 280856 306416 280862 306468
rect 295610 306416 295616 306468
rect 295668 306416 295674 306468
rect 305086 306416 305092 306468
rect 305144 306456 305150 306468
rect 305730 306456 305736 306468
rect 305144 306428 305736 306456
rect 305144 306416 305150 306428
rect 305730 306416 305736 306428
rect 305788 306416 305794 306468
rect 307294 306456 307300 306468
rect 306576 306428 307300 306456
rect 248506 306348 248512 306400
rect 248564 306388 248570 306400
rect 249242 306388 249248 306400
rect 248564 306360 249248 306388
rect 248564 306348 248570 306360
rect 249242 306348 249248 306360
rect 249300 306348 249306 306400
rect 264974 306348 264980 306400
rect 265032 306388 265038 306400
rect 265894 306388 265900 306400
rect 265032 306360 265900 306388
rect 265032 306348 265038 306360
rect 265894 306348 265900 306360
rect 265952 306348 265958 306400
rect 266630 306348 266636 306400
rect 266688 306388 266694 306400
rect 266998 306388 267004 306400
rect 266688 306360 267004 306388
rect 266688 306348 266694 306360
rect 266998 306348 267004 306360
rect 267056 306348 267062 306400
rect 272150 306348 272156 306400
rect 272208 306388 272214 306400
rect 272334 306388 272340 306400
rect 272208 306360 272340 306388
rect 272208 306348 272214 306360
rect 272334 306348 272340 306360
rect 272392 306348 272398 306400
rect 273714 306348 273720 306400
rect 273772 306388 273778 306400
rect 274450 306388 274456 306400
rect 273772 306360 274456 306388
rect 273772 306348 273778 306360
rect 274450 306348 274456 306360
rect 274508 306348 274514 306400
rect 279050 306348 279056 306400
rect 279108 306388 279114 306400
rect 279418 306388 279424 306400
rect 279108 306360 279424 306388
rect 279108 306348 279114 306360
rect 279418 306348 279424 306360
rect 279476 306348 279482 306400
rect 294138 306348 294144 306400
rect 294196 306388 294202 306400
rect 294874 306388 294880 306400
rect 294196 306360 294880 306388
rect 294196 306348 294202 306360
rect 294874 306348 294880 306360
rect 294932 306348 294938 306400
rect 295426 306348 295432 306400
rect 295484 306388 295490 306400
rect 296162 306388 296168 306400
rect 295484 306360 296168 306388
rect 295484 306348 295490 306360
rect 296162 306348 296168 306360
rect 296220 306348 296226 306400
rect 299566 306348 299572 306400
rect 299624 306388 299630 306400
rect 300578 306388 300584 306400
rect 299624 306360 300584 306388
rect 299624 306348 299630 306360
rect 300578 306348 300584 306360
rect 300636 306348 300642 306400
rect 301038 306348 301044 306400
rect 301096 306388 301102 306400
rect 302050 306388 302056 306400
rect 301096 306360 302056 306388
rect 301096 306348 301102 306360
rect 302050 306348 302056 306360
rect 302108 306348 302114 306400
rect 3326 306280 3332 306332
rect 3384 306320 3390 306332
rect 94498 306320 94504 306332
rect 3384 306292 94504 306320
rect 3384 306280 3390 306292
rect 94498 306280 94504 306292
rect 94556 306280 94562 306332
rect 169846 306280 169852 306332
rect 169904 306320 169910 306332
rect 243262 306320 243268 306332
rect 169904 306292 243268 306320
rect 169904 306280 169910 306292
rect 243262 306280 243268 306292
rect 243320 306280 243326 306332
rect 247126 306280 247132 306332
rect 247184 306320 247190 306332
rect 247862 306320 247868 306332
rect 247184 306292 247868 306320
rect 247184 306280 247190 306292
rect 247862 306280 247868 306292
rect 247920 306280 247926 306332
rect 248598 306280 248604 306332
rect 248656 306320 248662 306332
rect 249426 306320 249432 306332
rect 248656 306292 249432 306320
rect 248656 306280 248662 306292
rect 249426 306280 249432 306292
rect 249484 306280 249490 306332
rect 251726 306280 251732 306332
rect 251784 306320 251790 306332
rect 252094 306320 252100 306332
rect 251784 306292 252100 306320
rect 251784 306280 251790 306292
rect 252094 306280 252100 306292
rect 252152 306280 252158 306332
rect 253106 306280 253112 306332
rect 253164 306320 253170 306332
rect 253658 306320 253664 306332
rect 253164 306292 253664 306320
rect 253164 306280 253170 306292
rect 253658 306280 253664 306292
rect 253716 306280 253722 306332
rect 253934 306280 253940 306332
rect 253992 306320 253998 306332
rect 255130 306320 255136 306332
rect 253992 306292 255136 306320
rect 253992 306280 253998 306292
rect 255130 306280 255136 306292
rect 255188 306280 255194 306332
rect 255314 306280 255320 306332
rect 255372 306320 255378 306332
rect 255590 306320 255596 306332
rect 255372 306292 255596 306320
rect 255372 306280 255378 306292
rect 255590 306280 255596 306292
rect 255648 306280 255654 306332
rect 258534 306280 258540 306332
rect 258592 306320 258598 306332
rect 259362 306320 259368 306332
rect 258592 306292 259368 306320
rect 258592 306280 258598 306292
rect 259362 306280 259368 306292
rect 259420 306280 259426 306332
rect 259638 306280 259644 306332
rect 259696 306320 259702 306332
rect 260650 306320 260656 306332
rect 259696 306292 260656 306320
rect 259696 306280 259702 306292
rect 260650 306280 260656 306292
rect 260708 306280 260714 306332
rect 262398 306280 262404 306332
rect 262456 306320 262462 306332
rect 263134 306320 263140 306332
rect 262456 306292 263140 306320
rect 262456 306280 262462 306292
rect 263134 306280 263140 306292
rect 263192 306280 263198 306332
rect 265342 306280 265348 306332
rect 265400 306320 265406 306332
rect 266262 306320 266268 306332
rect 265400 306292 266268 306320
rect 265400 306280 265406 306292
rect 266262 306280 266268 306292
rect 266320 306280 266326 306332
rect 266538 306280 266544 306332
rect 266596 306320 266602 306332
rect 267366 306320 267372 306332
rect 266596 306292 267372 306320
rect 266596 306280 266602 306292
rect 267366 306280 267372 306292
rect 267424 306280 267430 306332
rect 267734 306280 267740 306332
rect 267792 306320 267798 306332
rect 268010 306320 268016 306332
rect 267792 306292 268016 306320
rect 267792 306280 267798 306292
rect 268010 306280 268016 306292
rect 268068 306280 268074 306332
rect 272058 306280 272064 306332
rect 272116 306320 272122 306332
rect 272518 306320 272524 306332
rect 272116 306292 272524 306320
rect 272116 306280 272122 306292
rect 272518 306280 272524 306292
rect 272576 306280 272582 306332
rect 273622 306280 273628 306332
rect 273680 306320 273686 306332
rect 274082 306320 274088 306332
rect 273680 306292 274088 306320
rect 273680 306280 273686 306292
rect 274082 306280 274088 306292
rect 274140 306280 274146 306332
rect 276198 306280 276204 306332
rect 276256 306320 276262 306332
rect 276750 306320 276756 306332
rect 276256 306292 276756 306320
rect 276256 306280 276262 306292
rect 276750 306280 276756 306292
rect 276808 306280 276814 306332
rect 277578 306280 277584 306332
rect 277636 306320 277642 306332
rect 278222 306320 278228 306332
rect 277636 306292 278228 306320
rect 277636 306280 277642 306292
rect 278222 306280 278228 306292
rect 278280 306280 278286 306332
rect 278866 306280 278872 306332
rect 278924 306320 278930 306332
rect 279142 306320 279148 306332
rect 278924 306292 279148 306320
rect 278924 306280 278930 306292
rect 279142 306280 279148 306292
rect 279200 306280 279206 306332
rect 294322 306280 294328 306332
rect 294380 306320 294386 306332
rect 295058 306320 295064 306332
rect 294380 306292 295064 306320
rect 294380 306280 294386 306292
rect 295058 306280 295064 306292
rect 295116 306280 295122 306332
rect 295518 306280 295524 306332
rect 295576 306320 295582 306332
rect 295978 306320 295984 306332
rect 295576 306292 295984 306320
rect 295576 306280 295582 306292
rect 295978 306280 295984 306292
rect 296036 306280 296042 306332
rect 296806 306280 296812 306332
rect 296864 306320 296870 306332
rect 297542 306320 297548 306332
rect 296864 306292 297548 306320
rect 296864 306280 296870 306292
rect 297542 306280 297548 306292
rect 297600 306280 297606 306332
rect 298554 306280 298560 306332
rect 298612 306320 298618 306332
rect 299198 306320 299204 306332
rect 298612 306292 299204 306320
rect 298612 306280 298618 306292
rect 299198 306280 299204 306292
rect 299256 306280 299262 306332
rect 299474 306280 299480 306332
rect 299532 306320 299538 306332
rect 300394 306320 300400 306332
rect 299532 306292 300400 306320
rect 299532 306280 299538 306292
rect 300394 306280 300400 306292
rect 300452 306280 300458 306332
rect 301130 306280 301136 306332
rect 301188 306320 301194 306332
rect 301498 306320 301504 306332
rect 301188 306292 301504 306320
rect 301188 306280 301194 306292
rect 301498 306280 301504 306292
rect 301556 306280 301562 306332
rect 302234 306280 302240 306332
rect 302292 306320 302298 306332
rect 303246 306320 303252 306332
rect 302292 306292 303252 306320
rect 302292 306280 302298 306292
rect 303246 306280 303252 306292
rect 303304 306280 303310 306332
rect 303798 306280 303804 306332
rect 303856 306320 303862 306332
rect 304350 306320 304356 306332
rect 303856 306292 304356 306320
rect 303856 306280 303862 306292
rect 304350 306280 304356 306292
rect 304408 306280 304414 306332
rect 305454 306320 305460 306332
rect 305196 306292 305460 306320
rect 305196 306264 305224 306292
rect 305454 306280 305460 306292
rect 305512 306280 305518 306332
rect 306576 306264 306604 306428
rect 307294 306416 307300 306428
rect 307352 306416 307358 306468
rect 307938 306416 307944 306468
rect 307996 306456 308002 306468
rect 308398 306456 308404 306468
rect 307996 306428 308404 306456
rect 307996 306416 308002 306428
rect 308398 306416 308404 306428
rect 308456 306416 308462 306468
rect 308122 306280 308128 306332
rect 308180 306320 308186 306332
rect 308582 306320 308588 306332
rect 308180 306292 308588 306320
rect 308180 306280 308186 306292
rect 308582 306280 308588 306292
rect 308640 306280 308646 306332
rect 215202 306212 215208 306264
rect 215260 306252 215266 306264
rect 288526 306252 288532 306264
rect 215260 306224 288532 306252
rect 215260 306212 215266 306224
rect 288526 306212 288532 306224
rect 288584 306212 288590 306264
rect 294230 306212 294236 306264
rect 294288 306252 294294 306264
rect 295242 306252 295248 306264
rect 294288 306224 295248 306252
rect 294288 306212 294294 306224
rect 295242 306212 295248 306224
rect 295300 306212 295306 306264
rect 303982 306212 303988 306264
rect 304040 306252 304046 306264
rect 304626 306252 304632 306264
rect 304040 306224 304632 306252
rect 304040 306212 304046 306224
rect 304626 306212 304632 306224
rect 304684 306212 304690 306264
rect 305178 306212 305184 306264
rect 305236 306212 305242 306264
rect 306558 306212 306564 306264
rect 306616 306212 306622 306264
rect 308214 306212 308220 306264
rect 308272 306252 308278 306264
rect 308766 306252 308772 306264
rect 308272 306224 308772 306252
rect 308272 306212 308278 306224
rect 308766 306212 308772 306224
rect 308824 306212 308830 306264
rect 309336 306252 309364 306552
rect 310606 306416 310612 306468
rect 310664 306456 310670 306468
rect 310882 306456 310888 306468
rect 310664 306428 310888 306456
rect 310664 306416 310670 306428
rect 310882 306416 310888 306428
rect 310940 306416 310946 306468
rect 311894 306416 311900 306468
rect 311952 306456 311958 306468
rect 312446 306456 312452 306468
rect 311952 306428 312452 306456
rect 311952 306416 311958 306428
rect 312446 306416 312452 306428
rect 312504 306416 312510 306468
rect 319070 306416 319076 306468
rect 319128 306456 319134 306468
rect 319346 306456 319352 306468
rect 319128 306428 319352 306456
rect 319128 306416 319134 306428
rect 319346 306416 319352 306428
rect 319404 306416 319410 306468
rect 313274 306348 313280 306400
rect 313332 306388 313338 306400
rect 313918 306388 313924 306400
rect 313332 306360 313924 306388
rect 313332 306348 313338 306360
rect 313918 306348 313924 306360
rect 313976 306348 313982 306400
rect 316034 306348 316040 306400
rect 316092 306388 316098 306400
rect 316218 306388 316224 306400
rect 316092 306360 316224 306388
rect 316092 306348 316098 306360
rect 316218 306348 316224 306360
rect 316276 306348 316282 306400
rect 317690 306348 317696 306400
rect 317748 306388 317754 306400
rect 318702 306388 318708 306400
rect 317748 306360 318708 306388
rect 317748 306348 317754 306360
rect 318702 306348 318708 306360
rect 318760 306348 318766 306400
rect 318794 306348 318800 306400
rect 318852 306388 318858 306400
rect 319438 306388 319444 306400
rect 318852 306360 319444 306388
rect 318852 306348 318858 306360
rect 319438 306348 319444 306360
rect 319496 306348 319502 306400
rect 320358 306348 320364 306400
rect 320416 306388 320422 306400
rect 320634 306388 320640 306400
rect 320416 306360 320640 306388
rect 320416 306348 320422 306360
rect 320634 306348 320640 306360
rect 320692 306348 320698 306400
rect 310974 306280 310980 306332
rect 311032 306320 311038 306332
rect 311618 306320 311624 306332
rect 311032 306292 311624 306320
rect 311032 306280 311038 306292
rect 311618 306280 311624 306292
rect 311676 306280 311682 306332
rect 313550 306280 313556 306332
rect 313608 306320 313614 306332
rect 313826 306320 313832 306332
rect 313608 306292 313832 306320
rect 313608 306280 313614 306292
rect 313826 306280 313832 306292
rect 313884 306280 313890 306332
rect 314746 306280 314752 306332
rect 314804 306320 314810 306332
rect 315482 306320 315488 306332
rect 314804 306292 315488 306320
rect 314804 306280 314810 306292
rect 315482 306280 315488 306292
rect 315540 306280 315546 306332
rect 317598 306280 317604 306332
rect 317656 306320 317662 306332
rect 318334 306320 318340 306332
rect 317656 306292 318340 306320
rect 317656 306280 317662 306292
rect 318334 306280 318340 306292
rect 318392 306280 318398 306332
rect 319162 306280 319168 306332
rect 319220 306320 319226 306332
rect 319806 306320 319812 306332
rect 319220 306292 319812 306320
rect 319220 306280 319226 306292
rect 319806 306280 319812 306292
rect 319864 306280 319870 306332
rect 320174 306280 320180 306332
rect 320232 306320 320238 306332
rect 321186 306320 321192 306332
rect 320232 306292 321192 306320
rect 320232 306280 320238 306292
rect 321186 306280 321192 306292
rect 321244 306280 321250 306332
rect 321830 306280 321836 306332
rect 321888 306320 321894 306332
rect 322658 306320 322664 306332
rect 321888 306292 322664 306320
rect 321888 306280 321894 306292
rect 322658 306280 322664 306292
rect 322716 306280 322722 306332
rect 322952 306264 322980 306564
rect 323302 306552 323308 306564
rect 323360 306552 323366 306604
rect 325786 306552 325792 306604
rect 325844 306592 325850 306604
rect 326430 306592 326436 306604
rect 325844 306564 326436 306592
rect 325844 306552 325850 306564
rect 326430 306552 326436 306564
rect 326488 306552 326494 306604
rect 328454 306552 328460 306604
rect 328512 306592 328518 306604
rect 329098 306592 329104 306604
rect 328512 306564 329104 306592
rect 328512 306552 328518 306564
rect 329098 306552 329104 306564
rect 329156 306552 329162 306604
rect 324406 306484 324412 306536
rect 324464 306524 324470 306536
rect 325234 306524 325240 306536
rect 324464 306496 325240 306524
rect 324464 306484 324470 306496
rect 325234 306484 325240 306496
rect 325292 306484 325298 306536
rect 340874 306484 340880 306536
rect 340932 306524 340938 306536
rect 341702 306524 341708 306536
rect 340932 306496 341708 306524
rect 340932 306484 340938 306496
rect 341702 306484 341708 306496
rect 341760 306484 341766 306536
rect 342732 306468 342760 306688
rect 360672 306468 360700 306688
rect 324774 306456 324780 306468
rect 324424 306428 324780 306456
rect 323210 306280 323216 306332
rect 323268 306320 323274 306332
rect 323486 306320 323492 306332
rect 323268 306292 323492 306320
rect 323268 306280 323274 306292
rect 323486 306280 323492 306292
rect 323544 306280 323550 306332
rect 324424 306264 324452 306428
rect 324774 306416 324780 306428
rect 324832 306416 324838 306468
rect 342714 306416 342720 306468
rect 342772 306416 342778 306468
rect 360654 306416 360660 306468
rect 360712 306416 360718 306468
rect 325786 306348 325792 306400
rect 325844 306388 325850 306400
rect 326890 306388 326896 306400
rect 325844 306360 326896 306388
rect 325844 306348 325850 306360
rect 326890 306348 326896 306360
rect 326948 306348 326954 306400
rect 340874 306348 340880 306400
rect 340932 306388 340938 306400
rect 341426 306388 341432 306400
rect 340932 306360 341432 306388
rect 340932 306348 340938 306360
rect 341426 306348 341432 306360
rect 341484 306348 341490 306400
rect 347774 306348 347780 306400
rect 347832 306388 347838 306400
rect 349062 306388 349068 306400
rect 347832 306360 349068 306388
rect 347832 306348 347838 306360
rect 349062 306348 349068 306360
rect 349120 306348 349126 306400
rect 325878 306280 325884 306332
rect 325936 306320 325942 306332
rect 326522 306320 326528 306332
rect 325936 306292 326528 306320
rect 325936 306280 325942 306292
rect 326522 306280 326528 306292
rect 326580 306280 326586 306332
rect 327442 306280 327448 306332
rect 327500 306320 327506 306332
rect 327626 306320 327632 306332
rect 327500 306292 327632 306320
rect 327500 306280 327506 306292
rect 327626 306280 327632 306292
rect 327684 306280 327690 306332
rect 328546 306280 328552 306332
rect 328604 306320 328610 306332
rect 329742 306320 329748 306332
rect 328604 306292 329748 306320
rect 328604 306280 328610 306292
rect 329742 306280 329748 306292
rect 329800 306280 329806 306332
rect 329834 306280 329840 306332
rect 329892 306320 329898 306332
rect 330386 306320 330392 306332
rect 329892 306292 330392 306320
rect 329892 306280 329898 306292
rect 330386 306280 330392 306292
rect 330444 306280 330450 306332
rect 341150 306280 341156 306332
rect 341208 306320 341214 306332
rect 342162 306320 342168 306332
rect 341208 306292 342168 306320
rect 341208 306280 341214 306292
rect 342162 306280 342168 306292
rect 342220 306280 342226 306332
rect 342622 306280 342628 306332
rect 342680 306320 342686 306332
rect 343266 306320 343272 306332
rect 342680 306292 343272 306320
rect 342680 306280 342686 306292
rect 343266 306280 343272 306292
rect 343324 306280 343330 306332
rect 343818 306280 343824 306332
rect 343876 306320 343882 306332
rect 344646 306320 344652 306332
rect 343876 306292 344652 306320
rect 343876 306280 343882 306292
rect 344646 306280 344652 306292
rect 344704 306280 344710 306332
rect 345014 306280 345020 306332
rect 345072 306320 345078 306332
rect 345750 306320 345756 306332
rect 345072 306292 345756 306320
rect 345072 306280 345078 306292
rect 345750 306280 345756 306292
rect 345808 306280 345814 306332
rect 347866 306280 347872 306332
rect 347924 306320 347930 306332
rect 348234 306320 348240 306332
rect 347924 306292 348240 306320
rect 347924 306280 347930 306292
rect 348234 306280 348240 306292
rect 348292 306280 348298 306332
rect 354858 306280 354864 306332
rect 354916 306320 354922 306332
rect 370406 306320 370412 306332
rect 354916 306292 370412 306320
rect 354916 306280 354922 306292
rect 370406 306280 370412 306292
rect 370464 306280 370470 306332
rect 309502 306252 309508 306264
rect 309336 306224 309508 306252
rect 309502 306212 309508 306224
rect 309560 306212 309566 306264
rect 310698 306212 310704 306264
rect 310756 306252 310762 306264
rect 311250 306252 311256 306264
rect 310756 306224 311256 306252
rect 310756 306212 310762 306224
rect 311250 306212 311256 306224
rect 311308 306212 311314 306264
rect 317414 306212 317420 306264
rect 317472 306252 317478 306264
rect 318518 306252 318524 306264
rect 317472 306224 318524 306252
rect 317472 306212 317478 306224
rect 318518 306212 318524 306224
rect 318576 306212 318582 306264
rect 321554 306212 321560 306264
rect 321612 306252 321618 306264
rect 322014 306252 322020 306264
rect 321612 306224 322020 306252
rect 321612 306212 321618 306224
rect 322014 306212 322020 306224
rect 322072 306212 322078 306264
rect 322934 306212 322940 306264
rect 322992 306212 322998 306264
rect 323394 306212 323400 306264
rect 323452 306252 323458 306264
rect 324038 306252 324044 306264
rect 323452 306224 324044 306252
rect 323452 306212 323458 306224
rect 324038 306212 324044 306224
rect 324096 306212 324102 306264
rect 324406 306212 324412 306264
rect 324464 306212 324470 306264
rect 324498 306212 324504 306264
rect 324556 306252 324562 306264
rect 325326 306252 325332 306264
rect 324556 306224 325332 306252
rect 324556 306212 324562 306224
rect 325326 306212 325332 306224
rect 325384 306212 325390 306264
rect 327074 306212 327080 306264
rect 327132 306252 327138 306264
rect 328270 306252 328276 306264
rect 327132 306224 328276 306252
rect 327132 306212 327138 306224
rect 328270 306212 328276 306224
rect 328328 306212 328334 306264
rect 328730 306212 328736 306264
rect 328788 306252 328794 306264
rect 329374 306252 329380 306264
rect 328788 306224 329380 306252
rect 328788 306212 328794 306224
rect 329374 306212 329380 306224
rect 329432 306212 329438 306264
rect 330018 306212 330024 306264
rect 330076 306252 330082 306264
rect 331122 306252 331128 306264
rect 330076 306224 331128 306252
rect 330076 306212 330082 306224
rect 331122 306212 331128 306224
rect 331180 306212 331186 306264
rect 340966 306212 340972 306264
rect 341024 306252 341030 306264
rect 341794 306252 341800 306264
rect 341024 306224 341800 306252
rect 341024 306212 341030 306224
rect 341794 306212 341800 306224
rect 341852 306212 341858 306264
rect 342346 306212 342352 306264
rect 342404 306252 342410 306264
rect 342898 306252 342904 306264
rect 342404 306224 342904 306252
rect 342404 306212 342410 306224
rect 342898 306212 342904 306224
rect 342956 306212 342962 306264
rect 343726 306212 343732 306264
rect 343784 306252 343790 306264
rect 344278 306252 344284 306264
rect 343784 306224 344284 306252
rect 343784 306212 343790 306224
rect 344278 306212 344284 306224
rect 344336 306212 344342 306264
rect 345198 306212 345204 306264
rect 345256 306252 345262 306264
rect 345382 306252 345388 306264
rect 345256 306224 345388 306252
rect 345256 306212 345262 306224
rect 345382 306212 345388 306224
rect 345440 306212 345446 306264
rect 352374 306212 352380 306264
rect 352432 306252 352438 306264
rect 360194 306252 360200 306264
rect 352432 306224 360200 306252
rect 352432 306212 352438 306224
rect 360194 306212 360200 306224
rect 360252 306212 360258 306264
rect 360286 306212 360292 306264
rect 360344 306252 360350 306264
rect 360838 306252 360844 306264
rect 360344 306224 360844 306252
rect 360344 306212 360350 306224
rect 360838 306212 360844 306224
rect 360896 306212 360902 306264
rect 218974 306144 218980 306196
rect 219032 306184 219038 306196
rect 293494 306184 293500 306196
rect 219032 306156 293500 306184
rect 219032 306144 219038 306156
rect 293494 306144 293500 306156
rect 293552 306144 293558 306196
rect 295610 306144 295616 306196
rect 295668 306184 295674 306196
rect 296346 306184 296352 306196
rect 295668 306156 296352 306184
rect 295668 306144 295674 306156
rect 296346 306144 296352 306156
rect 296404 306144 296410 306196
rect 309134 306144 309140 306196
rect 309192 306184 309198 306196
rect 310146 306184 310152 306196
rect 309192 306156 310152 306184
rect 309192 306144 309198 306156
rect 310146 306144 310152 306156
rect 310204 306144 310210 306196
rect 310790 306144 310796 306196
rect 310848 306184 310854 306196
rect 311802 306184 311808 306196
rect 310848 306156 311808 306184
rect 310848 306144 310854 306156
rect 311802 306144 311808 306156
rect 311860 306144 311866 306196
rect 311986 306144 311992 306196
rect 312044 306184 312050 306196
rect 313182 306184 313188 306196
rect 312044 306156 313188 306184
rect 312044 306144 312050 306156
rect 313182 306144 313188 306156
rect 313240 306144 313246 306196
rect 313550 306144 313556 306196
rect 313608 306184 313614 306196
rect 314286 306184 314292 306196
rect 313608 306156 314292 306184
rect 313608 306144 313614 306156
rect 314286 306144 314292 306156
rect 314344 306144 314350 306196
rect 314930 306144 314936 306196
rect 314988 306184 314994 306196
rect 315850 306184 315856 306196
rect 314988 306156 315856 306184
rect 314988 306144 314994 306156
rect 315850 306144 315856 306156
rect 315908 306144 315914 306196
rect 316402 306144 316408 306196
rect 316460 306184 316466 306196
rect 317138 306184 317144 306196
rect 316460 306156 317144 306184
rect 316460 306144 316466 306156
rect 317138 306144 317144 306156
rect 317196 306144 317202 306196
rect 317782 306144 317788 306196
rect 317840 306184 317846 306196
rect 318150 306184 318156 306196
rect 317840 306156 318156 306184
rect 317840 306144 317846 306156
rect 318150 306144 318156 306156
rect 318208 306144 318214 306196
rect 318978 306144 318984 306196
rect 319036 306184 319042 306196
rect 319622 306184 319628 306196
rect 319036 306156 319628 306184
rect 319036 306144 319042 306156
rect 319622 306144 319628 306156
rect 319680 306144 319686 306196
rect 321738 306144 321744 306196
rect 321796 306184 321802 306196
rect 322474 306184 322480 306196
rect 321796 306156 322480 306184
rect 321796 306144 321802 306156
rect 322474 306144 322480 306156
rect 322532 306144 322538 306196
rect 323026 306144 323032 306196
rect 323084 306184 323090 306196
rect 323854 306184 323860 306196
rect 323084 306156 323860 306184
rect 323084 306144 323090 306156
rect 323854 306144 323860 306156
rect 323912 306144 323918 306196
rect 324590 306144 324596 306196
rect 324648 306184 324654 306196
rect 325602 306184 325608 306196
rect 324648 306156 325608 306184
rect 324648 306144 324654 306156
rect 325602 306144 325608 306156
rect 325660 306144 325666 306196
rect 328822 306144 328828 306196
rect 328880 306184 328886 306196
rect 329558 306184 329564 306196
rect 328880 306156 329564 306184
rect 328880 306144 328886 306156
rect 329558 306144 329564 306156
rect 329616 306144 329622 306196
rect 341242 306144 341248 306196
rect 341300 306184 341306 306196
rect 341610 306184 341616 306196
rect 341300 306156 341616 306184
rect 341300 306144 341306 306156
rect 341610 306144 341616 306156
rect 341668 306144 341674 306196
rect 352190 306144 352196 306196
rect 352248 306184 352254 306196
rect 368658 306184 368664 306196
rect 352248 306156 368664 306184
rect 352248 306144 352254 306156
rect 368658 306144 368664 306156
rect 368716 306144 368722 306196
rect 216398 306076 216404 306128
rect 216456 306116 216462 306128
rect 291470 306116 291476 306128
rect 216456 306088 291476 306116
rect 216456 306076 216462 306088
rect 291470 306076 291476 306088
rect 291528 306076 291534 306128
rect 304994 306076 305000 306128
rect 305052 306116 305058 306128
rect 305362 306116 305368 306128
rect 305052 306088 305368 306116
rect 305052 306076 305058 306088
rect 305362 306076 305368 306088
rect 305420 306076 305426 306128
rect 305454 306076 305460 306128
rect 305512 306116 305518 306128
rect 306282 306116 306288 306128
rect 305512 306088 306288 306116
rect 305512 306076 305518 306088
rect 306282 306076 306288 306088
rect 306340 306076 306346 306128
rect 307938 306076 307944 306128
rect 307996 306116 308002 306128
rect 308950 306116 308956 306128
rect 307996 306088 308956 306116
rect 307996 306076 308002 306088
rect 308950 306076 308956 306088
rect 309008 306076 309014 306128
rect 313366 306076 313372 306128
rect 313424 306116 313430 306128
rect 314470 306116 314476 306128
rect 313424 306088 314476 306116
rect 313424 306076 313430 306088
rect 314470 306076 314476 306088
rect 314528 306076 314534 306128
rect 314654 306076 314660 306128
rect 314712 306116 314718 306128
rect 315114 306116 315120 306128
rect 314712 306088 315120 306116
rect 314712 306076 314718 306088
rect 315114 306076 315120 306088
rect 315172 306076 315178 306128
rect 318886 306076 318892 306128
rect 318944 306116 318950 306128
rect 319990 306116 319996 306128
rect 318944 306088 319996 306116
rect 318944 306076 318950 306088
rect 319990 306076 319996 306088
rect 320048 306076 320054 306128
rect 320266 306076 320272 306128
rect 320324 306116 320330 306128
rect 320634 306116 320640 306128
rect 320324 306088 320640 306116
rect 320324 306076 320330 306088
rect 320634 306076 320640 306088
rect 320692 306076 320698 306128
rect 321554 306076 321560 306128
rect 321612 306116 321618 306128
rect 322290 306116 322296 306128
rect 321612 306088 322296 306116
rect 321612 306076 321618 306088
rect 322290 306076 322296 306088
rect 322348 306076 322354 306128
rect 328638 306076 328644 306128
rect 328696 306116 328702 306128
rect 329190 306116 329196 306128
rect 328696 306088 329196 306116
rect 328696 306076 328702 306088
rect 329190 306076 329196 306088
rect 329248 306076 329254 306128
rect 341058 306076 341064 306128
rect 341116 306116 341122 306128
rect 341426 306116 341432 306128
rect 341116 306088 341432 306116
rect 341116 306076 341122 306088
rect 341426 306076 341432 306088
rect 341484 306076 341490 306128
rect 345198 306076 345204 306128
rect 345256 306116 345262 306128
rect 346210 306116 346216 306128
rect 345256 306088 346216 306116
rect 345256 306076 345262 306088
rect 346210 306076 346216 306088
rect 346268 306076 346274 306128
rect 354766 306076 354772 306128
rect 354824 306116 354830 306128
rect 371418 306116 371424 306128
rect 354824 306088 371424 306116
rect 354824 306076 354830 306088
rect 371418 306076 371424 306088
rect 371476 306076 371482 306128
rect 216306 306008 216312 306060
rect 216364 306048 216370 306060
rect 292942 306048 292948 306060
rect 216364 306020 292948 306048
rect 216364 306008 216370 306020
rect 292942 306008 292948 306020
rect 293000 306008 293006 306060
rect 320450 306008 320456 306060
rect 320508 306048 320514 306060
rect 321002 306048 321008 306060
rect 320508 306020 321008 306048
rect 320508 306008 320514 306020
rect 321002 306008 321008 306020
rect 321060 306008 321066 306060
rect 343910 306008 343916 306060
rect 343968 306008 343974 306060
rect 354950 306008 354956 306060
rect 355008 306048 355014 306060
rect 371694 306048 371700 306060
rect 355008 306020 371700 306048
rect 355008 306008 355014 306020
rect 371694 306008 371700 306020
rect 371752 306008 371758 306060
rect 213638 305940 213644 305992
rect 213696 305980 213702 305992
rect 294046 305980 294052 305992
rect 213696 305952 294052 305980
rect 213696 305940 213702 305952
rect 294046 305940 294052 305952
rect 294104 305940 294110 305992
rect 304994 305940 305000 305992
rect 305052 305980 305058 305992
rect 306098 305980 306104 305992
rect 305052 305952 306104 305980
rect 305052 305940 305058 305952
rect 306098 305940 306104 305952
rect 306156 305940 306162 305992
rect 306834 305940 306840 305992
rect 306892 305980 306898 305992
rect 307662 305980 307668 305992
rect 306892 305952 307668 305980
rect 306892 305940 306898 305952
rect 307662 305940 307668 305952
rect 307720 305940 307726 305992
rect 320266 305940 320272 305992
rect 320324 305980 320330 305992
rect 321370 305980 321376 305992
rect 320324 305952 321376 305980
rect 320324 305940 320330 305952
rect 321370 305940 321376 305952
rect 321428 305940 321434 305992
rect 327350 305940 327356 305992
rect 327408 305980 327414 305992
rect 327810 305980 327816 305992
rect 327408 305952 327816 305980
rect 327408 305940 327414 305952
rect 327810 305940 327816 305952
rect 327868 305940 327874 305992
rect 341058 305940 341064 305992
rect 341116 305980 341122 305992
rect 341978 305980 341984 305992
rect 341116 305952 341984 305980
rect 341116 305940 341122 305952
rect 341978 305940 341984 305952
rect 342036 305940 342042 305992
rect 216582 305872 216588 305924
rect 216640 305912 216646 305924
rect 298462 305912 298468 305924
rect 216640 305884 298468 305912
rect 216640 305872 216646 305884
rect 298462 305872 298468 305884
rect 298520 305872 298526 305924
rect 327442 305872 327448 305924
rect 327500 305912 327506 305924
rect 327718 305912 327724 305924
rect 327500 305884 327724 305912
rect 327500 305872 327506 305884
rect 327718 305872 327724 305884
rect 327776 305872 327782 305924
rect 170398 305804 170404 305856
rect 170456 305844 170462 305856
rect 253934 305844 253940 305856
rect 170456 305816 253940 305844
rect 170456 305804 170462 305816
rect 253934 305804 253940 305816
rect 253992 305804 253998 305856
rect 254026 305804 254032 305856
rect 254084 305844 254090 305856
rect 254210 305844 254216 305856
rect 254084 305816 254216 305844
rect 254084 305804 254090 305816
rect 254210 305804 254216 305816
rect 254268 305804 254274 305856
rect 255682 305804 255688 305856
rect 255740 305844 255746 305856
rect 255866 305844 255872 305856
rect 255740 305816 255872 305844
rect 255740 305804 255746 305816
rect 255866 305804 255872 305816
rect 255924 305804 255930 305856
rect 257154 305804 257160 305856
rect 257212 305844 257218 305856
rect 257430 305844 257436 305856
rect 257212 305816 257436 305844
rect 257212 305804 257218 305816
rect 257430 305804 257436 305816
rect 257488 305804 257494 305856
rect 258074 305804 258080 305856
rect 258132 305844 258138 305856
rect 258350 305844 258356 305856
rect 258132 305816 258356 305844
rect 258132 305804 258138 305816
rect 258350 305804 258356 305816
rect 258408 305804 258414 305856
rect 258442 305804 258448 305856
rect 258500 305844 258506 305856
rect 259178 305844 259184 305856
rect 258500 305816 259184 305844
rect 258500 305804 258506 305816
rect 259178 305804 259184 305816
rect 259236 305804 259242 305856
rect 262582 305804 262588 305856
rect 262640 305844 262646 305856
rect 263318 305844 263324 305856
rect 262640 305816 263324 305844
rect 262640 305804 262646 305816
rect 263318 305804 263324 305816
rect 263376 305804 263382 305856
rect 263594 305804 263600 305856
rect 263652 305844 263658 305856
rect 263778 305844 263784 305856
rect 263652 305816 263784 305844
rect 263652 305804 263658 305816
rect 263778 305804 263784 305816
rect 263836 305804 263842 305856
rect 264054 305804 264060 305856
rect 264112 305844 264118 305856
rect 264882 305844 264888 305856
rect 264112 305816 264888 305844
rect 264112 305804 264118 305816
rect 264882 305804 264888 305816
rect 264940 305804 264946 305856
rect 265066 305804 265072 305856
rect 265124 305844 265130 305856
rect 265250 305844 265256 305856
rect 265124 305816 265256 305844
rect 265124 305804 265130 305816
rect 265250 305804 265256 305816
rect 265308 305804 265314 305856
rect 266722 305804 266728 305856
rect 266780 305844 266786 305856
rect 267550 305844 267556 305856
rect 266780 305816 267556 305844
rect 266780 305804 266786 305816
rect 267550 305804 267556 305816
rect 267608 305804 267614 305856
rect 269114 305804 269120 305856
rect 269172 305844 269178 305856
rect 269482 305844 269488 305856
rect 269172 305816 269488 305844
rect 269172 305804 269178 305816
rect 269482 305804 269488 305816
rect 269540 305804 269546 305856
rect 269574 305804 269580 305856
rect 269632 305844 269638 305856
rect 270034 305844 270040 305856
rect 269632 305816 270040 305844
rect 269632 305804 269638 305816
rect 270034 305804 270040 305816
rect 270092 305804 270098 305856
rect 270586 305804 270592 305856
rect 270644 305844 270650 305856
rect 271046 305844 271052 305856
rect 270644 305816 271052 305844
rect 270644 305804 270650 305816
rect 271046 305804 271052 305816
rect 271104 305804 271110 305856
rect 272242 305804 272248 305856
rect 272300 305844 272306 305856
rect 273070 305844 273076 305856
rect 272300 305816 273076 305844
rect 272300 305804 272306 305816
rect 273070 305804 273076 305816
rect 273128 305804 273134 305856
rect 273346 305804 273352 305856
rect 273404 305844 273410 305856
rect 274266 305844 274272 305856
rect 273404 305816 274272 305844
rect 273404 305804 273410 305816
rect 274266 305804 274272 305816
rect 274324 305804 274330 305856
rect 274634 305804 274640 305856
rect 274692 305844 274698 305856
rect 275738 305844 275744 305856
rect 274692 305816 275744 305844
rect 274692 305804 274698 305816
rect 275738 305804 275744 305816
rect 275796 305804 275802 305856
rect 276290 305804 276296 305856
rect 276348 305844 276354 305856
rect 276842 305844 276848 305856
rect 276348 305816 276848 305844
rect 276348 305804 276354 305816
rect 276842 305804 276848 305816
rect 276900 305804 276906 305856
rect 277486 305804 277492 305856
rect 277544 305844 277550 305856
rect 277854 305844 277860 305856
rect 277544 305816 277860 305844
rect 277544 305804 277550 305816
rect 277854 305804 277860 305816
rect 277912 305804 277918 305856
rect 279234 305804 279240 305856
rect 279292 305844 279298 305856
rect 279970 305844 279976 305856
rect 279292 305816 279976 305844
rect 279292 305804 279298 305816
rect 279970 305804 279976 305816
rect 280028 305804 280034 305856
rect 280430 305804 280436 305856
rect 280488 305844 280494 305856
rect 281074 305844 281080 305856
rect 280488 305816 281080 305844
rect 280488 305804 280494 305816
rect 281074 305804 281080 305816
rect 281132 305804 281138 305856
rect 281810 305804 281816 305856
rect 281868 305844 281874 305856
rect 282270 305844 282276 305856
rect 281868 305816 282276 305844
rect 281868 305804 281874 305816
rect 282270 305804 282276 305816
rect 282328 305804 282334 305856
rect 293034 305804 293040 305856
rect 293092 305844 293098 305856
rect 293678 305844 293684 305856
rect 293092 305816 293684 305844
rect 293092 305804 293098 305816
rect 293678 305804 293684 305816
rect 293736 305804 293742 305856
rect 306374 305804 306380 305856
rect 306432 305844 306438 305856
rect 306926 305844 306932 305856
rect 306432 305816 306932 305844
rect 306432 305804 306438 305816
rect 306926 305804 306932 305816
rect 306984 305804 306990 305856
rect 343928 305844 343956 306008
rect 354674 305940 354680 305992
rect 354732 305980 354738 305992
rect 371510 305980 371516 305992
rect 354732 305952 371516 305980
rect 354732 305940 354738 305952
rect 371510 305940 371516 305952
rect 371568 305940 371574 305992
rect 352282 305872 352288 305924
rect 352340 305912 352346 305924
rect 370314 305912 370320 305924
rect 352340 305884 370320 305912
rect 352340 305872 352346 305884
rect 370314 305872 370320 305884
rect 370372 305872 370378 305924
rect 344094 305844 344100 305856
rect 343928 305816 344100 305844
rect 344094 305804 344100 305816
rect 344152 305804 344158 305856
rect 350810 305804 350816 305856
rect 350868 305844 350874 305856
rect 360286 305844 360292 305856
rect 350868 305816 360292 305844
rect 350868 305804 350874 305816
rect 360286 305804 360292 305816
rect 360344 305804 360350 305856
rect 360562 305804 360568 305856
rect 360620 305844 360626 305856
rect 361206 305844 361212 305856
rect 360620 305816 361212 305844
rect 360620 305804 360626 305816
rect 361206 305804 361212 305816
rect 361264 305804 361270 305856
rect 210970 305736 210976 305788
rect 211028 305776 211034 305788
rect 211028 305748 292574 305776
rect 211028 305736 211034 305748
rect 195974 305668 195980 305720
rect 196032 305708 196038 305720
rect 284846 305708 284852 305720
rect 196032 305680 284852 305708
rect 196032 305668 196038 305680
rect 284846 305668 284852 305680
rect 284904 305668 284910 305720
rect 292546 305708 292574 305748
rect 292942 305736 292948 305788
rect 293000 305776 293006 305788
rect 293862 305776 293868 305788
rect 293000 305748 293868 305776
rect 293000 305736 293006 305748
rect 293862 305736 293868 305748
rect 293920 305736 293926 305788
rect 342254 305736 342260 305788
rect 342312 305776 342318 305788
rect 343082 305776 343088 305788
rect 342312 305748 343088 305776
rect 342312 305736 342318 305748
rect 343082 305736 343088 305748
rect 343140 305736 343146 305788
rect 353386 305736 353392 305788
rect 353444 305776 353450 305788
rect 371602 305776 371608 305788
rect 353444 305748 371608 305776
rect 353444 305736 353450 305748
rect 371602 305736 371608 305748
rect 371660 305736 371666 305788
rect 295886 305708 295892 305720
rect 292546 305680 295892 305708
rect 295886 305668 295892 305680
rect 295944 305668 295950 305720
rect 306374 305668 306380 305720
rect 306432 305708 306438 305720
rect 307202 305708 307208 305720
rect 306432 305680 307208 305708
rect 306432 305668 306438 305680
rect 307202 305668 307208 305680
rect 307260 305668 307266 305720
rect 347130 305668 347136 305720
rect 347188 305708 347194 305720
rect 364978 305708 364984 305720
rect 347188 305680 364984 305708
rect 347188 305668 347194 305680
rect 364978 305668 364984 305680
rect 365036 305668 365042 305720
rect 178034 305600 178040 305652
rect 178092 305640 178098 305652
rect 275830 305640 275836 305652
rect 178092 305612 275836 305640
rect 178092 305600 178098 305612
rect 275830 305600 275836 305612
rect 275888 305600 275894 305652
rect 276290 305600 276296 305652
rect 276348 305640 276354 305652
rect 277118 305640 277124 305652
rect 276348 305612 277124 305640
rect 276348 305600 276354 305612
rect 277118 305600 277124 305612
rect 277176 305600 277182 305652
rect 277486 305600 277492 305652
rect 277544 305640 277550 305652
rect 278406 305640 278412 305652
rect 277544 305612 278412 305640
rect 277544 305600 277550 305612
rect 278406 305600 278412 305612
rect 278464 305600 278470 305652
rect 278866 305600 278872 305652
rect 278924 305640 278930 305652
rect 279602 305640 279608 305652
rect 278924 305612 279608 305640
rect 278924 305600 278930 305612
rect 279602 305600 279608 305612
rect 279660 305600 279666 305652
rect 280246 305600 280252 305652
rect 280304 305640 280310 305652
rect 280890 305640 280896 305652
rect 280304 305612 280896 305640
rect 280304 305600 280310 305612
rect 280890 305600 280896 305612
rect 280948 305600 280954 305652
rect 281718 305600 281724 305652
rect 281776 305640 281782 305652
rect 282822 305640 282828 305652
rect 281776 305612 282828 305640
rect 281776 305600 281782 305612
rect 282822 305600 282828 305612
rect 282880 305600 282886 305652
rect 353294 305600 353300 305652
rect 353352 305640 353358 305652
rect 371786 305640 371792 305652
rect 353352 305612 371792 305640
rect 353352 305600 353358 305612
rect 371786 305600 371792 305612
rect 371844 305600 371850 305652
rect 219066 305532 219072 305584
rect 219124 305572 219130 305584
rect 291286 305572 291292 305584
rect 219124 305544 291292 305572
rect 219124 305532 219130 305544
rect 291286 305532 291292 305544
rect 291344 305532 291350 305584
rect 353570 305532 353576 305584
rect 353628 305572 353634 305584
rect 368934 305572 368940 305584
rect 353628 305544 368940 305572
rect 353628 305532 353634 305544
rect 368934 305532 368940 305544
rect 368992 305532 368998 305584
rect 218882 305464 218888 305516
rect 218940 305504 218946 305516
rect 289814 305504 289820 305516
rect 218940 305476 289820 305504
rect 218940 305464 218946 305476
rect 289814 305464 289820 305476
rect 289872 305464 289878 305516
rect 356146 305464 356152 305516
rect 356204 305504 356210 305516
rect 367738 305504 367744 305516
rect 356204 305476 367744 305504
rect 356204 305464 356210 305476
rect 367738 305464 367744 305476
rect 367796 305464 367802 305516
rect 171686 305396 171692 305448
rect 171744 305436 171750 305448
rect 234982 305436 234988 305448
rect 171744 305408 234988 305436
rect 171744 305396 171750 305408
rect 234982 305396 234988 305408
rect 235040 305396 235046 305448
rect 251358 305396 251364 305448
rect 251416 305436 251422 305448
rect 251634 305436 251640 305448
rect 251416 305408 251640 305436
rect 251416 305396 251422 305408
rect 251634 305396 251640 305408
rect 251692 305396 251698 305448
rect 253014 305396 253020 305448
rect 253072 305436 253078 305448
rect 253842 305436 253848 305448
rect 253072 305408 253848 305436
rect 253072 305396 253078 305408
rect 253842 305396 253848 305408
rect 253900 305396 253906 305448
rect 254026 305396 254032 305448
rect 254084 305436 254090 305448
rect 254762 305436 254768 305448
rect 254084 305408 254768 305436
rect 254084 305396 254090 305408
rect 254762 305396 254768 305408
rect 254820 305396 254826 305448
rect 255682 305396 255688 305448
rect 255740 305436 255746 305448
rect 256326 305436 256332 305448
rect 255740 305408 256332 305436
rect 255740 305396 255746 305408
rect 256326 305396 256332 305408
rect 256384 305396 256390 305448
rect 257154 305396 257160 305448
rect 257212 305436 257218 305448
rect 257982 305436 257988 305448
rect 257212 305408 257988 305436
rect 257212 305396 257218 305408
rect 257982 305396 257988 305408
rect 258040 305396 258046 305448
rect 260834 305396 260840 305448
rect 260892 305436 260898 305448
rect 261294 305436 261300 305448
rect 260892 305408 261300 305436
rect 260892 305396 260898 305408
rect 261294 305396 261300 305408
rect 261352 305396 261358 305448
rect 263778 305396 263784 305448
rect 263836 305436 263842 305448
rect 264514 305436 264520 305448
rect 263836 305408 264520 305436
rect 263836 305396 263842 305408
rect 264514 305396 264520 305408
rect 264572 305396 264578 305448
rect 265066 305396 265072 305448
rect 265124 305436 265130 305448
rect 265618 305436 265624 305448
rect 265124 305408 265624 305436
rect 265124 305396 265130 305408
rect 265618 305396 265624 305408
rect 265676 305396 265682 305448
rect 269666 305396 269672 305448
rect 269724 305436 269730 305448
rect 270218 305436 270224 305448
rect 269724 305408 270224 305436
rect 269724 305396 269730 305408
rect 270218 305396 270224 305408
rect 270276 305396 270282 305448
rect 270770 305396 270776 305448
rect 270828 305436 270834 305448
rect 271414 305436 271420 305448
rect 270828 305408 271420 305436
rect 270828 305396 270834 305408
rect 271414 305396 271420 305408
rect 271472 305396 271478 305448
rect 276198 305396 276204 305448
rect 276256 305436 276262 305448
rect 277302 305436 277308 305448
rect 276256 305408 277308 305436
rect 276256 305396 276262 305408
rect 277302 305396 277308 305408
rect 277360 305396 277366 305448
rect 280154 305396 280160 305448
rect 280212 305436 280218 305448
rect 280522 305436 280528 305448
rect 280212 305408 280528 305436
rect 280212 305396 280218 305408
rect 280522 305396 280528 305408
rect 280580 305396 280586 305448
rect 350902 305396 350908 305448
rect 350960 305436 350966 305448
rect 362034 305436 362040 305448
rect 350960 305408 362040 305436
rect 350960 305396 350966 305408
rect 362034 305396 362040 305408
rect 362092 305396 362098 305448
rect 255498 305328 255504 305380
rect 255556 305368 255562 305380
rect 256510 305368 256516 305380
rect 255556 305340 256516 305368
rect 255556 305328 255562 305340
rect 256510 305328 256516 305340
rect 256568 305328 256574 305380
rect 261110 305328 261116 305380
rect 261168 305368 261174 305380
rect 262030 305368 262036 305380
rect 261168 305340 262036 305368
rect 261168 305328 261174 305340
rect 262030 305328 262036 305340
rect 262088 305328 262094 305380
rect 269298 305328 269304 305380
rect 269356 305368 269362 305380
rect 270402 305368 270408 305380
rect 269356 305340 270408 305368
rect 269356 305328 269362 305340
rect 270402 305328 270408 305340
rect 270460 305328 270466 305380
rect 270586 305328 270592 305380
rect 270644 305368 270650 305380
rect 271782 305368 271788 305380
rect 270644 305340 271788 305368
rect 270644 305328 270650 305340
rect 271782 305328 271788 305340
rect 271840 305328 271846 305380
rect 275830 305328 275836 305380
rect 275888 305368 275894 305380
rect 281534 305368 281540 305380
rect 275888 305340 281540 305368
rect 275888 305328 275894 305340
rect 281534 305328 281540 305340
rect 281592 305328 281598 305380
rect 360286 305328 360292 305380
rect 360344 305368 360350 305380
rect 368842 305368 368848 305380
rect 360344 305340 368848 305368
rect 360344 305328 360350 305340
rect 368842 305328 368848 305340
rect 368900 305328 368906 305380
rect 260834 305260 260840 305312
rect 260892 305300 260898 305312
rect 261846 305300 261852 305312
rect 260892 305272 261852 305300
rect 260892 305260 260898 305272
rect 261846 305260 261852 305272
rect 261904 305260 261910 305312
rect 360194 305260 360200 305312
rect 360252 305300 360258 305312
rect 368750 305300 368756 305312
rect 360252 305272 368756 305300
rect 360252 305260 360258 305272
rect 368750 305260 368756 305272
rect 368808 305260 368814 305312
rect 97258 305056 97264 305108
rect 97316 305096 97322 305108
rect 97534 305096 97540 305108
rect 97316 305068 97540 305096
rect 97316 305056 97322 305068
rect 97534 305056 97540 305068
rect 97592 305056 97598 305108
rect 97534 304920 97540 304972
rect 97592 304960 97598 304972
rect 97902 304960 97908 304972
rect 97592 304932 97908 304960
rect 97592 304920 97598 304932
rect 97902 304920 97908 304932
rect 97960 304920 97966 304972
rect 172330 304920 172336 304972
rect 172388 304960 172394 304972
rect 245194 304960 245200 304972
rect 172388 304932 245200 304960
rect 172388 304920 172394 304932
rect 245194 304920 245200 304932
rect 245252 304920 245258 304972
rect 314654 304648 314660 304700
rect 314712 304688 314718 304700
rect 315666 304688 315672 304700
rect 314712 304660 315672 304688
rect 314712 304648 314718 304660
rect 315666 304648 315672 304660
rect 315724 304648 315730 304700
rect 170030 304580 170036 304632
rect 170088 304620 170094 304632
rect 240042 304620 240048 304632
rect 170088 304592 240048 304620
rect 170088 304580 170094 304592
rect 240042 304580 240048 304592
rect 240100 304580 240106 304632
rect 171962 304512 171968 304564
rect 172020 304552 172026 304564
rect 245470 304552 245476 304564
rect 172020 304524 245476 304552
rect 172020 304512 172026 304524
rect 245470 304512 245476 304524
rect 245528 304512 245534 304564
rect 172238 304444 172244 304496
rect 172296 304484 172302 304496
rect 248874 304484 248880 304496
rect 172296 304456 248880 304484
rect 172296 304444 172302 304456
rect 248874 304444 248880 304456
rect 248932 304444 248938 304496
rect 207014 304376 207020 304428
rect 207072 304416 207078 304428
rect 285766 304416 285772 304428
rect 207072 304388 285772 304416
rect 207072 304376 207078 304388
rect 285766 304376 285772 304388
rect 285824 304376 285830 304428
rect 326430 304376 326436 304428
rect 326488 304416 326494 304428
rect 452654 304416 452660 304428
rect 326488 304388 452660 304416
rect 326488 304376 326494 304388
rect 452654 304376 452660 304388
rect 452712 304376 452718 304428
rect 171778 304308 171784 304360
rect 171836 304348 171842 304360
rect 256694 304348 256700 304360
rect 171836 304320 256700 304348
rect 171836 304308 171842 304320
rect 256694 304308 256700 304320
rect 256752 304308 256758 304360
rect 256878 304308 256884 304360
rect 256936 304348 256942 304360
rect 257062 304348 257068 304360
rect 256936 304320 257068 304348
rect 256936 304308 256942 304320
rect 257062 304308 257068 304320
rect 257120 304308 257126 304360
rect 263502 304308 263508 304360
rect 263560 304348 263566 304360
rect 263686 304348 263692 304360
rect 263560 304320 263692 304348
rect 263560 304308 263566 304320
rect 263686 304308 263692 304320
rect 263744 304308 263750 304360
rect 331766 304308 331772 304360
rect 331824 304348 331830 304360
rect 485038 304348 485044 304360
rect 331824 304320 485044 304348
rect 331824 304308 331830 304320
rect 485038 304308 485044 304320
rect 485096 304308 485102 304360
rect 189074 304240 189080 304292
rect 189132 304280 189138 304292
rect 283006 304280 283012 304292
rect 189132 304252 283012 304280
rect 189132 304240 189138 304252
rect 283006 304240 283012 304252
rect 283064 304240 283070 304292
rect 335906 304240 335912 304292
rect 335964 304280 335970 304292
rect 514018 304280 514024 304292
rect 335964 304252 514024 304280
rect 335964 304240 335970 304252
rect 514018 304240 514024 304252
rect 514076 304240 514082 304292
rect 256602 304172 256608 304224
rect 256660 304212 256666 304224
rect 256970 304212 256976 304224
rect 256660 304184 256976 304212
rect 256660 304172 256666 304184
rect 256970 304172 256976 304184
rect 257028 304172 257034 304224
rect 274818 303968 274824 304020
rect 274876 304008 274882 304020
rect 275922 304008 275928 304020
rect 274876 303980 275928 304008
rect 274876 303968 274882 303980
rect 275922 303968 275928 303980
rect 275980 303968 275986 304020
rect 302510 303968 302516 304020
rect 302568 304008 302574 304020
rect 303430 304008 303436 304020
rect 302568 303980 303436 304008
rect 302568 303968 302574 303980
rect 303430 303968 303436 303980
rect 303488 303968 303494 304020
rect 300946 303696 300952 303748
rect 301004 303736 301010 303748
rect 301866 303736 301872 303748
rect 301004 303708 301872 303736
rect 301004 303696 301010 303708
rect 301866 303696 301872 303708
rect 301924 303696 301930 303748
rect 342438 303696 342444 303748
rect 342496 303736 342502 303748
rect 343358 303736 343364 303748
rect 342496 303708 343364 303736
rect 342496 303696 342502 303708
rect 343358 303696 343364 303708
rect 343416 303696 343422 303748
rect 214650 303560 214656 303612
rect 214708 303600 214714 303612
rect 288434 303600 288440 303612
rect 214708 303572 288440 303600
rect 214708 303560 214714 303572
rect 288434 303560 288440 303572
rect 288492 303560 288498 303612
rect 344002 303560 344008 303612
rect 344060 303600 344066 303612
rect 344462 303600 344468 303612
rect 344060 303572 344468 303600
rect 344060 303560 344066 303572
rect 344462 303560 344468 303572
rect 344520 303560 344526 303612
rect 356054 303560 356060 303612
rect 356112 303600 356118 303612
rect 373442 303600 373448 303612
rect 356112 303572 373448 303600
rect 356112 303560 356118 303572
rect 373442 303560 373448 303572
rect 373500 303560 373506 303612
rect 215938 303492 215944 303544
rect 215996 303532 216002 303544
rect 290826 303532 290832 303544
rect 215996 303504 290832 303532
rect 215996 303492 216002 303504
rect 290826 303492 290832 303504
rect 290884 303492 290890 303544
rect 316126 303492 316132 303544
rect 316184 303532 316190 303544
rect 316954 303532 316960 303544
rect 316184 303504 316960 303532
rect 316184 303492 316190 303504
rect 316954 303492 316960 303504
rect 317012 303492 317018 303544
rect 350718 303492 350724 303544
rect 350776 303532 350782 303544
rect 370682 303532 370688 303544
rect 350776 303504 370688 303532
rect 350776 303492 350782 303504
rect 370682 303492 370688 303504
rect 370740 303492 370746 303544
rect 169938 303424 169944 303476
rect 169996 303464 170002 303476
rect 246022 303464 246028 303476
rect 169996 303436 246028 303464
rect 169996 303424 170002 303436
rect 246022 303424 246028 303436
rect 246080 303424 246086 303476
rect 352006 303424 352012 303476
rect 352064 303464 352070 303476
rect 372982 303464 372988 303476
rect 352064 303436 372988 303464
rect 352064 303424 352070 303436
rect 372982 303424 372988 303436
rect 373040 303424 373046 303476
rect 217962 303356 217968 303408
rect 218020 303396 218026 303408
rect 293218 303396 293224 303408
rect 218020 303368 293224 303396
rect 218020 303356 218026 303368
rect 293218 303356 293224 303368
rect 293276 303356 293282 303408
rect 352098 303356 352104 303408
rect 352156 303396 352162 303408
rect 373074 303396 373080 303408
rect 352156 303368 373080 303396
rect 352156 303356 352162 303368
rect 373074 303356 373080 303368
rect 373132 303356 373138 303408
rect 214742 303288 214748 303340
rect 214800 303328 214806 303340
rect 289906 303328 289912 303340
rect 214800 303300 289912 303328
rect 214800 303288 214806 303300
rect 289906 303288 289912 303300
rect 289964 303288 289970 303340
rect 348694 303288 348700 303340
rect 348752 303328 348758 303340
rect 370222 303328 370228 303340
rect 348752 303300 370228 303328
rect 348752 303288 348758 303300
rect 370222 303288 370228 303300
rect 370280 303288 370286 303340
rect 216030 303220 216036 303272
rect 216088 303260 216094 303272
rect 291194 303260 291200 303272
rect 216088 303232 291200 303260
rect 216088 303220 216094 303232
rect 291194 303220 291200 303232
rect 291252 303220 291258 303272
rect 350626 303220 350632 303272
rect 350684 303260 350690 303272
rect 372890 303260 372896 303272
rect 350684 303232 372896 303260
rect 350684 303220 350690 303232
rect 372890 303220 372896 303232
rect 372948 303220 372954 303272
rect 215018 303152 215024 303204
rect 215076 303192 215082 303204
rect 291378 303192 291384 303204
rect 215076 303164 291384 303192
rect 215076 303152 215082 303164
rect 291378 303152 291384 303164
rect 291436 303152 291442 303204
rect 349614 303152 349620 303204
rect 349672 303192 349678 303204
rect 373166 303192 373172 303204
rect 349672 303164 373172 303192
rect 349672 303152 349678 303164
rect 373166 303152 373172 303164
rect 373224 303152 373230 303204
rect 214558 303084 214564 303136
rect 214616 303124 214622 303136
rect 292574 303124 292580 303136
rect 214616 303096 292580 303124
rect 214616 303084 214622 303096
rect 292574 303084 292580 303096
rect 292632 303084 292638 303136
rect 347958 303084 347964 303136
rect 348016 303124 348022 303136
rect 372062 303124 372068 303136
rect 348016 303096 372068 303124
rect 348016 303084 348022 303096
rect 372062 303084 372068 303096
rect 372120 303084 372126 303136
rect 219158 303016 219164 303068
rect 219216 303056 219222 303068
rect 299014 303056 299020 303068
rect 219216 303028 299020 303056
rect 219216 303016 219222 303028
rect 299014 303016 299020 303028
rect 299072 303016 299078 303068
rect 348878 303016 348884 303068
rect 348936 303056 348942 303068
rect 373350 303056 373356 303068
rect 348936 303028 373356 303056
rect 348936 303016 348942 303028
rect 373350 303016 373356 303028
rect 373408 303016 373414 303068
rect 169754 302948 169760 303000
rect 169812 302988 169818 303000
rect 251542 302988 251548 303000
rect 169812 302960 251548 302988
rect 169812 302948 169818 302960
rect 251542 302948 251548 302960
rect 251600 302948 251606 303000
rect 301222 302948 301228 303000
rect 301280 302988 301286 303000
rect 363598 302988 363604 303000
rect 301280 302960 363604 302988
rect 301280 302948 301286 302960
rect 363598 302948 363604 302960
rect 363656 302948 363662 303000
rect 212166 302880 212172 302932
rect 212224 302920 212230 302932
rect 294506 302920 294512 302932
rect 212224 302892 294512 302920
rect 212224 302880 212230 302892
rect 294506 302880 294512 302892
rect 294564 302880 294570 302932
rect 299382 302880 299388 302932
rect 299440 302920 299446 302932
rect 365162 302920 365168 302932
rect 299440 302892 365168 302920
rect 299440 302880 299446 302892
rect 365162 302880 365168 302892
rect 365220 302880 365226 302932
rect 215110 302812 215116 302864
rect 215168 302852 215174 302864
rect 288618 302852 288624 302864
rect 215168 302824 288624 302852
rect 215168 302812 215174 302824
rect 288618 302812 288624 302824
rect 288676 302812 288682 302864
rect 303706 302812 303712 302864
rect 303764 302852 303770 302864
rect 304534 302852 304540 302864
rect 303764 302824 304540 302852
rect 303764 302812 303770 302824
rect 304534 302812 304540 302824
rect 304592 302812 304598 302864
rect 327166 302812 327172 302864
rect 327224 302852 327230 302864
rect 327902 302852 327908 302864
rect 327224 302824 327908 302852
rect 327224 302812 327230 302824
rect 327902 302812 327908 302824
rect 327960 302812 327966 302864
rect 349430 302812 349436 302864
rect 349488 302852 349494 302864
rect 366542 302852 366548 302864
rect 349488 302824 366548 302852
rect 349488 302812 349494 302824
rect 366542 302812 366548 302824
rect 366600 302812 366606 302864
rect 215846 302744 215852 302796
rect 215904 302784 215910 302796
rect 288802 302784 288808 302796
rect 215904 302756 288808 302784
rect 215904 302744 215910 302756
rect 288802 302744 288808 302756
rect 288860 302744 288866 302796
rect 352558 302744 352564 302796
rect 352616 302784 352622 302796
rect 369118 302784 369124 302796
rect 352616 302756 369124 302784
rect 352616 302744 352622 302756
rect 369118 302744 369124 302756
rect 369176 302744 369182 302796
rect 216490 302676 216496 302728
rect 216548 302716 216554 302728
rect 289170 302716 289176 302728
rect 216548 302688 289176 302716
rect 216548 302676 216554 302688
rect 289170 302676 289176 302688
rect 289228 302676 289234 302728
rect 350166 302676 350172 302728
rect 350224 302716 350230 302728
rect 363690 302716 363696 302728
rect 350224 302688 363696 302716
rect 350224 302676 350230 302688
rect 363690 302676 363696 302688
rect 363748 302676 363754 302728
rect 247678 302608 247684 302660
rect 247736 302648 247742 302660
rect 247954 302648 247960 302660
rect 247736 302620 247960 302648
rect 247736 302608 247742 302620
rect 247954 302608 247960 302620
rect 248012 302608 248018 302660
rect 329926 302608 329932 302660
rect 329984 302648 329990 302660
rect 330294 302648 330300 302660
rect 329984 302620 330300 302648
rect 329984 302608 329990 302620
rect 330294 302608 330300 302620
rect 330352 302608 330358 302660
rect 297174 302472 297180 302524
rect 297232 302512 297238 302524
rect 297910 302512 297916 302524
rect 297232 302484 297916 302512
rect 297232 302472 297238 302484
rect 297910 302472 297916 302484
rect 297968 302472 297974 302524
rect 345106 302336 345112 302388
rect 345164 302376 345170 302388
rect 345842 302376 345848 302388
rect 345164 302348 345848 302376
rect 345164 302336 345170 302348
rect 345842 302336 345848 302348
rect 345900 302336 345906 302388
rect 262306 302268 262312 302320
rect 262364 302308 262370 302320
rect 262364 302280 262812 302308
rect 262364 302268 262370 302280
rect 262784 302252 262812 302280
rect 262766 302200 262772 302252
rect 262824 302200 262830 302252
rect 172422 302132 172428 302184
rect 172480 302172 172486 302184
rect 240410 302172 240416 302184
rect 172480 302144 240416 302172
rect 172480 302132 172486 302144
rect 240410 302132 240416 302144
rect 240468 302132 240474 302184
rect 216214 302064 216220 302116
rect 216272 302104 216278 302116
rect 293126 302104 293132 302116
rect 216272 302076 293132 302104
rect 216272 302064 216278 302076
rect 293126 302064 293132 302076
rect 293184 302064 293190 302116
rect 216122 301996 216128 302048
rect 216180 302036 216186 302048
rect 296806 302036 296812 302048
rect 216180 302008 296812 302036
rect 216180 301996 216186 302008
rect 296806 301996 296812 302008
rect 296864 301996 296870 302048
rect 212442 301928 212448 301980
rect 212500 301968 212506 301980
rect 296530 301968 296536 301980
rect 212500 301940 296536 301968
rect 212500 301928 212506 301940
rect 296530 301928 296536 301940
rect 296588 301928 296594 301980
rect 212258 301860 212264 301912
rect 212316 301900 212322 301912
rect 296714 301900 296720 301912
rect 212316 301872 296720 301900
rect 212316 301860 212322 301872
rect 296714 301860 296720 301872
rect 296772 301860 296778 301912
rect 211062 301792 211068 301844
rect 211120 301832 211126 301844
rect 295518 301832 295524 301844
rect 211120 301804 295524 301832
rect 211120 301792 211126 301804
rect 295518 301792 295524 301804
rect 295576 301792 295582 301844
rect 210786 301724 210792 301776
rect 210844 301764 210850 301776
rect 295426 301764 295432 301776
rect 210844 301736 295432 301764
rect 210844 301724 210850 301736
rect 295426 301724 295432 301736
rect 295484 301724 295490 301776
rect 312262 301724 312268 301776
rect 312320 301764 312326 301776
rect 374086 301764 374092 301776
rect 312320 301736 374092 301764
rect 312320 301724 312326 301736
rect 374086 301724 374092 301736
rect 374144 301724 374150 301776
rect 218422 301656 218428 301708
rect 218480 301696 218486 301708
rect 349798 301696 349804 301708
rect 218480 301668 349804 301696
rect 218480 301656 218486 301668
rect 349798 301656 349804 301668
rect 349856 301656 349862 301708
rect 211706 301588 211712 301640
rect 211764 301628 211770 301640
rect 347958 301628 347964 301640
rect 211764 301600 347964 301628
rect 211764 301588 211770 301600
rect 347958 301588 347964 301600
rect 348016 301588 348022 301640
rect 210878 301520 210884 301572
rect 210936 301560 210942 301572
rect 295610 301560 295616 301572
rect 210936 301532 295616 301560
rect 210936 301520 210942 301532
rect 295610 301520 295616 301532
rect 295668 301520 295674 301572
rect 331582 301520 331588 301572
rect 331640 301560 331646 301572
rect 494054 301560 494060 301572
rect 331640 301532 494060 301560
rect 331640 301520 331646 301532
rect 494054 301520 494060 301532
rect 494112 301520 494118 301572
rect 193214 301452 193220 301504
rect 193272 301492 193278 301504
rect 282914 301492 282920 301504
rect 193272 301464 282920 301492
rect 193272 301452 193278 301464
rect 282914 301452 282920 301464
rect 282972 301452 282978 301504
rect 338666 301452 338672 301504
rect 338724 301492 338730 301504
rect 529934 301492 529940 301504
rect 338724 301464 529940 301492
rect 338724 301452 338730 301464
rect 529934 301452 529940 301464
rect 529992 301452 529998 301504
rect 97350 300772 97356 300824
rect 97408 300812 97414 300824
rect 249886 300812 249892 300824
rect 97408 300784 249892 300812
rect 97408 300772 97414 300784
rect 249886 300772 249892 300784
rect 249944 300772 249950 300824
rect 98638 300704 98644 300756
rect 98696 300744 98702 300756
rect 251358 300744 251364 300756
rect 98696 300716 251364 300744
rect 98696 300704 98702 300716
rect 251358 300704 251364 300716
rect 251416 300704 251422 300756
rect 97718 300636 97724 300688
rect 97776 300676 97782 300688
rect 246206 300676 246212 300688
rect 97776 300648 246212 300676
rect 97776 300636 97782 300648
rect 246206 300636 246212 300648
rect 246264 300636 246270 300688
rect 97810 300568 97816 300620
rect 97868 300608 97874 300620
rect 242802 300608 242808 300620
rect 97868 300580 242808 300608
rect 97868 300568 97874 300580
rect 242802 300568 242808 300580
rect 242860 300568 242866 300620
rect 296990 300568 296996 300620
rect 297048 300608 297054 300620
rect 297358 300608 297364 300620
rect 297048 300580 297364 300608
rect 297048 300568 297054 300580
rect 297358 300568 297364 300580
rect 297416 300568 297422 300620
rect 99098 300500 99104 300552
rect 99156 300540 99162 300552
rect 243078 300540 243084 300552
rect 99156 300512 243084 300540
rect 99156 300500 99162 300512
rect 243078 300500 243084 300512
rect 243136 300500 243142 300552
rect 97626 300432 97632 300484
rect 97684 300472 97690 300484
rect 242710 300472 242716 300484
rect 97684 300444 242716 300472
rect 97684 300432 97690 300444
rect 242710 300432 242716 300444
rect 242768 300432 242774 300484
rect 300210 300432 300216 300484
rect 300268 300472 300274 300484
rect 362310 300472 362316 300484
rect 300268 300444 362316 300472
rect 300268 300432 300274 300444
rect 362310 300432 362316 300444
rect 362368 300432 362374 300484
rect 99374 300364 99380 300416
rect 99432 300404 99438 300416
rect 240318 300404 240324 300416
rect 99432 300376 240324 300404
rect 99432 300364 99438 300376
rect 240318 300364 240324 300376
rect 240376 300364 240382 300416
rect 313826 300364 313832 300416
rect 313884 300404 313890 300416
rect 376754 300404 376760 300416
rect 313884 300376 376760 300404
rect 313884 300364 313890 300376
rect 376754 300364 376760 300376
rect 376812 300364 376818 300416
rect 99558 300296 99564 300348
rect 99616 300336 99622 300348
rect 240134 300336 240140 300348
rect 99616 300308 240140 300336
rect 99616 300296 99622 300308
rect 240134 300296 240140 300308
rect 240192 300296 240198 300348
rect 301222 300296 301228 300348
rect 301280 300336 301286 300348
rect 370590 300336 370596 300348
rect 301280 300308 370596 300336
rect 301280 300296 301286 300308
rect 370590 300296 370596 300308
rect 370648 300296 370654 300348
rect 99834 300228 99840 300280
rect 99892 300268 99898 300280
rect 238938 300268 238944 300280
rect 99892 300240 238944 300268
rect 99892 300228 99898 300240
rect 238938 300228 238944 300240
rect 238996 300228 239002 300280
rect 327626 300228 327632 300280
rect 327684 300268 327690 300280
rect 463694 300268 463700 300280
rect 327684 300240 463700 300268
rect 327684 300228 327690 300240
rect 463694 300228 463700 300240
rect 463752 300228 463758 300280
rect 99190 300160 99196 300212
rect 99248 300200 99254 300212
rect 237742 300200 237748 300212
rect 99248 300172 237748 300200
rect 99248 300160 99254 300172
rect 237742 300160 237748 300172
rect 237800 300160 237806 300212
rect 333146 300160 333152 300212
rect 333204 300200 333210 300212
rect 498286 300200 498292 300212
rect 333204 300172 498292 300200
rect 333204 300160 333210 300172
rect 498286 300160 498292 300172
rect 498344 300160 498350 300212
rect 99466 300092 99472 300144
rect 99524 300132 99530 300144
rect 236178 300132 236184 300144
rect 99524 300104 236184 300132
rect 99524 300092 99530 300104
rect 236178 300092 236184 300104
rect 236236 300092 236242 300144
rect 339954 300092 339960 300144
rect 340012 300132 340018 300144
rect 538858 300132 538864 300144
rect 340012 300104 538864 300132
rect 340012 300092 340018 300104
rect 538858 300092 538864 300104
rect 538916 300092 538922 300144
rect 210602 300024 210608 300076
rect 210660 300064 210666 300076
rect 347866 300064 347872 300076
rect 210660 300036 347872 300064
rect 210660 300024 210666 300036
rect 347866 300024 347872 300036
rect 347924 300024 347930 300076
rect 99006 299956 99012 300008
rect 99064 299996 99070 300008
rect 233326 299996 233332 300008
rect 99064 299968 233332 299996
rect 99064 299956 99070 299968
rect 233326 299956 233332 299968
rect 233384 299956 233390 300008
rect 217778 299888 217784 299940
rect 217836 299928 217842 299940
rect 348970 299928 348976 299940
rect 217836 299900 348976 299928
rect 217836 299888 217842 299900
rect 348970 299888 348976 299900
rect 349028 299888 349034 299940
rect 305546 299684 305552 299736
rect 305604 299724 305610 299736
rect 305914 299724 305920 299736
rect 305604 299696 305920 299724
rect 305604 299684 305610 299696
rect 305914 299684 305920 299696
rect 305972 299684 305978 299736
rect 98822 299412 98828 299464
rect 98880 299452 98886 299464
rect 247310 299452 247316 299464
rect 98880 299424 247316 299452
rect 98880 299412 98886 299424
rect 247310 299412 247316 299424
rect 247368 299412 247374 299464
rect 97902 299344 97908 299396
rect 97960 299384 97966 299396
rect 242986 299384 242992 299396
rect 97960 299356 242992 299384
rect 97960 299344 97966 299356
rect 242986 299344 242992 299356
rect 243044 299344 243050 299396
rect 99742 299276 99748 299328
rect 99800 299316 99806 299328
rect 240226 299316 240232 299328
rect 99800 299288 240232 299316
rect 99800 299276 99806 299288
rect 240226 299276 240232 299288
rect 240284 299276 240290 299328
rect 98914 299208 98920 299260
rect 98972 299248 98978 299260
rect 238018 299248 238024 299260
rect 98972 299220 238024 299248
rect 98972 299208 98978 299220
rect 238018 299208 238024 299220
rect 238076 299208 238082 299260
rect 114830 299140 114836 299192
rect 114888 299180 114894 299192
rect 244458 299180 244464 299192
rect 114888 299152 244464 299180
rect 114888 299140 114894 299152
rect 244458 299140 244464 299152
rect 244516 299140 244522 299192
rect 119982 299072 119988 299124
rect 120040 299112 120046 299124
rect 247126 299112 247132 299124
rect 120040 299084 247132 299112
rect 120040 299072 120046 299084
rect 247126 299072 247132 299084
rect 247184 299072 247190 299124
rect 130286 299004 130292 299056
rect 130344 299044 130350 299056
rect 249978 299044 249984 299056
rect 130344 299016 249984 299044
rect 130344 299004 130350 299016
rect 249978 299004 249984 299016
rect 250036 299004 250042 299056
rect 313642 299004 313648 299056
rect 313700 299044 313706 299056
rect 378134 299044 378140 299056
rect 313700 299016 378140 299044
rect 313700 299004 313706 299016
rect 378134 299004 378140 299016
rect 378192 299004 378198 299056
rect 125134 298936 125140 298988
rect 125192 298976 125198 298988
rect 238846 298976 238852 298988
rect 125192 298948 238852 298976
rect 125192 298936 125198 298948
rect 238846 298936 238852 298948
rect 238904 298936 238910 298988
rect 315114 298936 315120 298988
rect 315172 298976 315178 298988
rect 381538 298976 381544 298988
rect 315172 298948 381544 298976
rect 315172 298936 315178 298948
rect 381538 298936 381544 298948
rect 381596 298936 381602 298988
rect 140590 298868 140596 298920
rect 140648 298908 140654 298920
rect 250622 298908 250628 298920
rect 140648 298880 250628 298908
rect 140648 298868 140654 298880
rect 250622 298868 250628 298880
rect 250680 298868 250686 298920
rect 333054 298868 333060 298920
rect 333112 298908 333118 298920
rect 500218 298908 500224 298920
rect 333112 298880 500224 298908
rect 333112 298868 333118 298880
rect 500218 298868 500224 298880
rect 500276 298868 500282 298920
rect 143442 298800 143448 298852
rect 143500 298840 143506 298852
rect 248506 298840 248512 298852
rect 143500 298812 248512 298840
rect 143500 298800 143506 298812
rect 248506 298800 248512 298812
rect 248564 298800 248570 298852
rect 341426 298800 341432 298852
rect 341484 298840 341490 298852
rect 547966 298840 547972 298852
rect 341484 298812 547972 298840
rect 341484 298800 341490 298812
rect 547966 298800 547972 298812
rect 548024 298800 548030 298852
rect 133782 298732 133788 298784
rect 133840 298772 133846 298784
rect 243170 298772 243176 298784
rect 133840 298744 243176 298772
rect 133840 298732 133846 298744
rect 243170 298732 243176 298744
rect 243228 298732 243234 298784
rect 344830 298732 344836 298784
rect 344888 298772 344894 298784
rect 567838 298772 567844 298784
rect 344888 298744 567844 298772
rect 344888 298732 344894 298744
rect 567838 298732 567844 298744
rect 567896 298732 567902 298784
rect 156046 298664 156052 298716
rect 156104 298704 156110 298716
rect 251726 298704 251732 298716
rect 156104 298676 251732 298704
rect 156104 298664 156110 298676
rect 251726 298664 251732 298676
rect 251784 298664 251790 298716
rect 161198 298596 161204 298648
rect 161256 298636 161262 298648
rect 247770 298636 247776 298648
rect 161256 298608 247776 298636
rect 161256 298596 161262 298608
rect 247770 298596 247776 298608
rect 247828 298596 247834 298648
rect 163774 298528 163780 298580
rect 163832 298568 163838 298580
rect 234706 298568 234712 298580
rect 163832 298540 234712 298568
rect 163832 298528 163838 298540
rect 234706 298528 234712 298540
rect 234764 298528 234770 298580
rect 107102 298052 107108 298104
rect 107160 298092 107166 298104
rect 111150 298092 111156 298104
rect 107160 298064 111156 298092
rect 107160 298052 107166 298064
rect 111150 298052 111156 298064
rect 111208 298052 111214 298104
rect 166350 298052 166356 298104
rect 166408 298092 166414 298104
rect 170582 298092 170588 298104
rect 166408 298064 170588 298092
rect 166408 298052 166414 298064
rect 170582 298052 170588 298064
rect 170640 298052 170646 298104
rect 117406 297984 117412 298036
rect 117464 298024 117470 298036
rect 133782 298024 133788 298036
rect 117464 297996 133788 298024
rect 117464 297984 117470 297996
rect 133782 297984 133788 297996
rect 133840 297984 133846 298036
rect 158622 297984 158628 298036
rect 158680 298024 158686 298036
rect 169846 298024 169852 298036
rect 158680 297996 169852 298024
rect 158680 297984 158686 297996
rect 169846 297984 169852 297996
rect 169904 297984 169910 298036
rect 122558 297916 122564 297968
rect 122616 297956 122622 297968
rect 237650 297956 237656 297968
rect 122616 297928 237656 297956
rect 122616 297916 122622 297928
rect 237650 297916 237656 297928
rect 237708 297916 237714 297968
rect 138014 297848 138020 297900
rect 138072 297888 138078 297900
rect 239030 297888 239036 297900
rect 138072 297860 239036 297888
rect 138072 297848 138078 297860
rect 239030 297848 239036 297860
rect 239088 297848 239094 297900
rect 127710 297780 127716 297832
rect 127768 297820 127774 297832
rect 143442 297820 143448 297832
rect 127768 297792 143448 297820
rect 127768 297780 127774 297792
rect 143442 297780 143448 297792
rect 143500 297780 143506 297832
rect 148318 297780 148324 297832
rect 148376 297820 148382 297832
rect 236362 297820 236368 297832
rect 148376 297792 236368 297820
rect 148376 297780 148382 297792
rect 236362 297780 236368 297792
rect 236420 297780 236426 297832
rect 100018 297712 100024 297764
rect 100076 297752 100082 297764
rect 169938 297752 169944 297764
rect 100076 297724 169944 297752
rect 100076 297712 100082 297724
rect 169938 297712 169944 297724
rect 169996 297712 170002 297764
rect 213454 297712 213460 297764
rect 213512 297752 213518 297764
rect 293034 297752 293040 297764
rect 213512 297724 293040 297752
rect 213512 297712 213518 297724
rect 293034 297712 293040 297724
rect 293092 297712 293098 297764
rect 109678 297644 109684 297696
rect 109736 297684 109742 297696
rect 109736 297656 171134 297684
rect 109736 297644 109742 297656
rect 135438 297576 135444 297628
rect 135496 297616 135502 297628
rect 171106 297616 171134 297656
rect 214466 297644 214472 297696
rect 214524 297684 214530 297696
rect 294138 297684 294144 297696
rect 214524 297656 294144 297684
rect 214524 297644 214530 297656
rect 294138 297644 294144 297656
rect 294196 297644 294202 297696
rect 322198 297644 322204 297696
rect 322256 297684 322262 297696
rect 381630 297684 381636 297696
rect 322256 297656 381636 297684
rect 322256 297644 322262 297656
rect 381630 297644 381636 297656
rect 381688 297644 381694 297696
rect 172238 297616 172244 297628
rect 135496 297588 162900 297616
rect 171106 297588 172244 297616
rect 135496 297576 135502 297588
rect 143166 297508 143172 297560
rect 143224 297548 143230 297560
rect 162872 297548 162900 297588
rect 172238 297576 172244 297588
rect 172296 297576 172302 297628
rect 213822 297576 213828 297628
rect 213880 297616 213886 297628
rect 294414 297616 294420 297628
rect 213880 297588 294420 297616
rect 213880 297576 213886 297588
rect 294414 297576 294420 297588
rect 294472 297576 294478 297628
rect 319254 297576 319260 297628
rect 319312 297616 319318 297628
rect 412634 297616 412640 297628
rect 319312 297588 412640 297616
rect 319312 297576 319318 297588
rect 412634 297576 412640 297588
rect 412692 297576 412698 297628
rect 171962 297548 171968 297560
rect 143224 297520 161612 297548
rect 162872 297520 171968 297548
rect 143224 297508 143230 297520
rect 150894 297440 150900 297492
rect 150952 297480 150958 297492
rect 150952 297452 161474 297480
rect 150952 297440 150958 297452
rect 161446 297344 161474 297452
rect 161584 297412 161612 297520
rect 171962 297508 171968 297520
rect 172020 297508 172026 297560
rect 213178 297508 213184 297560
rect 213236 297548 213242 297560
rect 346578 297548 346584 297560
rect 213236 297520 346584 297548
rect 213236 297508 213242 297520
rect 346578 297508 346584 297520
rect 346636 297508 346642 297560
rect 213730 297440 213736 297492
rect 213788 297480 213794 297492
rect 294690 297480 294696 297492
rect 213788 297452 294696 297480
rect 213788 297440 213794 297452
rect 294690 297440 294696 297452
rect 294748 297440 294754 297492
rect 342806 297440 342812 297492
rect 342864 297480 342870 297492
rect 556154 297480 556160 297492
rect 342864 297452 556160 297480
rect 342864 297440 342870 297452
rect 556154 297440 556160 297452
rect 556212 297440 556218 297492
rect 171686 297412 171692 297424
rect 161584 297384 171692 297412
rect 171686 297372 171692 297384
rect 171744 297372 171750 297424
rect 210694 297372 210700 297424
rect 210752 297412 210758 297424
rect 292942 297412 292948 297424
rect 210752 297384 292948 297412
rect 210752 297372 210758 297384
rect 292942 297372 292948 297384
rect 293000 297372 293006 297424
rect 342714 297372 342720 297424
rect 342772 297412 342778 297424
rect 557534 297412 557540 297424
rect 342772 297384 557540 297412
rect 342772 297372 342778 297384
rect 557534 297372 557540 297384
rect 557592 297372 557598 297424
rect 170030 297344 170036 297356
rect 161446 297316 170036 297344
rect 170030 297304 170036 297316
rect 170088 297304 170094 297356
rect 212350 297304 212356 297356
rect 212408 297344 212414 297356
rect 291654 297344 291660 297356
rect 212408 297316 291660 297344
rect 212408 297304 212414 297316
rect 291654 297304 291660 297316
rect 291712 297304 291718 297356
rect 217870 297236 217876 297288
rect 217928 297276 217934 297288
rect 295794 297276 295800 297288
rect 217928 297248 295800 297276
rect 217928 297236 217934 297248
rect 295794 297236 295800 297248
rect 295852 297236 295858 297288
rect 218790 297168 218796 297220
rect 218848 297208 218854 297220
rect 294230 297208 294236 297220
rect 218848 297180 294236 297208
rect 218848 297168 218854 297180
rect 294230 297168 294236 297180
rect 294288 297168 294294 297220
rect 112254 297100 112260 297152
rect 112312 297140 112318 297152
rect 235902 297140 235908 297152
rect 112312 297112 235908 297140
rect 112312 297100 112318 297112
rect 235902 297100 235908 297112
rect 235960 297100 235966 297152
rect 132862 297032 132868 297084
rect 132920 297072 132926 297084
rect 251450 297072 251456 297084
rect 132920 297044 251456 297072
rect 132920 297032 132926 297044
rect 251450 297032 251456 297044
rect 251508 297032 251514 297084
rect 98730 296624 98736 296676
rect 98788 296664 98794 296676
rect 240502 296664 240508 296676
rect 98788 296636 240508 296664
rect 98788 296624 98794 296636
rect 240502 296624 240508 296636
rect 240560 296624 240566 296676
rect 103514 296556 103520 296608
rect 103572 296596 103578 296608
rect 234798 296596 234804 296608
rect 103572 296568 234804 296596
rect 103572 296556 103578 296568
rect 234798 296556 234804 296568
rect 234856 296556 234862 296608
rect 111150 296488 111156 296540
rect 111208 296528 111214 296540
rect 236454 296528 236460 296540
rect 111208 296500 236460 296528
rect 111208 296488 111214 296500
rect 236454 296488 236460 296500
rect 236512 296488 236518 296540
rect 153194 296420 153200 296472
rect 153252 296460 153258 296472
rect 248690 296460 248696 296472
rect 153252 296432 248696 296460
rect 153252 296420 153258 296432
rect 248690 296420 248696 296432
rect 248748 296420 248754 296472
rect 312170 296216 312176 296268
rect 312228 296256 312234 296268
rect 372614 296256 372620 296268
rect 312228 296228 372620 296256
rect 312228 296216 312234 296228
rect 372614 296216 372620 296228
rect 372672 296216 372678 296268
rect 322014 296148 322020 296200
rect 322072 296188 322078 296200
rect 421558 296188 421564 296200
rect 322072 296160 421564 296188
rect 322072 296148 322078 296160
rect 421558 296148 421564 296160
rect 421616 296148 421622 296200
rect 209774 296080 209780 296132
rect 209832 296120 209838 296132
rect 285674 296120 285680 296132
rect 209832 296092 285680 296120
rect 209832 296080 209838 296092
rect 285674 296080 285680 296092
rect 285732 296080 285738 296132
rect 320726 296080 320732 296132
rect 320784 296120 320790 296132
rect 422294 296120 422300 296132
rect 320784 296092 422300 296120
rect 320784 296080 320790 296092
rect 422294 296080 422300 296092
rect 422352 296080 422358 296132
rect 129734 296012 129740 296064
rect 129792 296052 129798 296064
rect 273806 296052 273812 296064
rect 129792 296024 273812 296052
rect 129792 296012 129798 296024
rect 273806 296012 273812 296024
rect 273864 296012 273870 296064
rect 335814 296012 335820 296064
rect 335872 296052 335878 296064
rect 516778 296052 516784 296064
rect 335872 296024 516784 296052
rect 335872 296012 335878 296024
rect 516778 296012 516784 296024
rect 516836 296012 516842 296064
rect 125594 295944 125600 295996
rect 125652 295984 125658 295996
rect 272426 295984 272432 295996
rect 125652 295956 272432 295984
rect 125652 295944 125658 295956
rect 272426 295944 272432 295956
rect 272484 295944 272490 295996
rect 344094 295944 344100 295996
rect 344152 295984 344158 295996
rect 563698 295984 563704 295996
rect 344152 295956 563704 295984
rect 344152 295944 344158 295956
rect 563698 295944 563704 295956
rect 563756 295944 563762 295996
rect 219342 295128 219348 295180
rect 219400 295168 219406 295180
rect 295702 295168 295708 295180
rect 219400 295140 295708 295168
rect 219400 295128 219406 295140
rect 295702 295128 295708 295140
rect 295760 295128 295766 295180
rect 209682 295060 209688 295112
rect 209740 295100 209746 295112
rect 287422 295100 287428 295112
rect 209740 295072 287428 295100
rect 209740 295060 209746 295072
rect 287422 295060 287428 295072
rect 287480 295060 287486 295112
rect 214926 294992 214932 295044
rect 214984 295032 214990 295044
rect 294322 295032 294328 295044
rect 214984 295004 294328 295032
rect 214984 294992 214990 295004
rect 294322 294992 294328 295004
rect 294380 294992 294386 295044
rect 215754 294924 215760 294976
rect 215812 294964 215818 294976
rect 296990 294964 296996 294976
rect 215812 294936 296996 294964
rect 215812 294924 215818 294936
rect 296990 294924 296996 294936
rect 297048 294924 297054 294976
rect 214374 294856 214380 294908
rect 214432 294896 214438 294908
rect 297082 294896 297088 294908
rect 214432 294868 297088 294896
rect 214432 294856 214438 294868
rect 297082 294856 297088 294868
rect 297140 294856 297146 294908
rect 213270 294788 213276 294840
rect 213328 294828 213334 294840
rect 296898 294828 296904 294840
rect 213328 294800 296904 294828
rect 213328 294788 213334 294800
rect 296898 294788 296904 294800
rect 296956 294788 296962 294840
rect 168374 294720 168380 294772
rect 168432 294760 168438 294772
rect 278774 294760 278780 294772
rect 168432 294732 278780 294760
rect 168432 294720 168438 294732
rect 278774 294720 278780 294732
rect 278832 294720 278838 294772
rect 315022 294720 315028 294772
rect 315080 294760 315086 294772
rect 387058 294760 387064 294772
rect 315080 294732 387064 294760
rect 315080 294720 315086 294732
rect 387058 294720 387064 294732
rect 387116 294720 387122 294772
rect 135254 294652 135260 294704
rect 135312 294692 135318 294704
rect 274726 294692 274732 294704
rect 135312 294664 274732 294692
rect 135312 294652 135318 294664
rect 274726 294652 274732 294664
rect 274784 294652 274790 294704
rect 326062 294652 326068 294704
rect 326120 294692 326126 294704
rect 457438 294692 457444 294704
rect 326120 294664 457444 294692
rect 326120 294652 326126 294664
rect 457438 294652 457444 294664
rect 457496 294652 457502 294704
rect 43438 294584 43444 294636
rect 43496 294624 43502 294636
rect 258626 294624 258632 294636
rect 43496 294596 258632 294624
rect 43496 294584 43502 294596
rect 258626 294584 258632 294596
rect 258684 294584 258690 294636
rect 337194 294584 337200 294636
rect 337252 294624 337258 294636
rect 525794 294624 525800 294636
rect 337252 294596 525800 294624
rect 337252 294584 337258 294596
rect 525794 294584 525800 294596
rect 525852 294584 525858 294636
rect 202874 293360 202880 293412
rect 202932 293400 202938 293412
rect 284662 293400 284668 293412
rect 202932 293372 284668 293400
rect 202932 293360 202938 293372
rect 284662 293360 284668 293372
rect 284720 293360 284726 293412
rect 329098 293360 329104 293412
rect 329156 293400 329162 293412
rect 467098 293400 467104 293412
rect 329156 293372 467104 293400
rect 329156 293360 329162 293372
rect 467098 293360 467104 293372
rect 467156 293360 467162 293412
rect 58618 293292 58624 293344
rect 58676 293332 58682 293344
rect 260834 293332 260840 293344
rect 58676 293304 260840 293332
rect 58676 293292 58682 293304
rect 260834 293292 260840 293304
rect 260892 293292 260898 293344
rect 335722 293292 335728 293344
rect 335780 293332 335786 293344
rect 509878 293332 509884 293344
rect 335780 293304 509884 293332
rect 335780 293292 335786 293304
rect 509878 293292 509884 293304
rect 509936 293292 509942 293344
rect 13078 293224 13084 293276
rect 13136 293264 13142 293276
rect 254302 293264 254308 293276
rect 13136 293236 254308 293264
rect 13136 293224 13142 293236
rect 254302 293224 254308 293236
rect 254360 293224 254366 293276
rect 338574 293224 338580 293276
rect 338632 293264 338638 293276
rect 527818 293264 527824 293276
rect 338632 293236 527824 293264
rect 338632 293224 338638 293236
rect 527818 293224 527824 293236
rect 527876 293224 527882 293276
rect 161474 292000 161480 292052
rect 161532 292040 161538 292052
rect 279142 292040 279148 292052
rect 161532 292012 279148 292040
rect 161532 292000 161538 292012
rect 279142 292000 279148 292012
rect 279200 292000 279206 292052
rect 128354 291932 128360 291984
rect 128412 291972 128418 291984
rect 271138 291972 271144 291984
rect 128412 291944 271144 291972
rect 128412 291932 128418 291944
rect 271138 291932 271144 291944
rect 271196 291932 271202 291984
rect 71038 291864 71044 291916
rect 71096 291904 71102 291916
rect 263594 291904 263600 291916
rect 71096 291876 263600 291904
rect 71096 291864 71102 291876
rect 263594 291864 263600 291876
rect 263652 291864 263658 291916
rect 317782 291864 317788 291916
rect 317840 291904 317846 291916
rect 405734 291904 405740 291916
rect 317840 291876 405740 291904
rect 317840 291864 317846 291876
rect 405734 291864 405740 291876
rect 405792 291864 405798 291916
rect 27614 291796 27620 291848
rect 27672 291836 27678 291848
rect 257430 291836 257436 291848
rect 27672 291808 257436 291836
rect 27672 291796 27678 291808
rect 257430 291796 257436 291808
rect 257488 291796 257494 291848
rect 338482 291796 338488 291848
rect 338540 291836 338546 291848
rect 534718 291836 534724 291848
rect 338540 291808 534724 291836
rect 338540 291796 338546 291808
rect 534718 291796 534724 291808
rect 534776 291796 534782 291848
rect 187694 290640 187700 290692
rect 187752 290680 187758 290692
rect 283282 290680 283288 290692
rect 187752 290652 283288 290680
rect 187752 290640 187758 290652
rect 283282 290640 283288 290652
rect 283340 290640 283346 290692
rect 317690 290640 317696 290692
rect 317748 290680 317754 290692
rect 408494 290680 408500 290692
rect 317748 290652 408500 290680
rect 317748 290640 317754 290652
rect 408494 290640 408500 290652
rect 408552 290640 408558 290692
rect 143534 290572 143540 290624
rect 143592 290612 143598 290624
rect 274634 290612 274640 290624
rect 143592 290584 274640 290612
rect 143592 290572 143598 290584
rect 274634 290572 274640 290584
rect 274692 290572 274698 290624
rect 320634 290572 320640 290624
rect 320692 290612 320698 290624
rect 418154 290612 418160 290624
rect 320692 290584 418160 290612
rect 320692 290572 320698 290584
rect 418154 290572 418160 290584
rect 418212 290572 418218 290624
rect 57238 290504 57244 290556
rect 57296 290544 57302 290556
rect 261294 290544 261300 290556
rect 57296 290516 261300 290544
rect 57296 290504 57302 290516
rect 261294 290504 261300 290516
rect 261352 290504 261358 290556
rect 341334 290504 341340 290556
rect 341392 290544 341398 290556
rect 542998 290544 543004 290556
rect 341392 290516 543004 290544
rect 341392 290504 341398 290516
rect 542998 290504 543004 290516
rect 543056 290504 543062 290556
rect 8294 290436 8300 290488
rect 8352 290476 8358 290488
rect 254210 290476 254216 290488
rect 8352 290448 254216 290476
rect 8352 290436 8358 290448
rect 254210 290436 254216 290448
rect 254268 290436 254274 290488
rect 341242 290436 341248 290488
rect 341300 290476 341306 290488
rect 549898 290476 549904 290488
rect 341300 290448 549904 290476
rect 341300 290436 341306 290448
rect 549898 290436 549904 290448
rect 549956 290436 549962 290488
rect 205634 289280 205640 289332
rect 205692 289320 205698 289332
rect 286042 289320 286048 289332
rect 205692 289292 286048 289320
rect 205692 289280 205698 289292
rect 286042 289280 286048 289292
rect 286100 289280 286106 289332
rect 132494 289212 132500 289264
rect 132552 289252 132558 289264
rect 273622 289252 273628 289264
rect 132552 289224 273628 289252
rect 132552 289212 132558 289224
rect 273622 289212 273628 289224
rect 273680 289212 273686 289264
rect 321922 289212 321928 289264
rect 321980 289252 321986 289264
rect 430574 289252 430580 289264
rect 321980 289224 430580 289252
rect 321980 289212 321986 289224
rect 430574 289212 430580 289224
rect 430632 289212 430638 289264
rect 103514 289144 103520 289196
rect 103572 289184 103578 289196
rect 269758 289184 269764 289196
rect 103572 289156 269764 289184
rect 103572 289144 103578 289156
rect 269758 289144 269764 289156
rect 269816 289144 269822 289196
rect 331490 289144 331496 289196
rect 331548 289184 331554 289196
rect 490006 289184 490012 289196
rect 331548 289156 490012 289184
rect 331548 289144 331554 289156
rect 490006 289144 490012 289156
rect 490064 289144 490070 289196
rect 9674 289076 9680 289128
rect 9732 289116 9738 289128
rect 254118 289116 254124 289128
rect 9732 289088 254124 289116
rect 9732 289076 9738 289088
rect 254118 289076 254124 289088
rect 254176 289076 254182 289128
rect 341150 289076 341156 289128
rect 341208 289116 341214 289128
rect 552658 289116 552664 289128
rect 341208 289088 552664 289116
rect 341208 289076 341214 289088
rect 552658 289076 552664 289088
rect 552716 289076 552722 289128
rect 313550 287920 313556 287972
rect 313608 287960 313614 287972
rect 382274 287960 382280 287972
rect 313608 287932 382280 287960
rect 313608 287920 313614 287932
rect 382274 287920 382280 287932
rect 382332 287920 382338 287972
rect 181438 287852 181444 287904
rect 181496 287892 181502 287904
rect 281902 287892 281908 287904
rect 181496 287864 281908 287892
rect 181496 287852 181502 287864
rect 281902 287852 281908 287864
rect 281960 287852 281966 287904
rect 327534 287852 327540 287904
rect 327592 287892 327598 287904
rect 460198 287892 460204 287904
rect 327592 287864 460204 287892
rect 327592 287852 327598 287864
rect 460198 287852 460204 287864
rect 460256 287852 460262 287904
rect 217686 287784 217692 287836
rect 217744 287824 217750 287836
rect 351178 287824 351184 287836
rect 217744 287796 351184 287824
rect 217744 287784 217750 287796
rect 351178 287784 351184 287796
rect 351236 287784 351242 287836
rect 139394 287716 139400 287768
rect 139452 287756 139458 287768
rect 275094 287756 275100 287768
rect 139452 287728 275100 287756
rect 139452 287716 139458 287728
rect 275094 287716 275100 287728
rect 275152 287716 275158 287768
rect 337102 287716 337108 287768
rect 337160 287756 337166 287768
rect 518158 287756 518164 287768
rect 337160 287728 518164 287756
rect 337160 287716 337166 287728
rect 518158 287716 518164 287728
rect 518216 287716 518222 287768
rect 22094 287648 22100 287700
rect 22152 287688 22158 287700
rect 255682 287688 255688 287700
rect 22152 287660 255688 287688
rect 22152 287648 22158 287660
rect 255682 287648 255688 287660
rect 255740 287648 255746 287700
rect 342622 287648 342628 287700
rect 342680 287688 342686 287700
rect 561674 287688 561680 287700
rect 342680 287660 561680 287688
rect 342680 287648 342686 287660
rect 561674 287648 561680 287660
rect 561732 287648 561738 287700
rect 203518 286560 203524 286612
rect 203576 286600 203582 286612
rect 283190 286600 283196 286612
rect 203576 286572 283196 286600
rect 203576 286560 203582 286572
rect 283190 286560 283196 286572
rect 283248 286560 283254 286612
rect 146294 286492 146300 286544
rect 146352 286532 146358 286544
rect 276566 286532 276572 286544
rect 146352 286504 276572 286532
rect 146352 286492 146358 286504
rect 276566 286492 276572 286504
rect 276624 286492 276630 286544
rect 46934 286424 46940 286476
rect 46992 286464 46998 286476
rect 259822 286464 259828 286476
rect 46992 286436 259828 286464
rect 46992 286424 46998 286436
rect 259822 286424 259828 286436
rect 259880 286424 259886 286476
rect 325970 286424 325976 286476
rect 326028 286464 326034 286476
rect 454678 286464 454684 286476
rect 326028 286436 454684 286464
rect 326028 286424 326034 286436
rect 454678 286424 454684 286436
rect 454736 286424 454742 286476
rect 40034 286356 40040 286408
rect 40092 286396 40098 286408
rect 258442 286396 258448 286408
rect 40092 286368 258448 286396
rect 40092 286356 40098 286368
rect 258442 286356 258448 286368
rect 258500 286356 258506 286408
rect 327442 286356 327448 286408
rect 327500 286396 327506 286408
rect 458818 286396 458824 286408
rect 327500 286368 458824 286396
rect 327500 286356 327506 286368
rect 458818 286356 458824 286368
rect 458876 286356 458882 286408
rect 18598 286288 18604 286340
rect 18656 286328 18662 286340
rect 252922 286328 252928 286340
rect 18656 286300 252928 286328
rect 18656 286288 18662 286300
rect 252922 286288 252928 286300
rect 252980 286288 252986 286340
rect 344002 286288 344008 286340
rect 344060 286328 344066 286340
rect 566458 286328 566464 286340
rect 344060 286300 566464 286328
rect 344060 286288 344066 286300
rect 566458 286288 566464 286300
rect 566516 286288 566522 286340
rect 150434 285132 150440 285184
rect 150492 285172 150498 285184
rect 276474 285172 276480 285184
rect 150492 285144 276480 285172
rect 150492 285132 150498 285144
rect 276474 285132 276480 285144
rect 276532 285132 276538 285184
rect 81434 285064 81440 285116
rect 81492 285104 81498 285116
rect 265526 285104 265532 285116
rect 81492 285076 265532 285104
rect 81492 285064 81498 285076
rect 265526 285064 265532 285076
rect 265584 285064 265590 285116
rect 311986 285064 311992 285116
rect 312044 285104 312050 285116
rect 371878 285104 371884 285116
rect 312044 285076 371884 285104
rect 312044 285064 312050 285076
rect 371878 285064 371884 285076
rect 371936 285064 371942 285116
rect 26234 284996 26240 285048
rect 26292 285036 26298 285048
rect 257062 285036 257068 285048
rect 26292 285008 257068 285036
rect 26292 284996 26298 285008
rect 257062 284996 257068 285008
rect 257120 284996 257126 285048
rect 329006 284996 329012 285048
rect 329064 285036 329070 285048
rect 471238 285036 471244 285048
rect 329064 285008 471244 285036
rect 329064 284996 329070 285008
rect 471238 284996 471244 285008
rect 471296 284996 471302 285048
rect 2774 284928 2780 284980
rect 2832 284968 2838 284980
rect 252830 284968 252836 284980
rect 2832 284940 252836 284968
rect 2832 284928 2838 284940
rect 252830 284928 252836 284940
rect 252888 284928 252894 284980
rect 345474 284928 345480 284980
rect 345532 284968 345538 284980
rect 575474 284968 575480 284980
rect 345532 284940 575480 284968
rect 345532 284928 345538 284940
rect 575474 284928 575480 284940
rect 575532 284928 575538 284980
rect 211154 283772 211160 283824
rect 211212 283812 211218 283824
rect 285858 283812 285864 283824
rect 211212 283784 285864 283812
rect 211212 283772 211218 283784
rect 285858 283772 285864 283784
rect 285916 283772 285922 283824
rect 314930 283772 314936 283824
rect 314988 283812 314994 283824
rect 390554 283812 390560 283824
rect 314988 283784 390560 283812
rect 314988 283772 314994 283784
rect 390554 283772 390560 283784
rect 390612 283772 390618 283824
rect 153194 283704 153200 283756
rect 153252 283744 153258 283756
rect 277854 283744 277860 283756
rect 153252 283716 277860 283744
rect 153252 283704 153258 283716
rect 277854 283704 277860 283716
rect 277912 283704 277918 283756
rect 324866 283704 324872 283756
rect 324924 283744 324930 283756
rect 442258 283744 442264 283756
rect 324924 283716 442264 283744
rect 324924 283704 324930 283716
rect 442258 283704 442264 283716
rect 442316 283704 442322 283756
rect 138014 283636 138020 283688
rect 138072 283676 138078 283688
rect 275002 283676 275008 283688
rect 138072 283648 275008 283676
rect 138072 283636 138078 283648
rect 275002 283636 275008 283648
rect 275060 283636 275066 283688
rect 337010 283636 337016 283688
rect 337068 283676 337074 283688
rect 522298 283676 522304 283688
rect 337068 283648 522304 283676
rect 337068 283636 337074 283648
rect 522298 283636 522304 283648
rect 522356 283636 522362 283688
rect 16574 283568 16580 283620
rect 16632 283608 16638 283620
rect 255590 283608 255596 283620
rect 16632 283580 255596 283608
rect 16632 283568 16638 283580
rect 255590 283568 255596 283580
rect 255648 283568 255654 283620
rect 338390 283568 338396 283620
rect 338448 283608 338454 283620
rect 531314 283608 531320 283620
rect 338448 283580 531320 283608
rect 338448 283568 338454 283580
rect 531314 283568 531320 283580
rect 531372 283568 531378 283620
rect 157334 282344 157340 282396
rect 157392 282384 157398 282396
rect 277762 282384 277768 282396
rect 157392 282356 277768 282384
rect 157392 282344 157398 282356
rect 277762 282344 277768 282356
rect 277820 282344 277826 282396
rect 313458 282344 313464 282396
rect 313516 282384 313522 282396
rect 374638 282384 374644 282396
rect 313516 282356 374644 282384
rect 313516 282344 313522 282356
rect 374638 282344 374644 282356
rect 374696 282344 374702 282396
rect 131114 282276 131120 282328
rect 131172 282316 131178 282328
rect 273530 282316 273536 282328
rect 131172 282288 273536 282316
rect 131172 282276 131178 282288
rect 273530 282276 273536 282288
rect 273588 282276 273594 282328
rect 319162 282276 319168 282328
rect 319220 282316 319226 282328
rect 414658 282316 414664 282328
rect 319220 282288 414664 282316
rect 319220 282276 319226 282288
rect 414658 282276 414664 282288
rect 414716 282276 414722 282328
rect 114554 282208 114560 282260
rect 114612 282248 114618 282260
rect 270954 282248 270960 282260
rect 114612 282220 270960 282248
rect 114612 282208 114618 282220
rect 270954 282208 270960 282220
rect 271012 282208 271018 282260
rect 327350 282208 327356 282260
rect 327408 282248 327414 282260
rect 464338 282248 464344 282260
rect 327408 282220 464344 282248
rect 327408 282208 327414 282220
rect 464338 282208 464344 282220
rect 464396 282208 464402 282260
rect 44174 282140 44180 282192
rect 44232 282180 44238 282192
rect 259730 282180 259736 282192
rect 44232 282152 259736 282180
rect 44232 282140 44238 282152
rect 259730 282140 259736 282152
rect 259788 282140 259794 282192
rect 342530 282140 342536 282192
rect 342588 282180 342594 282192
rect 556246 282180 556252 282192
rect 342588 282152 556252 282180
rect 342588 282140 342594 282152
rect 556246 282140 556252 282152
rect 556304 282140 556310 282192
rect 198734 280984 198740 281036
rect 198792 281024 198798 281036
rect 284570 281024 284576 281036
rect 198792 280996 284576 281024
rect 198792 280984 198798 280996
rect 284570 280984 284576 280996
rect 284628 280984 284634 281036
rect 126974 280916 126980 280968
rect 127032 280956 127038 280968
rect 272242 280956 272248 280968
rect 127032 280928 272248 280956
rect 127032 280916 127038 280928
rect 272242 280916 272248 280928
rect 272300 280916 272306 280968
rect 107654 280848 107660 280900
rect 107712 280888 107718 280900
rect 269574 280888 269580 280900
rect 107712 280860 269580 280888
rect 107712 280848 107718 280860
rect 269574 280848 269580 280860
rect 269632 280848 269638 280900
rect 320542 280848 320548 280900
rect 320600 280888 320606 280900
rect 417418 280888 417424 280900
rect 320600 280860 417424 280888
rect 320600 280848 320606 280860
rect 417418 280848 417424 280860
rect 417476 280848 417482 280900
rect 34514 280780 34520 280832
rect 34572 280820 34578 280832
rect 258350 280820 258356 280832
rect 34572 280792 258356 280820
rect 34572 280780 34578 280792
rect 258350 280780 258356 280792
rect 258408 280780 258414 280832
rect 345382 280780 345388 280832
rect 345440 280820 345446 280832
rect 571978 280820 571984 280832
rect 345440 280792 571984 280820
rect 345440 280780 345446 280792
rect 571978 280780 571984 280792
rect 572036 280780 572042 280832
rect 165614 279624 165620 279676
rect 165672 279664 165678 279676
rect 279050 279664 279056 279676
rect 165672 279636 279056 279664
rect 165672 279624 165678 279636
rect 279050 279624 279056 279636
rect 279108 279624 279114 279676
rect 97994 279556 98000 279608
rect 98052 279596 98058 279608
rect 268194 279596 268200 279608
rect 98052 279568 268200 279596
rect 98052 279556 98058 279568
rect 268194 279556 268200 279568
rect 268252 279556 268258 279608
rect 317598 279556 317604 279608
rect 317656 279596 317662 279608
rect 407114 279596 407120 279608
rect 317656 279568 407120 279596
rect 317656 279556 317662 279568
rect 407114 279556 407120 279568
rect 407172 279556 407178 279608
rect 71774 279488 71780 279540
rect 71832 279528 71838 279540
rect 264146 279528 264152 279540
rect 71832 279500 264152 279528
rect 71832 279488 71838 279500
rect 264146 279488 264152 279500
rect 264204 279488 264210 279540
rect 320450 279488 320456 279540
rect 320508 279528 320514 279540
rect 423674 279528 423680 279540
rect 320508 279500 423680 279528
rect 320508 279488 320514 279500
rect 423674 279488 423680 279500
rect 423732 279488 423738 279540
rect 38654 279420 38660 279472
rect 38712 279460 38718 279472
rect 257338 279460 257344 279472
rect 38712 279432 257344 279460
rect 38712 279420 38718 279432
rect 257338 279420 257344 279432
rect 257396 279420 257402 279472
rect 332962 279420 332968 279472
rect 333020 279460 333026 279472
rect 493318 279460 493324 279472
rect 333020 279432 493324 279460
rect 333020 279420 333026 279432
rect 493318 279420 493324 279432
rect 493376 279420 493382 279472
rect 188338 278264 188344 278316
rect 188396 278304 188402 278316
rect 281810 278304 281816 278316
rect 188396 278276 281816 278304
rect 188396 278264 188402 278276
rect 281810 278264 281816 278276
rect 281868 278264 281874 278316
rect 147674 278196 147680 278248
rect 147732 278236 147738 278248
rect 276382 278236 276388 278248
rect 147732 278208 276388 278236
rect 147732 278196 147738 278208
rect 276382 278196 276388 278208
rect 276440 278196 276446 278248
rect 102134 278128 102140 278180
rect 102192 278168 102198 278180
rect 269482 278168 269488 278180
rect 102192 278140 269488 278168
rect 102192 278128 102198 278140
rect 269482 278128 269488 278140
rect 269540 278128 269546 278180
rect 319070 278128 319076 278180
rect 319128 278168 319134 278180
rect 409874 278168 409880 278180
rect 319128 278140 409880 278168
rect 319128 278128 319134 278140
rect 409874 278128 409880 278140
rect 409932 278128 409938 278180
rect 78674 278060 78680 278112
rect 78732 278100 78738 278112
rect 265434 278100 265440 278112
rect 78732 278072 265440 278100
rect 78732 278060 78738 278072
rect 265434 278060 265440 278072
rect 265492 278060 265498 278112
rect 321830 278060 321836 278112
rect 321888 278100 321894 278112
rect 428458 278100 428464 278112
rect 321888 278072 428464 278100
rect 321888 278060 321894 278072
rect 428458 278060 428464 278072
rect 428516 278060 428522 278112
rect 35894 277992 35900 278044
rect 35952 278032 35958 278044
rect 258258 278032 258264 278044
rect 35952 278004 258264 278032
rect 35952 277992 35958 278004
rect 258258 277992 258264 278004
rect 258316 277992 258322 278044
rect 341058 277992 341064 278044
rect 341116 278032 341122 278044
rect 553394 278032 553400 278044
rect 341116 278004 553400 278032
rect 341116 277992 341122 278004
rect 553394 277992 553400 278004
rect 553452 277992 553458 278044
rect 196618 276836 196624 276888
rect 196676 276876 196682 276888
rect 281718 276876 281724 276888
rect 196676 276848 281724 276876
rect 196676 276836 196682 276848
rect 281718 276836 281724 276848
rect 281776 276836 281782 276888
rect 136634 276768 136640 276820
rect 136692 276808 136698 276820
rect 274910 276808 274916 276820
rect 136692 276780 274916 276808
rect 136692 276768 136698 276780
rect 274910 276768 274916 276780
rect 274968 276768 274974 276820
rect 325878 276768 325884 276820
rect 325936 276808 325942 276820
rect 445018 276808 445024 276820
rect 325936 276780 445024 276808
rect 325936 276768 325942 276780
rect 445018 276768 445024 276780
rect 445076 276768 445082 276820
rect 111794 276700 111800 276752
rect 111852 276740 111858 276752
rect 270862 276740 270868 276752
rect 111852 276712 270868 276740
rect 111852 276700 111858 276712
rect 270862 276700 270868 276712
rect 270920 276700 270926 276752
rect 324774 276700 324780 276752
rect 324832 276740 324838 276752
rect 448514 276740 448520 276752
rect 324832 276712 448520 276740
rect 324832 276700 324838 276712
rect 448514 276700 448520 276712
rect 448572 276700 448578 276752
rect 27706 276632 27712 276684
rect 27764 276672 27770 276684
rect 256970 276672 256976 276684
rect 27764 276644 256976 276672
rect 27764 276632 27770 276644
rect 256970 276632 256976 276644
rect 257028 276632 257034 276684
rect 335630 276632 335636 276684
rect 335688 276672 335694 276684
rect 511258 276672 511264 276684
rect 335688 276644 511264 276672
rect 335688 276632 335694 276644
rect 511258 276632 511264 276644
rect 511316 276632 511322 276684
rect 193306 275544 193312 275596
rect 193364 275584 193370 275596
rect 283098 275584 283104 275596
rect 193364 275556 283104 275584
rect 193364 275544 193370 275556
rect 283098 275544 283104 275556
rect 283156 275544 283162 275596
rect 127066 275476 127072 275528
rect 127124 275516 127130 275528
rect 273438 275516 273444 275528
rect 127124 275488 273444 275516
rect 127124 275476 127130 275488
rect 273438 275476 273444 275488
rect 273496 275476 273502 275528
rect 317506 275476 317512 275528
rect 317564 275516 317570 275528
rect 404354 275516 404360 275528
rect 317564 275488 404360 275516
rect 317564 275476 317570 275488
rect 404354 275476 404360 275488
rect 404412 275476 404418 275528
rect 115934 275408 115940 275460
rect 115992 275448 115998 275460
rect 270770 275448 270776 275460
rect 115992 275420 270776 275448
rect 115992 275408 115998 275420
rect 270770 275408 270776 275420
rect 270828 275408 270834 275460
rect 324682 275408 324688 275460
rect 324740 275448 324746 275460
rect 448606 275448 448612 275460
rect 324740 275420 448612 275448
rect 324740 275408 324746 275420
rect 448606 275408 448612 275420
rect 448664 275408 448670 275460
rect 96614 275340 96620 275392
rect 96672 275380 96678 275392
rect 268102 275380 268108 275392
rect 96672 275352 268108 275380
rect 96672 275340 96678 275352
rect 268102 275340 268108 275352
rect 268160 275340 268166 275392
rect 328914 275340 328920 275392
rect 328972 275380 328978 275392
rect 468478 275380 468484 275392
rect 328972 275352 468484 275380
rect 328972 275340 328978 275352
rect 468478 275340 468484 275352
rect 468536 275340 468542 275392
rect 42794 275272 42800 275324
rect 42852 275312 42858 275324
rect 250530 275312 250536 275324
rect 42852 275284 250536 275312
rect 42852 275272 42858 275284
rect 250530 275272 250536 275284
rect 250588 275272 250594 275324
rect 336918 275272 336924 275324
rect 336976 275312 336982 275324
rect 525058 275312 525064 275324
rect 336976 275284 525064 275312
rect 336976 275272 336982 275284
rect 525058 275272 525064 275284
rect 525116 275272 525122 275324
rect 197354 274184 197360 274236
rect 197412 274224 197418 274236
rect 284478 274224 284484 274236
rect 197412 274196 284484 274224
rect 197412 274184 197418 274196
rect 284478 274184 284484 274196
rect 284536 274184 284542 274236
rect 162854 274116 162860 274168
rect 162912 274156 162918 274168
rect 278958 274156 278964 274168
rect 162912 274128 278964 274156
rect 162912 274116 162918 274128
rect 278958 274116 278964 274128
rect 279016 274116 279022 274168
rect 324590 274116 324596 274168
rect 324648 274156 324654 274168
rect 446398 274156 446404 274168
rect 324648 274128 446404 274156
rect 324648 274116 324654 274128
rect 446398 274116 446404 274128
rect 446456 274116 446462 274168
rect 113174 274048 113180 274100
rect 113232 274088 113238 274100
rect 270678 274088 270684 274100
rect 113232 274060 270684 274088
rect 113232 274048 113238 274060
rect 270678 274048 270684 274060
rect 270736 274048 270742 274100
rect 327258 274048 327264 274100
rect 327316 274088 327322 274100
rect 460934 274088 460940 274100
rect 327316 274060 460940 274088
rect 327316 274048 327322 274060
rect 460934 274048 460940 274060
rect 460992 274048 460998 274100
rect 93854 273980 93860 274032
rect 93912 274020 93918 274032
rect 268010 274020 268016 274032
rect 93912 273992 268016 274020
rect 93912 273980 93918 273992
rect 268010 273980 268016 273992
rect 268068 273980 268074 274032
rect 325786 273980 325792 274032
rect 325844 274020 325850 274032
rect 459554 274020 459560 274032
rect 325844 273992 459560 274020
rect 325844 273980 325850 273992
rect 459554 273980 459560 273992
rect 459612 273980 459618 274032
rect 14458 273912 14464 273964
rect 14516 273952 14522 273964
rect 254026 273952 254032 273964
rect 14516 273924 254032 273952
rect 14516 273912 14522 273924
rect 254026 273912 254032 273924
rect 254084 273912 254090 273964
rect 338298 273912 338304 273964
rect 338356 273952 338362 273964
rect 531406 273952 531412 273964
rect 338356 273924 531412 273952
rect 338356 273912 338362 273924
rect 531406 273912 531412 273924
rect 531464 273912 531470 273964
rect 201494 272756 201500 272808
rect 201552 272796 201558 272808
rect 284386 272796 284392 272808
rect 201552 272768 284392 272796
rect 201552 272756 201558 272768
rect 284386 272756 284392 272768
rect 284444 272756 284450 272808
rect 180794 272688 180800 272740
rect 180852 272728 180858 272740
rect 281626 272728 281632 272740
rect 180852 272700 281632 272728
rect 180852 272688 180858 272700
rect 281626 272688 281632 272700
rect 281684 272688 281690 272740
rect 99374 272620 99380 272672
rect 99432 272660 99438 272672
rect 260098 272660 260104 272672
rect 99432 272632 260104 272660
rect 99432 272620 99438 272632
rect 260098 272620 260104 272632
rect 260156 272620 260162 272672
rect 84194 272552 84200 272604
rect 84252 272592 84258 272604
rect 265342 272592 265348 272604
rect 84252 272564 265348 272592
rect 84252 272552 84258 272564
rect 265342 272552 265348 272564
rect 265400 272552 265406 272604
rect 53834 272484 53840 272536
rect 53892 272524 53898 272536
rect 261202 272524 261208 272536
rect 53892 272496 261208 272524
rect 53892 272484 53898 272496
rect 261202 272484 261208 272496
rect 261260 272484 261266 272536
rect 328822 272484 328828 272536
rect 328880 272524 328886 272536
rect 475378 272524 475384 272536
rect 328880 272496 475384 272524
rect 328880 272484 328886 272496
rect 475378 272484 475384 272496
rect 475436 272484 475442 272536
rect 211798 271328 211804 271380
rect 211856 271368 211862 271380
rect 286226 271368 286232 271380
rect 211856 271340 286232 271368
rect 211856 271328 211862 271340
rect 286226 271328 286232 271340
rect 286284 271328 286290 271380
rect 166994 271260 167000 271312
rect 167052 271300 167058 271312
rect 278866 271300 278872 271312
rect 167052 271272 278872 271300
rect 167052 271260 167058 271272
rect 278866 271260 278872 271272
rect 278924 271260 278930 271312
rect 102226 271192 102232 271244
rect 102284 271232 102290 271244
rect 269390 271232 269396 271244
rect 102284 271204 269396 271232
rect 102284 271192 102290 271204
rect 269390 271192 269396 271204
rect 269448 271192 269454 271244
rect 314838 271192 314844 271244
rect 314896 271232 314902 271244
rect 386414 271232 386420 271244
rect 314896 271204 386420 271232
rect 314896 271192 314902 271204
rect 386414 271192 386420 271204
rect 386472 271192 386478 271244
rect 57974 271124 57980 271176
rect 58032 271164 58038 271176
rect 261110 271164 261116 271176
rect 58032 271136 261116 271164
rect 58032 271124 58038 271136
rect 261110 271124 261116 271136
rect 261168 271124 261174 271176
rect 335538 271124 335544 271176
rect 335596 271164 335602 271176
rect 517514 271164 517520 271176
rect 335596 271136 517520 271164
rect 335596 271124 335602 271136
rect 517514 271124 517520 271136
rect 517572 271124 517578 271176
rect 151814 269968 151820 270020
rect 151872 270008 151878 270020
rect 276290 270008 276296 270020
rect 151872 269980 276296 270008
rect 151872 269968 151878 269980
rect 276290 269968 276296 269980
rect 276348 269968 276354 270020
rect 318058 269968 318064 270020
rect 318116 270008 318122 270020
rect 400214 270008 400220 270020
rect 318116 269980 400220 270008
rect 318116 269968 318122 269980
rect 400214 269968 400220 269980
rect 400272 269968 400278 270020
rect 110414 269900 110420 269952
rect 110472 269940 110478 269952
rect 269298 269940 269304 269952
rect 110472 269912 269304 269940
rect 110472 269900 110478 269912
rect 269298 269900 269304 269912
rect 269356 269900 269362 269952
rect 320358 269900 320364 269952
rect 320416 269940 320422 269952
rect 420914 269940 420920 269952
rect 320416 269912 420920 269940
rect 320416 269900 320422 269912
rect 420914 269900 420920 269912
rect 420972 269900 420978 269952
rect 93946 269832 93952 269884
rect 94004 269872 94010 269884
rect 267918 269872 267924 269884
rect 94004 269844 267924 269872
rect 94004 269832 94010 269844
rect 267918 269832 267924 269844
rect 267976 269832 267982 269884
rect 331398 269832 331404 269884
rect 331456 269872 331462 269884
rect 486418 269872 486424 269884
rect 331456 269844 486424 269872
rect 331456 269832 331462 269844
rect 486418 269832 486424 269844
rect 486476 269832 486482 269884
rect 75914 269764 75920 269816
rect 75972 269804 75978 269816
rect 264054 269804 264060 269816
rect 75972 269776 264060 269804
rect 75972 269764 75978 269776
rect 264054 269764 264060 269776
rect 264112 269764 264118 269816
rect 340966 269764 340972 269816
rect 341024 269804 341030 269816
rect 552014 269804 552020 269816
rect 341024 269776 552020 269804
rect 341024 269764 341030 269776
rect 552014 269764 552020 269776
rect 552072 269764 552078 269816
rect 151906 268472 151912 268524
rect 151964 268512 151970 268524
rect 276198 268512 276204 268524
rect 151964 268484 276204 268512
rect 151964 268472 151970 268484
rect 276198 268472 276204 268484
rect 276256 268472 276262 268524
rect 143626 268404 143632 268456
rect 143684 268444 143690 268456
rect 274818 268444 274824 268456
rect 143684 268416 274824 268444
rect 143684 268404 143690 268416
rect 274818 268404 274824 268416
rect 274876 268404 274882 268456
rect 328638 268404 328644 268456
rect 328696 268444 328702 268456
rect 473446 268444 473452 268456
rect 328696 268416 473452 268444
rect 328696 268404 328702 268416
rect 473446 268404 473452 268416
rect 473504 268404 473510 268456
rect 77294 268336 77300 268388
rect 77352 268376 77358 268388
rect 265250 268376 265256 268388
rect 77352 268348 265256 268376
rect 77352 268336 77358 268348
rect 265250 268336 265256 268348
rect 265308 268336 265314 268388
rect 328730 268336 328736 268388
rect 328788 268376 328794 268388
rect 474734 268376 474740 268388
rect 328788 268348 474740 268376
rect 328788 268336 328794 268348
rect 474734 268336 474740 268348
rect 474792 268336 474798 268388
rect 2958 267656 2964 267708
rect 3016 267696 3022 267708
rect 225598 267696 225604 267708
rect 3016 267668 225604 267696
rect 3016 267656 3022 267668
rect 225598 267656 225604 267668
rect 225656 267656 225662 267708
rect 317414 267248 317420 267300
rect 317472 267288 317478 267300
rect 407206 267288 407212 267300
rect 317472 267260 407212 267288
rect 317472 267248 317478 267260
rect 407206 267248 407212 267260
rect 407264 267248 407270 267300
rect 217318 267180 217324 267232
rect 217376 267220 217382 267232
rect 351086 267220 351092 267232
rect 217376 267192 351092 267220
rect 217376 267180 217382 267192
rect 351086 267180 351092 267192
rect 351144 267180 351150 267232
rect 332870 267112 332876 267164
rect 332928 267152 332934 267164
rect 495434 267152 495440 267164
rect 332928 267124 495440 267152
rect 332928 267112 332934 267124
rect 495434 267112 495440 267124
rect 495492 267112 495498 267164
rect 340874 267044 340880 267096
rect 340932 267084 340938 267096
rect 549254 267084 549260 267096
rect 340932 267056 549260 267084
rect 340932 267044 340938 267056
rect 549254 267044 549260 267056
rect 549312 267044 549318 267096
rect 70394 266976 70400 267028
rect 70452 267016 70458 267028
rect 263962 267016 263968 267028
rect 70452 266988 263968 267016
rect 70452 266976 70458 266988
rect 263962 266976 263968 266988
rect 264020 266976 264026 267028
rect 343910 266976 343916 267028
rect 343968 267016 343974 267028
rect 565814 267016 565820 267028
rect 343968 266988 565820 267016
rect 343968 266976 343974 266988
rect 565814 266976 565820 266988
rect 565872 266976 565878 267028
rect 191834 265888 191840 265940
rect 191892 265928 191898 265940
rect 283466 265928 283472 265940
rect 191892 265900 283472 265928
rect 191892 265888 191898 265900
rect 283466 265888 283472 265900
rect 283524 265888 283530 265940
rect 133874 265820 133880 265872
rect 133932 265860 133938 265872
rect 273346 265860 273352 265872
rect 133932 265832 273352 265860
rect 133932 265820 133938 265832
rect 273346 265820 273352 265832
rect 273404 265820 273410 265872
rect 313366 265820 313372 265872
rect 313424 265860 313430 265872
rect 382366 265860 382372 265872
rect 313424 265832 382372 265860
rect 313424 265820 313430 265832
rect 382366 265820 382372 265832
rect 382424 265820 382430 265872
rect 121454 265752 121460 265804
rect 121512 265792 121518 265804
rect 272150 265792 272156 265804
rect 121512 265764 272156 265792
rect 121512 265752 121518 265764
rect 272150 265752 272156 265764
rect 272208 265752 272214 265804
rect 331306 265752 331312 265804
rect 331364 265792 331370 265804
rect 491294 265792 491300 265804
rect 331364 265764 491300 265792
rect 331364 265752 331370 265764
rect 491294 265752 491300 265764
rect 491352 265752 491358 265804
rect 39298 265684 39304 265736
rect 39356 265724 39362 265736
rect 258166 265724 258172 265736
rect 39356 265696 258172 265724
rect 39356 265684 39362 265696
rect 258166 265684 258172 265696
rect 258224 265684 258230 265736
rect 338206 265684 338212 265736
rect 338264 265724 338270 265736
rect 535454 265724 535460 265736
rect 338264 265696 535460 265724
rect 338264 265684 338270 265696
rect 535454 265684 535460 265696
rect 535512 265684 535518 265736
rect 11054 265616 11060 265668
rect 11112 265656 11118 265668
rect 247678 265656 247684 265668
rect 11112 265628 247684 265656
rect 11112 265616 11118 265628
rect 247678 265616 247684 265628
rect 247736 265616 247742 265668
rect 342438 265616 342444 265668
rect 342496 265656 342502 265668
rect 560938 265656 560944 265668
rect 342496 265628 560944 265656
rect 342496 265616 342502 265628
rect 560938 265616 560944 265628
rect 560996 265616 561002 265668
rect 314746 264392 314752 264444
rect 314804 264432 314810 264444
rect 389174 264432 389180 264444
rect 314804 264404 389180 264432
rect 314804 264392 314810 264404
rect 389174 264392 389180 264404
rect 389232 264392 389238 264444
rect 154574 264324 154580 264376
rect 154632 264364 154638 264376
rect 277670 264364 277676 264376
rect 154632 264336 277676 264364
rect 154632 264324 154638 264336
rect 277670 264324 277676 264336
rect 277728 264324 277734 264376
rect 323486 264324 323492 264376
rect 323544 264364 323550 264376
rect 440234 264364 440240 264376
rect 323544 264336 440240 264364
rect 323544 264324 323550 264336
rect 440234 264324 440240 264336
rect 440292 264324 440298 264376
rect 149054 264256 149060 264308
rect 149112 264296 149118 264308
rect 276106 264296 276112 264308
rect 149112 264268 276112 264296
rect 149112 264256 149118 264268
rect 276106 264256 276112 264268
rect 276164 264256 276170 264308
rect 323578 264256 323584 264308
rect 323636 264296 323642 264308
rect 442994 264296 443000 264308
rect 323636 264268 443000 264296
rect 323636 264256 323642 264268
rect 442994 264256 443000 264268
rect 443052 264256 443058 264308
rect 69014 264188 69020 264240
rect 69072 264228 69078 264240
rect 263870 264228 263876 264240
rect 69072 264200 263876 264228
rect 69072 264188 69078 264200
rect 263870 264188 263876 264200
rect 263928 264188 263934 264240
rect 345290 264188 345296 264240
rect 345348 264228 345354 264240
rect 574094 264228 574100 264240
rect 345348 264200 574100 264228
rect 345348 264188 345354 264200
rect 574094 264188 574100 264200
rect 574152 264188 574158 264240
rect 316586 263100 316592 263152
rect 316644 263140 316650 263152
rect 393314 263140 393320 263152
rect 316644 263112 393320 263140
rect 316644 263100 316650 263112
rect 393314 263100 393320 263112
rect 393372 263100 393378 263152
rect 316494 263032 316500 263084
rect 316552 263072 316558 263084
rect 397454 263072 397460 263084
rect 316552 263044 397460 263072
rect 316552 263032 316558 263044
rect 397454 263032 397460 263044
rect 397512 263032 397518 263084
rect 142154 262964 142160 263016
rect 142212 263004 142218 263016
rect 275278 263004 275284 263016
rect 142212 262976 275284 263004
rect 142212 262964 142218 262976
rect 275278 262964 275284 262976
rect 275336 262964 275342 263016
rect 323302 262964 323308 263016
rect 323360 263004 323366 263016
rect 436094 263004 436100 263016
rect 323360 262976 436100 263004
rect 323360 262964 323366 262976
rect 436094 262964 436100 262976
rect 436152 262964 436158 263016
rect 52454 262896 52460 262948
rect 52512 262936 52518 262948
rect 261018 262936 261024 262948
rect 52512 262908 261024 262936
rect 52512 262896 52518 262908
rect 261018 262896 261024 262908
rect 261076 262896 261082 262948
rect 323394 262896 323400 262948
rect 323452 262936 323458 262948
rect 441614 262936 441620 262948
rect 323452 262908 441620 262936
rect 323452 262896 323458 262908
rect 441614 262896 441620 262908
rect 441672 262896 441678 262948
rect 7558 262828 7564 262880
rect 7616 262868 7622 262880
rect 252738 262868 252744 262880
rect 7616 262840 252744 262868
rect 7616 262828 7622 262840
rect 252738 262828 252744 262840
rect 252796 262828 252802 262880
rect 324498 262828 324504 262880
rect 324556 262868 324562 262880
rect 449894 262868 449900 262880
rect 324556 262840 449900 262868
rect 324556 262828 324562 262840
rect 449894 262828 449900 262840
rect 449952 262828 449958 262880
rect 314654 261808 314660 261860
rect 314712 261848 314718 261860
rect 390646 261848 390652 261860
rect 314712 261820 390652 261848
rect 314712 261808 314718 261820
rect 390646 261808 390652 261820
rect 390704 261808 390710 261860
rect 212534 261740 212540 261792
rect 212592 261780 212598 261792
rect 287330 261780 287336 261792
rect 212592 261752 287336 261780
rect 212592 261740 212598 261752
rect 287330 261740 287336 261752
rect 287388 261740 287394 261792
rect 316402 261740 316408 261792
rect 316460 261780 316466 261792
rect 398834 261780 398840 261792
rect 316460 261752 398840 261780
rect 316460 261740 316466 261752
rect 398834 261740 398840 261752
rect 398892 261740 398898 261792
rect 158714 261672 158720 261724
rect 158772 261712 158778 261724
rect 277578 261712 277584 261724
rect 158772 261684 277584 261712
rect 158772 261672 158778 261684
rect 277578 261672 277584 261684
rect 277636 261672 277642 261724
rect 323210 261672 323216 261724
rect 323268 261712 323274 261724
rect 438854 261712 438860 261724
rect 323268 261684 438860 261712
rect 323268 261672 323274 261684
rect 438854 261672 438860 261684
rect 438912 261672 438918 261724
rect 144914 261604 144920 261656
rect 144972 261644 144978 261656
rect 276014 261644 276020 261656
rect 144972 261616 276020 261644
rect 144972 261604 144978 261616
rect 276014 261604 276020 261616
rect 276072 261604 276078 261656
rect 334618 261604 334624 261656
rect 334676 261644 334682 261656
rect 506474 261644 506480 261656
rect 334676 261616 506480 261644
rect 334676 261604 334682 261616
rect 506474 261604 506480 261616
rect 506532 261604 506538 261656
rect 73154 261536 73160 261588
rect 73212 261576 73218 261588
rect 263778 261576 263784 261588
rect 73212 261548 263784 261576
rect 73212 261536 73218 261548
rect 263778 261536 263784 261548
rect 263836 261536 263842 261588
rect 334526 261536 334532 261588
rect 334584 261576 334590 261588
rect 510614 261576 510620 261588
rect 334584 261548 510620 261576
rect 334584 261536 334590 261548
rect 510614 261536 510620 261548
rect 510672 261536 510678 261588
rect 13814 261468 13820 261520
rect 13872 261508 13878 261520
rect 254394 261508 254400 261520
rect 13872 261480 254400 261508
rect 13872 261468 13878 261480
rect 254394 261468 254400 261480
rect 254452 261468 254458 261520
rect 343818 261468 343824 261520
rect 343876 261508 343882 261520
rect 569954 261508 569960 261520
rect 343876 261480 569960 261508
rect 343876 261468 343882 261480
rect 569954 261468 569960 261480
rect 570012 261468 570018 261520
rect 124214 260380 124220 260432
rect 124272 260420 124278 260432
rect 251910 260420 251916 260432
rect 124272 260392 251916 260420
rect 124272 260380 124278 260392
rect 251910 260380 251916 260392
rect 251968 260380 251974 260432
rect 63494 260312 63500 260364
rect 63552 260352 63558 260364
rect 262674 260352 262680 260364
rect 63552 260324 262680 260352
rect 63552 260312 63558 260324
rect 262674 260312 262680 260324
rect 262732 260312 262738 260364
rect 316218 260312 316224 260364
rect 316276 260352 316282 260364
rect 391934 260352 391940 260364
rect 316276 260324 391940 260352
rect 316276 260312 316282 260324
rect 391934 260312 391940 260324
rect 391992 260312 391998 260364
rect 39390 260244 39396 260296
rect 39448 260284 39454 260296
rect 256878 260284 256884 260296
rect 39448 260256 256884 260284
rect 39448 260244 39454 260256
rect 256878 260244 256884 260256
rect 256936 260244 256942 260296
rect 316310 260244 316316 260296
rect 316368 260284 316374 260296
rect 396074 260284 396080 260296
rect 316368 260256 396080 260284
rect 316368 260244 316374 260256
rect 396074 260244 396080 260256
rect 396132 260244 396138 260296
rect 30374 260176 30380 260228
rect 30432 260216 30438 260228
rect 257246 260216 257252 260228
rect 30432 260188 257252 260216
rect 30432 260176 30438 260188
rect 257246 260176 257252 260188
rect 257304 260176 257310 260228
rect 339862 260176 339868 260228
rect 339920 260216 339926 260228
rect 542354 260216 542360 260228
rect 339920 260188 542360 260216
rect 339920 260176 339926 260188
rect 542354 260176 542360 260188
rect 542412 260176 542418 260228
rect 19334 260108 19340 260160
rect 19392 260148 19398 260160
rect 246298 260148 246304 260160
rect 19392 260120 246304 260148
rect 19392 260108 19398 260120
rect 246298 260108 246304 260120
rect 246356 260108 246362 260160
rect 342346 260108 342352 260160
rect 342404 260148 342410 260160
rect 558914 260148 558920 260160
rect 342404 260120 558920 260148
rect 342404 260108 342410 260120
rect 558914 260108 558920 260120
rect 558972 260108 558978 260160
rect 362218 259360 362224 259412
rect 362276 259400 362282 259412
rect 579798 259400 579804 259412
rect 362276 259372 579804 259400
rect 362276 259360 362282 259372
rect 579798 259360 579804 259372
rect 579856 259360 579862 259412
rect 176654 258816 176660 258868
rect 176712 258856 176718 258868
rect 266998 258856 267004 258868
rect 176712 258828 267004 258856
rect 176712 258816 176718 258828
rect 266998 258816 267004 258828
rect 267056 258816 267062 258868
rect 323118 258816 323124 258868
rect 323176 258856 323182 258868
rect 434714 258856 434720 258868
rect 323176 258828 434720 258856
rect 323176 258816 323182 258828
rect 434714 258816 434720 258828
rect 434772 258816 434778 258868
rect 217594 258748 217600 258800
rect 217652 258788 217658 258800
rect 346486 258788 346492 258800
rect 217652 258760 346492 258788
rect 217652 258748 217658 258760
rect 346486 258748 346492 258760
rect 346544 258748 346550 258800
rect 173894 258680 173900 258732
rect 173952 258720 173958 258732
rect 280614 258720 280620 258732
rect 173952 258692 280620 258720
rect 173952 258680 173958 258692
rect 280614 258680 280620 258692
rect 280672 258680 280678 258732
rect 339770 258680 339776 258732
rect 339828 258720 339834 258732
rect 539686 258720 539692 258732
rect 339828 258692 539692 258720
rect 339828 258680 339834 258692
rect 539686 258680 539692 258692
rect 539744 258680 539750 258732
rect 218606 257592 218612 257644
rect 218664 257632 218670 257644
rect 287238 257632 287244 257644
rect 218664 257604 287244 257632
rect 218664 257592 218670 257604
rect 287238 257592 287244 257604
rect 287296 257592 287302 257644
rect 117314 257524 117320 257576
rect 117372 257564 117378 257576
rect 251818 257564 251824 257576
rect 117372 257536 251824 257564
rect 117372 257524 117378 257536
rect 251818 257524 251824 257536
rect 251876 257524 251882 257576
rect 106274 257456 106280 257508
rect 106332 257496 106338 257508
rect 261478 257496 261484 257508
rect 106332 257468 261484 257496
rect 106332 257456 106338 257468
rect 261478 257456 261484 257468
rect 261536 257456 261542 257508
rect 334434 257456 334440 257508
rect 334492 257496 334498 257508
rect 509234 257496 509240 257508
rect 334492 257468 509240 257496
rect 334492 257456 334498 257468
rect 509234 257456 509240 257468
rect 509292 257456 509298 257508
rect 25590 257388 25596 257440
rect 25648 257428 25654 257440
rect 255406 257428 255412 257440
rect 25648 257400 255412 257428
rect 25648 257388 25654 257400
rect 255406 257388 255412 257400
rect 255464 257388 255470 257440
rect 339678 257388 339684 257440
rect 339736 257428 339742 257440
rect 540974 257428 540980 257440
rect 339736 257400 540980 257428
rect 339736 257388 339742 257400
rect 540974 257388 540980 257400
rect 541032 257388 541038 257440
rect 23474 257320 23480 257372
rect 23532 257360 23538 257372
rect 255498 257360 255504 257372
rect 23532 257332 255504 257360
rect 23532 257320 23538 257332
rect 255498 257320 255504 257332
rect 255556 257320 255562 257372
rect 339586 257320 339592 257372
rect 339644 257360 339650 257372
rect 545114 257360 545120 257372
rect 339644 257332 545120 257360
rect 339644 257320 339650 257332
rect 545114 257320 545120 257332
rect 545172 257320 545178 257372
rect 318978 256368 318984 256420
rect 319036 256408 319042 256420
rect 413278 256408 413284 256420
rect 319036 256380 413284 256408
rect 319036 256368 319042 256380
rect 413278 256368 413284 256380
rect 413336 256368 413342 256420
rect 217134 256300 217140 256352
rect 217192 256340 217198 256352
rect 348418 256340 348424 256352
rect 217192 256312 348424 256340
rect 217192 256300 217198 256312
rect 348418 256300 348424 256312
rect 348476 256300 348482 256352
rect 122834 256232 122840 256284
rect 122892 256272 122898 256284
rect 272058 256272 272064 256284
rect 122892 256244 272064 256272
rect 122892 256232 122898 256244
rect 272058 256232 272064 256244
rect 272116 256232 272122 256284
rect 320266 256232 320272 256284
rect 320324 256272 320330 256284
rect 425054 256272 425060 256284
rect 320324 256244 425060 256272
rect 320324 256232 320330 256244
rect 425054 256232 425060 256244
rect 425112 256232 425118 256284
rect 118694 256164 118700 256216
rect 118752 256204 118758 256216
rect 271966 256204 271972 256216
rect 118752 256176 271972 256204
rect 118752 256164 118758 256176
rect 271966 256164 271972 256176
rect 272024 256164 272030 256216
rect 321738 256164 321744 256216
rect 321796 256204 321802 256216
rect 431954 256204 431960 256216
rect 321796 256176 431960 256204
rect 321796 256164 321802 256176
rect 431954 256164 431960 256176
rect 432012 256164 432018 256216
rect 92474 256096 92480 256148
rect 92532 256136 92538 256148
rect 266722 256136 266728 256148
rect 92532 256108 266728 256136
rect 92532 256096 92538 256108
rect 266722 256096 266728 256108
rect 266780 256096 266786 256148
rect 323026 256096 323032 256148
rect 323084 256136 323090 256148
rect 440326 256136 440332 256148
rect 323084 256108 440332 256136
rect 323084 256096 323090 256108
rect 440326 256096 440332 256108
rect 440384 256096 440390 256148
rect 77386 256028 77392 256080
rect 77444 256068 77450 256080
rect 265158 256068 265164 256080
rect 77444 256040 265164 256068
rect 77444 256028 77450 256040
rect 265158 256028 265164 256040
rect 265216 256028 265222 256080
rect 325694 256028 325700 256080
rect 325752 256068 325758 256080
rect 454034 256068 454040 256080
rect 325752 256040 454040 256068
rect 325752 256028 325758 256040
rect 454034 256028 454040 256040
rect 454092 256028 454098 256080
rect 17954 255960 17960 256012
rect 18012 256000 18018 256012
rect 255866 256000 255872 256012
rect 18012 255972 255872 256000
rect 18012 255960 18018 255972
rect 255866 255960 255872 255972
rect 255924 255960 255930 256012
rect 334342 255960 334348 256012
rect 334400 256000 334406 256012
rect 506566 256000 506572 256012
rect 334400 255972 506572 256000
rect 334400 255960 334406 255972
rect 506566 255960 506572 255972
rect 506624 255960 506630 256012
rect 169754 254872 169760 254924
rect 169812 254912 169818 254924
rect 280522 254912 280528 254924
rect 169812 254884 280528 254912
rect 169812 254872 169818 254884
rect 280522 254872 280528 254884
rect 280580 254872 280586 254924
rect 217410 254804 217416 254856
rect 217468 254844 217474 254856
rect 345198 254844 345204 254856
rect 217468 254816 345204 254844
rect 217468 254804 217474 254816
rect 345198 254804 345204 254816
rect 345256 254804 345262 254856
rect 3326 254736 3332 254788
rect 3384 254776 3390 254788
rect 8938 254776 8944 254788
rect 3384 254748 8944 254776
rect 3384 254736 3390 254748
rect 8938 254736 8944 254748
rect 8996 254736 9002 254788
rect 95234 254736 95240 254788
rect 95292 254776 95298 254788
rect 267826 254776 267832 254788
rect 95292 254748 267832 254776
rect 95292 254736 95298 254748
rect 267826 254736 267832 254748
rect 267884 254736 267890 254788
rect 316126 254736 316132 254788
rect 316184 254776 316190 254788
rect 398926 254776 398932 254788
rect 316184 254748 398932 254776
rect 316184 254736 316190 254748
rect 398926 254736 398932 254748
rect 398984 254736 398990 254788
rect 91094 254668 91100 254720
rect 91152 254708 91158 254720
rect 266538 254708 266544 254720
rect 91152 254680 266544 254708
rect 91152 254668 91158 254680
rect 266538 254668 266544 254680
rect 266596 254668 266602 254720
rect 324406 254668 324412 254720
rect 324464 254708 324470 254720
rect 443638 254708 443644 254720
rect 324464 254680 443644 254708
rect 324464 254668 324470 254680
rect 443638 254668 443644 254680
rect 443696 254668 443702 254720
rect 88334 254600 88340 254652
rect 88392 254640 88398 254652
rect 264238 254640 264244 254652
rect 88392 254612 264244 254640
rect 88392 254600 88398 254612
rect 264238 254600 264244 254612
rect 264296 254600 264302 254652
rect 343634 254600 343640 254652
rect 343692 254640 343698 254652
rect 564526 254640 564532 254652
rect 343692 254612 564532 254640
rect 343692 254600 343698 254612
rect 564526 254600 564532 254612
rect 564584 254600 564590 254652
rect 86954 254532 86960 254584
rect 87012 254572 87018 254584
rect 266630 254572 266636 254584
rect 87012 254544 266636 254572
rect 87012 254532 87018 254544
rect 266630 254532 266636 254544
rect 266688 254532 266694 254584
rect 343726 254532 343732 254584
rect 343784 254572 343790 254584
rect 567194 254572 567200 254584
rect 343784 254544 567200 254572
rect 343784 254532 343790 254544
rect 567194 254532 567200 254544
rect 567252 254532 567258 254584
rect 302602 253784 302608 253836
rect 302660 253824 302666 253836
rect 360286 253824 360292 253836
rect 302660 253796 360292 253824
rect 302660 253784 302666 253796
rect 360286 253784 360292 253796
rect 360344 253784 360350 253836
rect 304074 253716 304080 253768
rect 304132 253756 304138 253768
rect 367186 253756 367192 253768
rect 304132 253728 367192 253756
rect 304132 253716 304138 253728
rect 367186 253716 367192 253728
rect 367244 253716 367250 253768
rect 301130 253648 301136 253700
rect 301188 253688 301194 253700
rect 364518 253688 364524 253700
rect 301188 253660 364524 253688
rect 301188 253648 301194 253660
rect 364518 253648 364524 253660
rect 364576 253648 364582 253700
rect 301038 253580 301044 253632
rect 301096 253620 301102 253632
rect 368474 253620 368480 253632
rect 301096 253592 368480 253620
rect 301096 253580 301102 253592
rect 368474 253580 368480 253592
rect 368532 253580 368538 253632
rect 176746 253512 176752 253564
rect 176804 253552 176810 253564
rect 280430 253552 280436 253564
rect 176804 253524 280436 253552
rect 176804 253512 176810 253524
rect 280430 253512 280436 253524
rect 280488 253512 280494 253564
rect 316034 253512 316040 253564
rect 316092 253552 316098 253564
rect 394694 253552 394700 253564
rect 316092 253524 394700 253552
rect 316092 253512 316098 253524
rect 394694 253512 394700 253524
rect 394752 253512 394758 253564
rect 218514 253444 218520 253496
rect 218572 253484 218578 253496
rect 347774 253484 347780 253496
rect 218572 253456 347780 253484
rect 218572 253444 218578 253456
rect 347774 253444 347780 253456
rect 347832 253444 347838 253496
rect 118786 253376 118792 253428
rect 118844 253416 118850 253428
rect 270586 253416 270592 253428
rect 118844 253388 270592 253416
rect 118844 253376 118850 253388
rect 270586 253376 270592 253388
rect 270644 253376 270650 253428
rect 322934 253376 322940 253428
rect 322992 253416 322998 253428
rect 437474 253416 437480 253428
rect 322992 253388 437480 253416
rect 322992 253376 322998 253388
rect 437474 253376 437480 253388
rect 437532 253376 437538 253428
rect 110506 253308 110512 253360
rect 110564 253348 110570 253360
rect 271046 253348 271052 253360
rect 110564 253320 271052 253348
rect 110564 253308 110570 253320
rect 271046 253308 271052 253320
rect 271104 253308 271110 253360
rect 332778 253308 332784 253360
rect 332836 253348 332842 253360
rect 496078 253348 496084 253360
rect 332836 253320 496084 253348
rect 332836 253308 332842 253320
rect 496078 253308 496084 253320
rect 496136 253308 496142 253360
rect 85574 253240 85580 253292
rect 85632 253280 85638 253292
rect 266446 253280 266452 253292
rect 85632 253252 266452 253280
rect 85632 253240 85638 253252
rect 266446 253240 266452 253252
rect 266504 253240 266510 253292
rect 332686 253240 332692 253292
rect 332744 253280 332750 253292
rect 499574 253280 499580 253292
rect 332744 253252 499580 253280
rect 332744 253240 332750 253252
rect 499574 253240 499580 253252
rect 499632 253240 499638 253292
rect 80054 253172 80060 253224
rect 80112 253212 80118 253224
rect 265066 253212 265072 253224
rect 80112 253184 265072 253212
rect 80112 253172 80118 253184
rect 265066 253172 265072 253184
rect 265124 253172 265130 253224
rect 336826 253172 336832 253224
rect 336884 253212 336890 253224
rect 528554 253212 528560 253224
rect 336884 253184 528560 253212
rect 336884 253172 336890 253184
rect 528554 253172 528560 253184
rect 528612 253172 528618 253224
rect 172514 252084 172520 252136
rect 172572 252124 172578 252136
rect 280338 252124 280344 252136
rect 172572 252096 280344 252124
rect 172572 252084 172578 252096
rect 280338 252084 280344 252096
rect 280396 252084 280402 252136
rect 321646 252084 321652 252136
rect 321704 252124 321710 252136
rect 427814 252124 427820 252136
rect 321704 252096 427820 252124
rect 321704 252084 321710 252096
rect 427814 252084 427820 252096
rect 427872 252084 427878 252136
rect 160186 252016 160192 252068
rect 160244 252056 160250 252068
rect 277486 252056 277492 252068
rect 160244 252028 277492 252056
rect 160244 252016 160250 252028
rect 277486 252016 277492 252028
rect 277544 252016 277550 252068
rect 321554 252016 321560 252068
rect 321612 252056 321618 252068
rect 432046 252056 432052 252068
rect 321612 252028 432052 252056
rect 321612 252016 321618 252028
rect 432046 252016 432052 252028
rect 432104 252016 432110 252068
rect 155954 251948 155960 252000
rect 156012 251988 156018 252000
rect 277394 251988 277400 252000
rect 156012 251960 277400 251988
rect 156012 251948 156018 251960
rect 277394 251948 277400 251960
rect 277452 251948 277458 252000
rect 327166 251948 327172 252000
rect 327224 251988 327230 252000
rect 466454 251988 466460 252000
rect 327224 251960 466460 251988
rect 327224 251948 327230 251960
rect 466454 251948 466460 251960
rect 466512 251948 466518 252000
rect 49694 251880 49700 251932
rect 49752 251920 49758 251932
rect 259638 251920 259644 251932
rect 49752 251892 259644 251920
rect 49752 251880 49758 251892
rect 259638 251880 259644 251892
rect 259696 251880 259702 251932
rect 339494 251880 339500 251932
rect 339552 251920 339558 251932
rect 538214 251920 538220 251932
rect 339552 251892 538220 251920
rect 339552 251880 339558 251892
rect 538214 251880 538220 251892
rect 538272 251880 538278 251932
rect 46198 251812 46204 251864
rect 46256 251852 46262 251864
rect 259546 251852 259552 251864
rect 46256 251824 259552 251852
rect 46256 251812 46262 251824
rect 259546 251812 259552 251824
rect 259604 251812 259610 251864
rect 345106 251812 345112 251864
rect 345164 251852 345170 251864
rect 578234 251852 578240 251864
rect 345164 251824 578240 251852
rect 345164 251812 345170 251824
rect 578234 251812 578240 251824
rect 578292 251812 578298 251864
rect 309502 251132 309508 251184
rect 309560 251172 309566 251184
rect 365806 251172 365812 251184
rect 309560 251144 365812 251172
rect 309560 251132 309566 251144
rect 365806 251132 365812 251144
rect 365864 251132 365870 251184
rect 306742 251064 306748 251116
rect 306800 251104 306806 251116
rect 363230 251104 363236 251116
rect 306800 251076 363236 251104
rect 306800 251064 306806 251076
rect 363230 251064 363236 251076
rect 363288 251064 363294 251116
rect 306834 250996 306840 251048
rect 306892 251036 306898 251048
rect 364610 251036 364616 251048
rect 306892 251008 364616 251036
rect 306892 250996 306898 251008
rect 364610 250996 364616 251008
rect 364668 250996 364674 251048
rect 306926 250928 306932 250980
rect 306984 250968 306990 250980
rect 364702 250968 364708 250980
rect 306984 250940 364708 250968
rect 306984 250928 306990 250940
rect 364702 250928 364708 250940
rect 364760 250928 364766 250980
rect 305546 250860 305552 250912
rect 305604 250900 305610 250912
rect 363322 250900 363328 250912
rect 305604 250872 363328 250900
rect 305604 250860 305610 250872
rect 363322 250860 363328 250872
rect 363380 250860 363386 250912
rect 209866 250792 209872 250844
rect 209924 250832 209930 250844
rect 286134 250832 286140 250844
rect 209924 250804 286140 250832
rect 209924 250792 209930 250804
rect 286134 250792 286140 250804
rect 286192 250792 286198 250844
rect 311894 250792 311900 250844
rect 311952 250832 311958 250844
rect 371234 250832 371240 250844
rect 311952 250804 371240 250832
rect 311952 250792 311958 250804
rect 371234 250792 371240 250804
rect 371292 250792 371298 250844
rect 135346 250724 135352 250776
rect 135404 250764 135410 250776
rect 273714 250764 273720 250776
rect 135404 250736 273720 250764
rect 135404 250724 135410 250736
rect 273714 250724 273720 250736
rect 273772 250724 273778 250776
rect 303890 250724 303896 250776
rect 303948 250764 303954 250776
rect 365898 250764 365904 250776
rect 303948 250736 365904 250764
rect 303948 250724 303954 250736
rect 365898 250724 365904 250736
rect 365956 250724 365962 250776
rect 60734 250656 60740 250708
rect 60792 250696 60798 250708
rect 255958 250696 255964 250708
rect 60792 250668 255964 250696
rect 60792 250656 60798 250668
rect 255958 250656 255964 250668
rect 256016 250656 256022 250708
rect 318886 250656 318892 250708
rect 318944 250696 318950 250708
rect 416774 250696 416780 250708
rect 318944 250668 416780 250696
rect 318944 250656 318950 250668
rect 416774 250656 416780 250668
rect 416832 250656 416838 250708
rect 67634 250588 67640 250640
rect 67692 250628 67698 250640
rect 263686 250628 263692 250640
rect 67692 250600 263692 250628
rect 67692 250588 67698 250600
rect 263686 250588 263692 250600
rect 263744 250588 263750 250640
rect 330294 250588 330300 250640
rect 330352 250628 330358 250640
rect 484394 250628 484400 250640
rect 330352 250600 484400 250628
rect 330352 250588 330358 250600
rect 484394 250588 484400 250600
rect 484452 250588 484458 250640
rect 66254 250520 66260 250572
rect 66312 250560 66318 250572
rect 262582 250560 262588 250572
rect 66312 250532 262588 250560
rect 66312 250520 66318 250532
rect 262582 250520 262588 250532
rect 262640 250520 262646 250572
rect 334250 250520 334256 250572
rect 334308 250560 334314 250572
rect 503714 250560 503720 250572
rect 334308 250532 503720 250560
rect 334308 250520 334314 250532
rect 503714 250520 503720 250532
rect 503772 250520 503778 250572
rect 52546 250452 52552 250504
rect 52604 250492 52610 250504
rect 260926 250492 260932 250504
rect 52604 250464 260932 250492
rect 52604 250452 52610 250464
rect 260926 250452 260932 250464
rect 260984 250452 260990 250504
rect 345014 250452 345020 250504
rect 345072 250492 345078 250504
rect 576854 250492 576860 250504
rect 345072 250464 576860 250492
rect 345072 250452 345078 250464
rect 576854 250452 576860 250464
rect 576912 250452 576918 250504
rect 309594 250384 309600 250436
rect 309652 250424 309658 250436
rect 365714 250424 365720 250436
rect 309652 250396 365720 250424
rect 309652 250384 309658 250396
rect 365714 250384 365720 250396
rect 365772 250384 365778 250436
rect 305638 250316 305644 250368
rect 305696 250356 305702 250368
rect 360194 250356 360200 250368
rect 305696 250328 360200 250356
rect 305696 250316 305702 250328
rect 360194 250316 360200 250328
rect 360252 250316 360258 250368
rect 318794 249432 318800 249484
rect 318852 249472 318858 249484
rect 414014 249472 414020 249484
rect 318852 249444 414020 249472
rect 318852 249432 318858 249444
rect 414014 249432 414020 249444
rect 414072 249432 414078 249484
rect 185026 249364 185032 249416
rect 185084 249404 185090 249416
rect 282178 249404 282184 249416
rect 185084 249376 282184 249404
rect 185084 249364 185090 249376
rect 282178 249364 282184 249376
rect 282236 249364 282242 249416
rect 340138 249364 340144 249416
rect 340196 249404 340202 249416
rect 455414 249404 455420 249416
rect 340196 249376 455420 249404
rect 340196 249364 340202 249376
rect 455414 249364 455420 249376
rect 455472 249364 455478 249416
rect 217226 249296 217232 249348
rect 217284 249336 217290 249348
rect 346394 249336 346400 249348
rect 217284 249308 346400 249336
rect 217284 249296 217290 249308
rect 346394 249296 346400 249308
rect 346452 249296 346458 249348
rect 82814 249228 82820 249280
rect 82872 249268 82878 249280
rect 264974 249268 264980 249280
rect 82872 249240 264980 249268
rect 82872 249228 82878 249240
rect 264974 249228 264980 249240
rect 265032 249228 265038 249280
rect 327074 249228 327080 249280
rect 327132 249268 327138 249280
rect 467834 249268 467840 249280
rect 327132 249240 467840 249268
rect 327132 249228 327138 249240
rect 467834 249228 467840 249240
rect 467892 249228 467898 249280
rect 74534 249160 74540 249212
rect 74592 249200 74598 249212
rect 264330 249200 264336 249212
rect 74592 249172 264336 249200
rect 74592 249160 74598 249172
rect 264330 249160 264336 249172
rect 264388 249160 264394 249212
rect 328546 249160 328552 249212
rect 328604 249200 328610 249212
rect 477494 249200 477500 249212
rect 328604 249172 477500 249200
rect 328604 249160 328610 249172
rect 477494 249160 477500 249172
rect 477552 249160 477558 249212
rect 62114 249092 62120 249144
rect 62172 249132 62178 249144
rect 262490 249132 262496 249144
rect 62172 249104 262496 249132
rect 62172 249092 62178 249104
rect 262490 249092 262496 249104
rect 262548 249092 262554 249144
rect 334158 249092 334164 249144
rect 334216 249132 334222 249144
rect 511994 249132 512000 249144
rect 334216 249104 512000 249132
rect 334216 249092 334222 249104
rect 511994 249092 512000 249104
rect 512052 249092 512058 249144
rect 57330 249024 57336 249076
rect 57388 249064 57394 249076
rect 261386 249064 261392 249076
rect 57388 249036 261392 249064
rect 57388 249024 57394 249036
rect 261386 249024 261392 249036
rect 261444 249024 261450 249076
rect 335446 249024 335452 249076
rect 335504 249064 335510 249076
rect 520274 249064 520280 249076
rect 335504 249036 520280 249064
rect 335504 249024 335510 249036
rect 520274 249024 520280 249036
rect 520332 249024 520338 249076
rect 306650 248344 306656 248396
rect 306708 248384 306714 248396
rect 362954 248384 362960 248396
rect 306708 248356 362960 248384
rect 306708 248344 306714 248356
rect 362954 248344 362960 248356
rect 363012 248344 363018 248396
rect 302418 248276 302424 248328
rect 302476 248316 302482 248328
rect 359458 248316 359464 248328
rect 302476 248288 359464 248316
rect 302476 248276 302482 248288
rect 359458 248276 359464 248288
rect 359516 248276 359522 248328
rect 306558 248208 306564 248260
rect 306616 248248 306622 248260
rect 364426 248248 364432 248260
rect 306616 248220 364432 248248
rect 306616 248208 306622 248220
rect 364426 248208 364432 248220
rect 364484 248208 364490 248260
rect 305086 248140 305092 248192
rect 305144 248180 305150 248192
rect 363046 248180 363052 248192
rect 305144 248152 363052 248180
rect 305144 248140 305150 248152
rect 363046 248140 363052 248152
rect 363104 248140 363110 248192
rect 305454 248072 305460 248124
rect 305512 248112 305518 248124
rect 364334 248112 364340 248124
rect 305512 248084 364340 248112
rect 305512 248072 305518 248084
rect 364334 248072 364340 248084
rect 364392 248072 364398 248124
rect 201586 248004 201592 248056
rect 201644 248044 201650 248056
rect 284754 248044 284760 248056
rect 201644 248016 284760 248044
rect 201644 248004 201650 248016
rect 284754 248004 284760 248016
rect 284812 248004 284818 248056
rect 302510 248004 302516 248056
rect 302568 248044 302574 248056
rect 361942 248044 361948 248056
rect 302568 248016 361948 248044
rect 302568 248004 302574 248016
rect 361942 248004 361948 248016
rect 362000 248004 362006 248056
rect 140774 247936 140780 247988
rect 140832 247976 140838 247988
rect 275186 247976 275192 247988
rect 140832 247948 275192 247976
rect 140832 247936 140838 247948
rect 275186 247936 275192 247948
rect 275244 247936 275250 247988
rect 302326 247936 302332 247988
rect 302384 247976 302390 247988
rect 372706 247976 372712 247988
rect 302384 247948 372712 247976
rect 302384 247936 302390 247948
rect 372706 247936 372712 247948
rect 372764 247936 372770 247988
rect 89714 247868 89720 247920
rect 89772 247908 89778 247920
rect 253198 247908 253204 247920
rect 89772 247880 253204 247908
rect 89772 247868 89778 247880
rect 253198 247868 253204 247880
rect 253256 247868 253262 247920
rect 320174 247868 320180 247920
rect 320232 247908 320238 247920
rect 423766 247908 423772 247920
rect 320232 247880 423772 247908
rect 320232 247868 320238 247880
rect 423766 247868 423772 247880
rect 423824 247868 423830 247920
rect 41414 247800 41420 247852
rect 41472 247840 41478 247852
rect 258534 247840 258540 247852
rect 41472 247812 258540 247840
rect 41472 247800 41478 247812
rect 258534 247800 258540 247812
rect 258592 247800 258598 247852
rect 332594 247800 332600 247852
rect 332652 247840 332658 247852
rect 502334 247840 502340 247852
rect 332652 247812 502340 247840
rect 332652 247800 332658 247812
rect 502334 247800 502340 247812
rect 502392 247800 502398 247852
rect 35158 247732 35164 247784
rect 35216 247772 35222 247784
rect 257154 247772 257160 247784
rect 35216 247744 257160 247772
rect 35216 247732 35222 247744
rect 257154 247732 257160 247744
rect 257212 247732 257218 247784
rect 333974 247732 333980 247784
rect 334032 247772 334038 247784
rect 505094 247772 505100 247784
rect 334032 247744 505100 247772
rect 334032 247732 334038 247744
rect 505094 247732 505100 247744
rect 505152 247732 505158 247784
rect 4154 247664 4160 247716
rect 4212 247704 4218 247716
rect 252646 247704 252652 247716
rect 4212 247676 252652 247704
rect 4212 247664 4218 247676
rect 252646 247664 252652 247676
rect 252704 247664 252710 247716
rect 334066 247664 334072 247716
rect 334124 247704 334130 247716
rect 507854 247704 507860 247716
rect 334124 247676 507860 247704
rect 334124 247664 334130 247676
rect 507854 247664 507860 247676
rect 507912 247664 507918 247716
rect 308030 247596 308036 247648
rect 308088 247636 308094 247648
rect 363138 247636 363144 247648
rect 308088 247608 363144 247636
rect 308088 247596 308094 247608
rect 363138 247596 363144 247608
rect 363196 247596 363202 247648
rect 303706 247528 303712 247580
rect 303764 247568 303770 247580
rect 356698 247568 356704 247580
rect 303764 247540 356704 247568
rect 303764 247528 303770 247540
rect 356698 247528 356704 247540
rect 356756 247528 356762 247580
rect 355686 247460 355692 247512
rect 355744 247500 355750 247512
rect 369854 247500 369860 247512
rect 355744 247472 369860 247500
rect 355744 247460 355750 247472
rect 369854 247460 369860 247472
rect 369912 247460 369918 247512
rect 211890 246780 211896 246832
rect 211948 246820 211954 246832
rect 262306 246820 262312 246832
rect 211948 246792 262312 246820
rect 211948 246780 211954 246792
rect 262306 246780 262312 246792
rect 262364 246780 262370 246832
rect 175274 246712 175280 246764
rect 175332 246752 175338 246764
rect 280246 246752 280252 246764
rect 175332 246724 280252 246752
rect 175332 246712 175338 246724
rect 280246 246712 280252 246724
rect 280304 246712 280310 246764
rect 120074 246644 120080 246696
rect 120132 246684 120138 246696
rect 272334 246684 272340 246696
rect 120132 246656 272340 246684
rect 120132 246644 120138 246656
rect 272334 246644 272340 246656
rect 272392 246644 272398 246696
rect 328454 246644 328460 246696
rect 328512 246684 328518 246696
rect 471974 246684 471980 246696
rect 328512 246656 471980 246684
rect 328512 246644 328518 246656
rect 471974 246644 471980 246656
rect 472032 246644 472038 246696
rect 104894 246576 104900 246628
rect 104952 246616 104958 246628
rect 269206 246616 269212 246628
rect 104952 246588 269212 246616
rect 104952 246576 104958 246588
rect 269206 246576 269212 246588
rect 269264 246576 269270 246628
rect 330110 246576 330116 246628
rect 330168 246616 330174 246628
rect 480254 246616 480260 246628
rect 330168 246588 480260 246616
rect 330168 246576 330174 246588
rect 480254 246576 480260 246588
rect 480312 246576 480318 246628
rect 85666 246508 85672 246560
rect 85724 246548 85730 246560
rect 266814 246548 266820 246560
rect 85724 246520 266820 246548
rect 85724 246508 85730 246520
rect 266814 246508 266820 246520
rect 266872 246508 266878 246560
rect 330202 246508 330208 246560
rect 330260 246548 330266 246560
rect 483014 246548 483020 246560
rect 330260 246520 483020 246548
rect 330260 246508 330266 246520
rect 483014 246508 483020 246520
rect 483072 246508 483078 246560
rect 64874 246440 64880 246492
rect 64932 246480 64938 246492
rect 262398 246480 262404 246492
rect 64932 246452 262404 246480
rect 64932 246440 64938 246452
rect 262398 246440 262404 246452
rect 262456 246440 262462 246492
rect 330018 246440 330024 246492
rect 330076 246480 330082 246492
rect 485774 246480 485780 246492
rect 330076 246452 485780 246480
rect 330076 246440 330082 246452
rect 485774 246440 485780 246452
rect 485832 246440 485838 246492
rect 48314 246372 48320 246424
rect 48372 246412 48378 246424
rect 260006 246412 260012 246424
rect 48372 246384 260012 246412
rect 48372 246372 48378 246384
rect 260006 246372 260012 246384
rect 260064 246372 260070 246424
rect 331214 246372 331220 246424
rect 331272 246412 331278 246424
rect 492674 246412 492680 246424
rect 331272 246384 492680 246412
rect 331272 246372 331278 246384
rect 492674 246372 492680 246384
rect 492732 246372 492738 246424
rect 6914 246304 6920 246356
rect 6972 246344 6978 246356
rect 253014 246344 253020 246356
rect 6972 246316 253020 246344
rect 6972 246304 6978 246316
rect 253014 246304 253020 246316
rect 253072 246304 253078 246356
rect 335354 246304 335360 246356
rect 335412 246344 335418 246356
rect 516134 246344 516140 246356
rect 335412 246316 516140 246344
rect 335412 246304 335418 246316
rect 516134 246304 516140 246316
rect 516192 246304 516198 246356
rect 355410 245556 355416 245608
rect 355468 245596 355474 245608
rect 372798 245596 372804 245608
rect 355468 245568 372804 245596
rect 355468 245556 355474 245568
rect 372798 245556 372804 245568
rect 372856 245556 372862 245608
rect 307938 245488 307944 245540
rect 307996 245528 308002 245540
rect 361574 245528 361580 245540
rect 307996 245500 361580 245528
rect 307996 245488 308002 245500
rect 361574 245488 361580 245500
rect 361632 245488 361638 245540
rect 307754 245420 307760 245472
rect 307812 245460 307818 245472
rect 361758 245460 361764 245472
rect 307812 245432 361764 245460
rect 307812 245420 307818 245432
rect 361758 245420 361764 245432
rect 361816 245420 361822 245472
rect 307846 245352 307852 245404
rect 307904 245392 307910 245404
rect 361850 245392 361856 245404
rect 307904 245364 361856 245392
rect 307904 245352 307910 245364
rect 361850 245352 361856 245364
rect 361908 245352 361914 245404
rect 198090 245284 198096 245336
rect 198148 245324 198154 245336
rect 283374 245324 283380 245336
rect 198148 245296 283380 245324
rect 198148 245284 198154 245296
rect 283374 245284 283380 245296
rect 283432 245284 283438 245336
rect 306374 245284 306380 245336
rect 306432 245324 306438 245336
rect 361666 245324 361672 245336
rect 306432 245296 361672 245324
rect 306432 245284 306438 245296
rect 361666 245284 361672 245296
rect 361724 245284 361730 245336
rect 171226 245216 171232 245268
rect 171284 245256 171290 245268
rect 280706 245256 280712 245268
rect 171284 245228 280712 245256
rect 171284 245216 171290 245228
rect 280706 245216 280712 245228
rect 280764 245216 280770 245268
rect 302234 245216 302240 245268
rect 302292 245256 302298 245268
rect 360930 245256 360936 245268
rect 302292 245228 360936 245256
rect 302292 245216 302298 245228
rect 360930 245216 360936 245228
rect 360988 245216 360994 245268
rect 168466 245148 168472 245200
rect 168524 245188 168530 245200
rect 279234 245188 279240 245200
rect 168524 245160 279240 245188
rect 168524 245148 168530 245160
rect 279234 245148 279240 245160
rect 279292 245148 279298 245200
rect 324314 245148 324320 245200
rect 324372 245188 324378 245200
rect 445754 245188 445760 245200
rect 324372 245160 445760 245188
rect 324372 245148 324378 245160
rect 445754 245148 445760 245160
rect 445812 245148 445818 245200
rect 109034 245080 109040 245132
rect 109092 245120 109098 245132
rect 269666 245120 269672 245132
rect 109092 245092 269672 245120
rect 109092 245080 109098 245092
rect 269666 245080 269672 245092
rect 269724 245080 269730 245132
rect 329926 245080 329932 245132
rect 329984 245120 329990 245132
rect 481726 245120 481732 245132
rect 329984 245092 481732 245120
rect 329984 245080 329990 245092
rect 481726 245080 481732 245092
rect 481784 245080 481790 245132
rect 100754 245012 100760 245064
rect 100812 245052 100818 245064
rect 268286 245052 268292 245064
rect 100812 245024 268292 245052
rect 100812 245012 100818 245024
rect 268286 245012 268292 245024
rect 268344 245012 268350 245064
rect 329834 245012 329840 245064
rect 329892 245052 329898 245064
rect 481634 245052 481640 245064
rect 329892 245024 481640 245052
rect 329892 245012 329898 245024
rect 481634 245012 481640 245024
rect 481692 245012 481698 245064
rect 60826 244944 60832 244996
rect 60884 244984 60890 244996
rect 262766 244984 262772 244996
rect 60884 244956 262772 244984
rect 60884 244944 60890 244956
rect 262766 244944 262772 244956
rect 262824 244944 262830 244996
rect 338114 244944 338120 244996
rect 338172 244984 338178 244996
rect 534074 244984 534080 244996
rect 338172 244956 534080 244984
rect 338172 244944 338178 244956
rect 534074 244944 534080 244956
rect 534132 244944 534138 244996
rect 31754 244876 31760 244928
rect 31812 244916 31818 244928
rect 250438 244916 250444 244928
rect 31812 244888 250444 244916
rect 31812 244876 31818 244888
rect 250438 244876 250444 244888
rect 250496 244876 250502 244928
rect 342254 244876 342260 244928
rect 342312 244916 342318 244928
rect 560294 244916 560300 244928
rect 342312 244888 560300 244916
rect 342312 244876 342318 244888
rect 560294 244876 560300 244888
rect 560352 244876 560358 244928
rect 355318 244808 355324 244860
rect 355376 244848 355382 244860
rect 365990 244848 365996 244860
rect 355376 244820 365996 244848
rect 355376 244808 355382 244820
rect 365990 244808 365996 244820
rect 366048 244808 366054 244860
rect 355594 244740 355600 244792
rect 355652 244780 355658 244792
rect 364794 244780 364800 244792
rect 355652 244752 364800 244780
rect 355652 244740 355658 244752
rect 364794 244740 364800 244752
rect 364852 244740 364858 244792
rect 355502 244604 355508 244656
rect 355560 244644 355566 244656
rect 358170 244644 358176 244656
rect 355560 244616 358176 244644
rect 355560 244604 355566 244616
rect 358170 244604 358176 244616
rect 358228 244604 358234 244656
rect 356974 243924 356980 243976
rect 357032 243964 357038 243976
rect 367922 243964 367928 243976
rect 357032 243936 367928 243964
rect 357032 243924 357038 243936
rect 367922 243924 367928 243936
rect 367980 243924 367986 243976
rect 299658 243856 299664 243908
rect 299716 243896 299722 243908
rect 362402 243896 362408 243908
rect 299716 243868 362408 243896
rect 299716 243856 299722 243868
rect 362402 243856 362408 243868
rect 362460 243856 362466 243908
rect 299474 243788 299480 243840
rect 299532 243828 299538 243840
rect 362218 243828 362224 243840
rect 299532 243800 362224 243828
rect 299532 243788 299538 243800
rect 362218 243788 362224 243800
rect 362276 243788 362282 243840
rect 298554 243720 298560 243772
rect 298612 243760 298618 243772
rect 361022 243760 361028 243772
rect 298612 243732 361028 243760
rect 298612 243720 298618 243732
rect 361022 243720 361028 243732
rect 361080 243720 361086 243772
rect 300854 243652 300860 243704
rect 300912 243692 300918 243704
rect 363782 243692 363788 243704
rect 300912 243664 363788 243692
rect 300912 243652 300918 243664
rect 363782 243652 363788 243664
rect 363840 243652 363846 243704
rect 219250 243584 219256 243636
rect 219308 243624 219314 243636
rect 297174 243624 297180 243636
rect 219308 243596 297180 243624
rect 219308 243584 219314 243596
rect 297174 243584 297180 243596
rect 297232 243584 297238 243636
rect 300946 243584 300952 243636
rect 301004 243624 301010 243636
rect 366082 243624 366088 243636
rect 301004 243596 366088 243624
rect 301004 243584 301010 243596
rect 366082 243584 366088 243596
rect 366140 243584 366146 243636
rect 217502 243516 217508 243568
rect 217560 243556 217566 243568
rect 297266 243556 297272 243568
rect 217560 243528 297272 243556
rect 217560 243516 217566 243528
rect 297266 243516 297272 243528
rect 297324 243516 297330 243568
rect 299566 243516 299572 243568
rect 299624 243556 299630 243568
rect 369302 243556 369308 243568
rect 299624 243528 369308 243556
rect 299624 243516 299630 243528
rect 369302 243516 369308 243528
rect 369360 243516 369366 243568
rect 356790 242156 356796 242208
rect 356848 242196 356854 242208
rect 369210 242196 369216 242208
rect 356848 242168 369216 242196
rect 356848 242156 356854 242168
rect 369210 242156 369216 242168
rect 369268 242156 369274 242208
rect 577590 206932 577596 206984
rect 577648 206972 577654 206984
rect 579614 206972 579620 206984
rect 577648 206944 579620 206972
rect 577648 206932 577654 206944
rect 579614 206932 579620 206944
rect 579672 206932 579678 206984
rect 3050 202784 3056 202836
rect 3108 202824 3114 202836
rect 196710 202824 196716 202836
rect 3108 202796 196716 202824
rect 3108 202784 3114 202796
rect 196710 202784 196716 202796
rect 196768 202784 196774 202836
rect 214374 195644 214380 195696
rect 214432 195684 214438 195696
rect 217318 195684 217324 195696
rect 214432 195656 217324 195684
rect 214432 195644 214438 195656
rect 217318 195644 217324 195656
rect 217376 195644 217382 195696
rect 215754 193128 215760 193180
rect 215812 193168 215818 193180
rect 218698 193168 218704 193180
rect 215812 193140 218704 193168
rect 215812 193128 215818 193140
rect 218698 193128 218704 193140
rect 218756 193128 218762 193180
rect 3510 188980 3516 189032
rect 3568 189020 3574 189032
rect 203610 189020 203616 189032
rect 3568 188992 203616 189020
rect 3568 188980 3574 188992
rect 203610 188980 203616 188992
rect 203668 188980 203674 189032
rect 210602 188980 210608 189032
rect 210660 189020 210666 189032
rect 216674 189020 216680 189032
rect 210660 188992 216680 189020
rect 210660 188980 210666 188992
rect 216674 188980 216680 188992
rect 216732 188980 216738 189032
rect 374730 179324 374736 179376
rect 374788 179364 374794 179376
rect 580166 179364 580172 179376
rect 374788 179336 580172 179364
rect 374788 179324 374794 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 371970 166948 371976 167000
rect 372028 166988 372034 167000
rect 579614 166988 579620 167000
rect 372028 166960 579620 166988
rect 372028 166948 372034 166960
rect 579614 166948 579620 166960
rect 579672 166948 579678 167000
rect 213638 159604 213644 159656
rect 213696 159644 213702 159656
rect 256694 159644 256700 159656
rect 213696 159616 256700 159644
rect 213696 159604 213702 159616
rect 256694 159604 256700 159616
rect 256752 159604 256758 159656
rect 214466 159536 214472 159588
rect 214524 159576 214530 159588
rect 260834 159576 260840 159588
rect 214524 159548 260840 159576
rect 214524 159536 214530 159548
rect 260834 159536 260840 159548
rect 260892 159536 260898 159588
rect 322934 159536 322940 159588
rect 322992 159576 322998 159588
rect 358078 159576 358084 159588
rect 322992 159548 358084 159576
rect 322992 159536 322998 159548
rect 358078 159536 358084 159548
rect 358136 159536 358142 159588
rect 217870 159468 217876 159520
rect 217928 159508 217934 159520
rect 264974 159508 264980 159520
rect 217928 159480 264980 159508
rect 217928 159468 217934 159480
rect 264974 159468 264980 159480
rect 265032 159468 265038 159520
rect 320082 159468 320088 159520
rect 320140 159508 320146 159520
rect 357986 159508 357992 159520
rect 320140 159480 357992 159508
rect 320140 159468 320146 159480
rect 357986 159468 357992 159480
rect 358044 159468 358050 159520
rect 212166 159400 212172 159452
rect 212224 159440 212230 159452
rect 259454 159440 259460 159452
rect 212224 159412 259460 159440
rect 212224 159400 212230 159412
rect 259454 159400 259460 159412
rect 259512 159400 259518 159452
rect 314654 159400 314660 159452
rect 314712 159440 314718 159452
rect 357894 159440 357900 159452
rect 314712 159412 357900 159440
rect 314712 159400 314718 159412
rect 357894 159400 357900 159412
rect 357952 159400 357958 159452
rect 214834 159332 214840 159384
rect 214892 159372 214898 159384
rect 282914 159372 282920 159384
rect 214892 159344 282920 159372
rect 214892 159332 214898 159344
rect 282914 159332 282920 159344
rect 282972 159332 282978 159384
rect 310422 159332 310428 159384
rect 310480 159372 310486 159384
rect 357710 159372 357716 159384
rect 310480 159344 357716 159372
rect 310480 159332 310486 159344
rect 357710 159332 357716 159344
rect 357768 159332 357774 159384
rect 300946 159264 300952 159316
rect 301004 159304 301010 159316
rect 357802 159304 357808 159316
rect 301004 159276 357808 159304
rect 301004 159264 301010 159276
rect 357802 159264 357808 159276
rect 357860 159264 357866 159316
rect 279234 159196 279240 159248
rect 279292 159236 279298 159248
rect 360746 159236 360752 159248
rect 279292 159208 360752 159236
rect 279292 159196 279298 159208
rect 360746 159196 360752 159208
rect 360804 159196 360810 159248
rect 278130 159128 278136 159180
rect 278188 159168 278194 159180
rect 360654 159168 360660 159180
rect 278188 159140 360660 159168
rect 278188 159128 278194 159140
rect 360654 159128 360660 159140
rect 360712 159128 360718 159180
rect 275830 159060 275836 159112
rect 275888 159100 275894 159112
rect 359274 159100 359280 159112
rect 275888 159072 359280 159100
rect 275888 159060 275894 159072
rect 359274 159060 359280 159072
rect 359332 159060 359338 159112
rect 277026 158992 277032 159044
rect 277084 159032 277090 159044
rect 360838 159032 360844 159044
rect 277084 159004 360844 159032
rect 277084 158992 277090 159004
rect 360838 158992 360844 159004
rect 360896 158992 360902 159044
rect 274450 158924 274456 158976
rect 274508 158964 274514 158976
rect 359366 158964 359372 158976
rect 274508 158936 359372 158964
rect 274508 158924 274514 158936
rect 359366 158924 359372 158936
rect 359424 158924 359430 158976
rect 267642 158856 267648 158908
rect 267700 158896 267706 158908
rect 370498 158896 370504 158908
rect 267700 158868 370504 158896
rect 267700 158856 267706 158868
rect 370498 158856 370504 158868
rect 370556 158856 370562 158908
rect 262858 158788 262864 158840
rect 262916 158828 262922 158840
rect 366358 158828 366364 158840
rect 262916 158800 366364 158828
rect 262916 158788 262922 158800
rect 366358 158788 366364 158800
rect 366416 158788 366422 158840
rect 211706 158720 211712 158772
rect 211764 158760 211770 158772
rect 239582 158760 239588 158772
rect 211764 158732 239588 158760
rect 211764 158720 211770 158732
rect 239582 158720 239588 158732
rect 239640 158720 239646 158772
rect 258534 158720 258540 158772
rect 258592 158760 258598 158772
rect 363690 158760 363696 158772
rect 258592 158732 363696 158760
rect 258592 158720 258598 158732
rect 363690 158720 363696 158732
rect 363748 158720 363754 158772
rect 213178 158652 213184 158704
rect 213236 158692 213242 158704
rect 238110 158692 238116 158704
rect 213236 158664 238116 158692
rect 213236 158652 213242 158664
rect 238110 158652 238116 158664
rect 238168 158652 238174 158704
rect 308674 158652 308680 158704
rect 308732 158692 308738 158704
rect 320082 158692 320088 158704
rect 308732 158664 320088 158692
rect 308732 158652 308738 158664
rect 320082 158652 320088 158664
rect 320140 158652 320146 158704
rect 211982 158584 211988 158636
rect 212040 158624 212046 158636
rect 230474 158624 230480 158636
rect 212040 158596 230480 158624
rect 212040 158584 212046 158596
rect 230474 158584 230480 158596
rect 230532 158584 230538 158636
rect 306098 158584 306104 158636
rect 306156 158624 306162 158636
rect 314654 158624 314660 158636
rect 306156 158596 314660 158624
rect 306156 158584 306162 158596
rect 314654 158584 314660 158596
rect 314712 158584 314718 158636
rect 215938 158516 215944 158568
rect 215996 158556 216002 158568
rect 235994 158556 236000 158568
rect 215996 158528 236000 158556
rect 215996 158516 216002 158528
rect 235994 158516 236000 158528
rect 236052 158516 236058 158568
rect 259546 158516 259552 158568
rect 259604 158556 259610 158568
rect 367830 158556 367836 158568
rect 259604 158528 367836 158556
rect 259604 158516 259610 158528
rect 367830 158516 367836 158528
rect 367888 158516 367894 158568
rect 213362 158448 213368 158500
rect 213420 158488 213426 158500
rect 234706 158488 234712 158500
rect 213420 158460 234712 158488
rect 213420 158448 213426 158460
rect 234706 158448 234712 158460
rect 234764 158448 234770 158500
rect 265986 158448 265992 158500
rect 266044 158488 266050 158500
rect 369118 158488 369124 158500
rect 266044 158460 369124 158488
rect 266044 158448 266050 158460
rect 369118 158448 369124 158460
rect 369176 158448 369182 158500
rect 219066 158380 219072 158432
rect 219124 158420 219130 158432
rect 242986 158420 242992 158432
rect 219124 158392 242992 158420
rect 219124 158380 219130 158392
rect 242986 158380 242992 158392
rect 243044 158380 243050 158432
rect 268746 158380 268752 158432
rect 268804 158420 268810 158432
rect 357434 158420 357440 158432
rect 268804 158392 357440 158420
rect 268804 158380 268810 158392
rect 357434 158380 357440 158392
rect 357492 158380 357498 158432
rect 216030 158312 216036 158364
rect 216088 158352 216094 158364
rect 242894 158352 242900 158364
rect 216088 158324 242900 158352
rect 216088 158312 216094 158324
rect 242894 158312 242900 158324
rect 242952 158312 242958 158364
rect 270218 158312 270224 158364
rect 270276 158352 270282 158364
rect 357618 158352 357624 158364
rect 270276 158324 357624 158352
rect 270276 158312 270282 158324
rect 357618 158312 357624 158324
rect 357676 158312 357682 158364
rect 216398 158244 216404 158296
rect 216456 158284 216462 158296
rect 245654 158284 245660 158296
rect 216456 158256 245660 158284
rect 216456 158244 216462 158256
rect 245654 158244 245660 158256
rect 245712 158244 245718 158296
rect 271138 158244 271144 158296
rect 271196 158284 271202 158296
rect 357526 158284 357532 158296
rect 271196 158256 357532 158284
rect 271196 158244 271202 158256
rect 357526 158244 357532 158256
rect 357584 158244 357590 158296
rect 214558 158176 214564 158228
rect 214616 158216 214622 158228
rect 247034 158216 247040 158228
rect 214616 158188 247040 158216
rect 214616 158176 214622 158188
rect 247034 158176 247040 158188
rect 247092 158176 247098 158228
rect 298922 158176 298928 158228
rect 298980 158216 298986 158228
rect 373442 158216 373448 158228
rect 298980 158188 373448 158216
rect 298980 158176 298986 158188
rect 373442 158176 373448 158188
rect 373500 158176 373506 158228
rect 217962 158108 217968 158160
rect 218020 158148 218026 158160
rect 251174 158148 251180 158160
rect 218020 158120 251180 158148
rect 218020 158108 218026 158120
rect 251174 158108 251180 158120
rect 251232 158108 251238 158160
rect 303522 158108 303528 158160
rect 303580 158148 303586 158160
rect 310422 158148 310428 158160
rect 303580 158120 310428 158148
rect 303580 158108 303586 158120
rect 310422 158108 310428 158120
rect 310480 158108 310486 158160
rect 321186 158108 321192 158160
rect 321244 158148 321250 158160
rect 360378 158148 360384 158160
rect 321244 158120 360384 158148
rect 321244 158108 321250 158120
rect 360378 158108 360384 158120
rect 360436 158108 360442 158160
rect 216306 158040 216312 158092
rect 216364 158080 216370 158092
rect 249794 158080 249800 158092
rect 216364 158052 249800 158080
rect 216364 158040 216370 158052
rect 249794 158040 249800 158052
rect 249852 158040 249858 158092
rect 313458 158040 313464 158092
rect 313516 158080 313522 158092
rect 358998 158080 359004 158092
rect 313516 158052 359004 158080
rect 313516 158040 313522 158052
rect 358998 158040 359004 158052
rect 359056 158040 359062 158092
rect 218974 157972 218980 158024
rect 219032 158012 219038 158024
rect 252554 158012 252560 158024
rect 219032 157984 252560 158012
rect 219032 157972 219038 157984
rect 252554 157972 252560 157984
rect 252612 157972 252618 158024
rect 315850 157972 315856 158024
rect 315908 158012 315914 158024
rect 359090 158012 359096 158024
rect 315908 157984 359096 158012
rect 315908 157972 315914 157984
rect 359090 157972 359096 157984
rect 359148 157972 359154 158024
rect 214742 157904 214748 157956
rect 214800 157944 214806 157956
rect 233234 157944 233240 157956
rect 214800 157916 233240 157944
rect 214800 157904 214806 157916
rect 233234 157904 233240 157916
rect 233292 157904 233298 157956
rect 318610 157904 318616 157956
rect 318668 157944 318674 157956
rect 359182 157944 359188 157956
rect 318668 157916 359188 157944
rect 318668 157904 318674 157916
rect 359182 157904 359188 157916
rect 359240 157904 359246 157956
rect 218882 157836 218888 157888
rect 218940 157876 218946 157888
rect 234614 157876 234620 157888
rect 218940 157848 234620 157876
rect 218940 157836 218946 157848
rect 234614 157836 234620 157848
rect 234672 157836 234678 157888
rect 272242 157836 272248 157888
rect 272300 157876 272306 157888
rect 322934 157876 322940 157888
rect 272300 157848 322940 157876
rect 272300 157836 272306 157848
rect 322934 157836 322940 157848
rect 322992 157836 322998 157888
rect 323394 157836 323400 157888
rect 323452 157876 323458 157888
rect 360470 157876 360476 157888
rect 323452 157848 360476 157876
rect 323452 157836 323458 157848
rect 360470 157836 360476 157848
rect 360528 157836 360534 157888
rect 215846 157768 215852 157820
rect 215904 157808 215910 157820
rect 229094 157808 229100 157820
rect 215904 157780 229100 157808
rect 215904 157768 215910 157780
rect 229094 157768 229100 157780
rect 229152 157768 229158 157820
rect 325970 157768 325976 157820
rect 326028 157808 326034 157820
rect 360562 157808 360568 157820
rect 326028 157780 360568 157808
rect 326028 157768 326034 157780
rect 360562 157768 360568 157780
rect 360620 157768 360626 157820
rect 240686 157700 240692 157752
rect 240744 157740 240750 157752
rect 373350 157740 373356 157752
rect 240744 157712 373356 157740
rect 240744 157700 240750 157712
rect 373350 157700 373356 157712
rect 373408 157700 373414 157752
rect 256602 157632 256608 157684
rect 256660 157672 256666 157684
rect 366542 157672 366548 157684
rect 256660 157644 366548 157672
rect 256660 157632 256666 157644
rect 366542 157632 366548 157644
rect 366600 157632 366606 157684
rect 261754 157360 261760 157412
rect 261812 157400 261818 157412
rect 317046 157400 317052 157412
rect 261812 157372 317052 157400
rect 261812 157360 261818 157372
rect 317046 157360 317052 157372
rect 317104 157360 317110 157412
rect 250162 157292 250168 157344
rect 250220 157332 250226 157344
rect 368842 157332 368848 157344
rect 250220 157304 368848 157332
rect 250220 157292 250226 157304
rect 368842 157292 368848 157304
rect 368900 157292 368906 157344
rect 248322 157224 248328 157276
rect 248380 157264 248386 157276
rect 364978 157264 364984 157276
rect 248380 157236 364984 157264
rect 248380 157224 248386 157236
rect 364978 157224 364984 157236
rect 365036 157224 365042 157276
rect 257154 157156 257160 157208
rect 257212 157196 257218 157208
rect 367646 157196 367652 157208
rect 257212 157168 367652 157196
rect 257212 157156 257218 157168
rect 367646 157156 367652 157168
rect 367704 157156 367710 157208
rect 255958 157088 255964 157140
rect 256016 157128 256022 157140
rect 364886 157128 364892 157140
rect 256016 157100 364892 157128
rect 256016 157088 256022 157100
rect 364886 157088 364892 157100
rect 364944 157088 364950 157140
rect 258626 157020 258632 157072
rect 258684 157060 258690 157072
rect 367554 157060 367560 157072
rect 258684 157032 367560 157060
rect 258684 157020 258690 157032
rect 367554 157020 367560 157032
rect 367612 157020 367618 157072
rect 260650 156952 260656 157004
rect 260708 156992 260714 157004
rect 367462 156992 367468 157004
rect 260708 156964 367468 156992
rect 260708 156952 260714 156964
rect 367462 156952 367468 156964
rect 367520 156952 367526 157004
rect 276106 156884 276112 156936
rect 276164 156924 276170 156936
rect 368934 156924 368940 156936
rect 276164 156896 368940 156924
rect 276164 156884 276170 156896
rect 368934 156884 368940 156896
rect 368992 156884 368998 156936
rect 281350 156816 281356 156868
rect 281408 156856 281414 156868
rect 371786 156856 371792 156868
rect 281408 156828 371792 156856
rect 281408 156816 281414 156828
rect 371786 156816 371792 156828
rect 371844 156816 371850 156868
rect 286226 156748 286232 156800
rect 286284 156788 286290 156800
rect 371694 156788 371700 156800
rect 286284 156760 371700 156788
rect 286284 156748 286290 156760
rect 371694 156748 371700 156760
rect 371752 156748 371758 156800
rect 273346 156680 273352 156732
rect 273404 156720 273410 156732
rect 358814 156720 358820 156732
rect 273404 156692 358820 156720
rect 273404 156680 273410 156692
rect 358814 156680 358820 156692
rect 358872 156680 358878 156732
rect 291010 156612 291016 156664
rect 291068 156652 291074 156664
rect 370406 156652 370412 156664
rect 291068 156624 370412 156652
rect 291068 156612 291074 156624
rect 370406 156612 370412 156624
rect 370464 156612 370470 156664
rect 296254 156544 296260 156596
rect 296312 156584 296318 156596
rect 359550 156584 359556 156596
rect 296312 156556 359556 156584
rect 296312 156544 296318 156556
rect 359550 156544 359556 156556
rect 359608 156544 359614 156596
rect 317046 156476 317052 156528
rect 317104 156516 317110 156528
rect 370682 156516 370688 156528
rect 317104 156488 370688 156516
rect 317104 156476 317110 156488
rect 370682 156476 370688 156488
rect 370740 156476 370746 156528
rect 311250 156408 311256 156460
rect 311308 156448 311314 156460
rect 358906 156448 358912 156460
rect 311308 156420 358912 156448
rect 311308 156408 311314 156420
rect 358906 156408 358912 156420
rect 358964 156408 358970 156460
rect 245378 155864 245384 155916
rect 245436 155904 245442 155916
rect 366174 155904 366180 155916
rect 245436 155876 366180 155904
rect 245436 155864 245442 155876
rect 366174 155864 366180 155876
rect 366232 155864 366238 155916
rect 212074 155796 212080 155848
rect 212132 155836 212138 155848
rect 237374 155836 237380 155848
rect 212132 155808 237380 155836
rect 212132 155796 212138 155808
rect 237374 155796 237380 155808
rect 237432 155796 237438 155848
rect 253566 155796 253572 155848
rect 253624 155836 253630 155848
rect 368658 155836 368664 155848
rect 253624 155808 368664 155836
rect 253624 155796 253630 155808
rect 368658 155796 368664 155808
rect 368716 155796 368722 155848
rect 213546 155728 213552 155780
rect 213604 155768 213610 155780
rect 241514 155768 241520 155780
rect 213604 155740 241520 155768
rect 213604 155728 213610 155740
rect 241514 155728 241520 155740
rect 241572 155728 241578 155780
rect 252094 155728 252100 155780
rect 252152 155768 252158 155780
rect 362034 155768 362040 155780
rect 252152 155740 362040 155768
rect 252152 155728 252158 155740
rect 362034 155728 362040 155740
rect 362092 155728 362098 155780
rect 216214 155660 216220 155712
rect 216272 155700 216278 155712
rect 248414 155700 248420 155712
rect 216272 155672 248420 155700
rect 216272 155660 216278 155672
rect 248414 155660 248420 155672
rect 248472 155660 248478 155712
rect 261938 155660 261944 155712
rect 261996 155700 262002 155712
rect 367370 155700 367376 155712
rect 261996 155672 367376 155700
rect 261996 155660 262002 155672
rect 367370 155660 367376 155672
rect 367428 155660 367434 155712
rect 210970 155592 210976 155644
rect 211028 155632 211034 155644
rect 267826 155632 267832 155644
rect 211028 155604 267832 155632
rect 211028 155592 211034 155604
rect 267826 155592 267832 155604
rect 267884 155592 267890 155644
rect 268930 155592 268936 155644
rect 268988 155632 268994 155644
rect 373074 155632 373080 155644
rect 268988 155604 373080 155632
rect 268988 155592 268994 155604
rect 373074 155592 373080 155604
rect 373132 155592 373138 155644
rect 213454 155524 213460 155576
rect 213512 155564 213518 155576
rect 253934 155564 253940 155576
rect 213512 155536 253940 155564
rect 213512 155524 213518 155536
rect 253934 155524 253940 155536
rect 253992 155524 253998 155576
rect 266722 155524 266728 155576
rect 266780 155564 266786 155576
rect 369946 155564 369952 155576
rect 266780 155536 369952 155564
rect 266780 155524 266786 155536
rect 369946 155524 369952 155536
rect 370004 155524 370010 155576
rect 210878 155456 210884 155508
rect 210936 155496 210942 155508
rect 270494 155496 270500 155508
rect 210936 155468 270500 155496
rect 210936 155456 210942 155468
rect 270494 155456 270500 155468
rect 270552 155456 270558 155508
rect 271046 155456 271052 155508
rect 271104 155496 271110 155508
rect 372982 155496 372988 155508
rect 271104 155468 372988 155496
rect 271104 155456 271110 155468
rect 372982 155456 372988 155468
rect 373040 155456 373046 155508
rect 210694 155388 210700 155440
rect 210752 155428 210758 155440
rect 255314 155428 255320 155440
rect 210752 155400 255320 155428
rect 210752 155388 210758 155400
rect 255314 155388 255320 155400
rect 255372 155388 255378 155440
rect 265986 155388 265992 155440
rect 266044 155428 266050 155440
rect 367278 155428 367284 155440
rect 266044 155400 367284 155428
rect 266044 155388 266050 155400
rect 367278 155388 367284 155400
rect 367336 155388 367342 155440
rect 218790 155320 218796 155372
rect 218848 155360 218854 155372
rect 263594 155360 263600 155372
rect 218848 155332 263600 155360
rect 218848 155320 218854 155332
rect 263594 155320 263600 155332
rect 263652 155320 263658 155372
rect 264422 155320 264428 155372
rect 264480 155360 264486 155372
rect 363506 155360 363512 155372
rect 264480 155332 363512 155360
rect 264480 155320 264486 155332
rect 363506 155320 363512 155332
rect 363564 155320 363570 155372
rect 212258 155252 212264 155304
rect 212316 155292 212322 155304
rect 273254 155292 273260 155304
rect 212316 155264 273260 155292
rect 212316 155252 212322 155264
rect 273254 155252 273260 155264
rect 273312 155252 273318 155304
rect 274450 155252 274456 155304
rect 274508 155292 274514 155304
rect 368750 155292 368756 155304
rect 274508 155264 368756 155292
rect 274508 155252 274514 155264
rect 368750 155252 368756 155264
rect 368808 155252 368814 155304
rect 213270 155184 213276 155236
rect 213328 155224 213334 155236
rect 274634 155224 274640 155236
rect 213328 155196 274640 155224
rect 213328 155184 213334 155196
rect 274634 155184 274640 155196
rect 274692 155184 274698 155236
rect 278682 155184 278688 155236
rect 278740 155224 278746 155236
rect 371602 155224 371608 155236
rect 278740 155196 371608 155224
rect 278740 155184 278746 155196
rect 371602 155184 371608 155196
rect 371660 155184 371666 155236
rect 217502 155116 217508 155168
rect 217560 155156 217566 155168
rect 278774 155156 278780 155168
rect 217560 155128 278780 155156
rect 217560 155116 217566 155128
rect 278774 155116 278780 155128
rect 278832 155116 278838 155168
rect 284110 155116 284116 155168
rect 284168 155156 284174 155168
rect 371510 155156 371516 155168
rect 284168 155128 371516 155156
rect 284168 155116 284174 155128
rect 371510 155116 371516 155128
rect 371568 155116 371574 155168
rect 219158 155048 219164 155100
rect 219216 155088 219222 155100
rect 287054 155088 287060 155100
rect 219216 155060 287060 155088
rect 219216 155048 219222 155060
rect 287054 155048 287060 155060
rect 287112 155048 287118 155100
rect 288250 155048 288256 155100
rect 288308 155088 288314 155100
rect 371418 155088 371424 155100
rect 288308 155060 371424 155088
rect 288308 155048 288314 155060
rect 371418 155048 371424 155060
rect 371476 155048 371482 155100
rect 216122 154980 216128 155032
rect 216180 155020 216186 155032
rect 277394 155020 277400 155032
rect 216180 154992 277400 155020
rect 216180 154980 216186 154992
rect 277394 154980 277400 154992
rect 277452 154980 277458 155032
rect 293586 154980 293592 155032
rect 293644 155020 293650 155032
rect 367738 155020 367744 155032
rect 293644 154992 367744 155020
rect 293644 154980 293650 154992
rect 367738 154980 367744 154992
rect 367796 154980 367802 155032
rect 253658 154504 253664 154556
rect 253716 154544 253722 154556
rect 370222 154544 370228 154556
rect 253716 154516 370228 154544
rect 253716 154504 253722 154516
rect 370222 154504 370228 154516
rect 370280 154504 370286 154556
rect 263962 154436 263968 154488
rect 264020 154476 264026 154488
rect 372890 154476 372896 154488
rect 264020 154448 372896 154476
rect 264020 154436 264026 154448
rect 372890 154436 372896 154448
rect 372948 154436 372954 154488
rect 299474 153960 299480 154012
rect 299532 154000 299538 154012
rect 363598 154000 363604 154012
rect 299532 153972 363604 154000
rect 299532 153960 299538 153972
rect 363598 153960 363604 153972
rect 363656 153960 363662 154012
rect 295334 153892 295340 153944
rect 295392 153932 295398 153944
rect 362218 153932 362224 153944
rect 295392 153904 362224 153932
rect 295392 153892 295398 153904
rect 362218 153892 362224 153904
rect 362276 153892 362282 153944
rect 288434 153824 288440 153876
rect 288492 153864 288498 153876
rect 361022 153864 361028 153876
rect 288492 153836 361028 153864
rect 288492 153824 288498 153836
rect 361022 153824 361028 153836
rect 361080 153824 361086 153876
rect 345750 152532 345756 152584
rect 345808 152572 345814 152584
rect 369210 152572 369216 152584
rect 345808 152544 369216 152572
rect 345808 152532 345814 152544
rect 369210 152532 369216 152544
rect 369268 152532 369274 152584
rect 300854 152464 300860 152516
rect 300912 152504 300918 152516
rect 370590 152504 370596 152516
rect 300912 152476 370596 152504
rect 300912 152464 300918 152476
rect 370590 152464 370596 152476
rect 370648 152464 370654 152516
rect 3510 150356 3516 150408
rect 3568 150396 3574 150408
rect 197998 150396 198004 150408
rect 3568 150368 198004 150396
rect 3568 150356 3574 150368
rect 197998 150356 198004 150368
rect 198056 150356 198062 150408
rect 3510 137912 3516 137964
rect 3568 137952 3574 137964
rect 206278 137952 206284 137964
rect 3568 137924 206284 137952
rect 3568 137912 3574 137924
rect 206278 137912 206284 137924
rect 206336 137912 206342 137964
rect 3418 97928 3424 97980
rect 3476 97968 3482 97980
rect 192478 97968 192484 97980
rect 3476 97940 192484 97968
rect 3476 97928 3482 97940
rect 192478 97928 192484 97940
rect 192536 97928 192542 97980
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 200758 85524 200764 85536
rect 3200 85496 200764 85524
rect 3200 85484 3206 85496
rect 200758 85484 200764 85496
rect 200816 85484 200822 85536
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 207658 71720 207664 71732
rect 3476 71692 207664 71720
rect 3476 71680 3482 71692
rect 207658 71680 207664 71692
rect 207716 71680 207722 71732
rect 373258 60664 373264 60716
rect 373316 60704 373322 60716
rect 580166 60704 580172 60716
rect 373316 60676 580172 60704
rect 373316 60664 373322 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 25498 59344 25504 59356
rect 3108 59316 25504 59344
rect 3108 59304 3114 59316
rect 25498 59304 25504 59316
rect 25556 59304 25562 59356
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 199378 45540 199384 45552
rect 3476 45512 199384 45540
rect 3476 45500 3482 45512
rect 199378 45500 199384 45512
rect 199436 45500 199442 45552
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 95878 33096 95884 33108
rect 3568 33068 95884 33096
rect 3568 33056 3574 33068
rect 95878 33056 95884 33068
rect 95936 33056 95942 33108
rect 577498 33056 577504 33108
rect 577556 33096 577562 33108
rect 579614 33096 579620 33108
rect 577556 33068 579620 33096
rect 577556 33056 577562 33068
rect 579614 33056 579620 33068
rect 579672 33056 579678 33108
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 64138 20652 64144 20664
rect 3476 20624 64144 20652
rect 3476 20612 3482 20624
rect 64138 20612 64144 20624
rect 64196 20612 64202 20664
rect 160094 11704 160100 11756
rect 160152 11744 160158 11756
rect 161290 11744 161296 11756
rect 160152 11716 161296 11744
rect 160152 11704 160158 11716
rect 161290 11704 161296 11716
rect 161348 11704 161354 11756
rect 176654 11704 176660 11756
rect 176712 11744 176718 11756
rect 177850 11744 177856 11756
rect 176712 11716 177856 11744
rect 176712 11704 176718 11716
rect 177850 11704 177856 11716
rect 177908 11704 177914 11756
rect 184934 11704 184940 11756
rect 184992 11744 184998 11756
rect 186130 11744 186136 11756
rect 184992 11716 186136 11744
rect 184992 11704 184998 11716
rect 186130 11704 186136 11716
rect 186188 11704 186194 11756
rect 234614 11704 234620 11756
rect 234672 11744 234678 11756
rect 235810 11744 235816 11756
rect 234672 11716 235816 11744
rect 234672 11704 234678 11716
rect 235810 11704 235816 11716
rect 235868 11704 235874 11756
rect 242894 11704 242900 11756
rect 242952 11744 242958 11756
rect 244090 11744 244096 11756
rect 242952 11716 244096 11744
rect 242952 11704 242958 11716
rect 244090 11704 244096 11716
rect 244148 11704 244154 11756
rect 316218 9256 316224 9308
rect 316276 9296 316282 9308
rect 363414 9296 363420 9308
rect 316276 9268 363420 9296
rect 316276 9256 316282 9268
rect 363414 9256 363420 9268
rect 363472 9256 363478 9308
rect 319714 9188 319720 9240
rect 319772 9228 319778 9240
rect 367186 9228 367192 9240
rect 319772 9200 367192 9228
rect 319772 9188 319778 9200
rect 367186 9188 367192 9200
rect 367244 9188 367250 9240
rect 312630 9120 312636 9172
rect 312688 9160 312694 9172
rect 360286 9160 360292 9172
rect 312688 9132 360292 9160
rect 312688 9120 312694 9132
rect 360286 9120 360292 9132
rect 360344 9120 360350 9172
rect 305546 9052 305552 9104
rect 305604 9092 305610 9104
rect 366082 9092 366088 9104
rect 305604 9064 366088 9092
rect 305604 9052 305610 9064
rect 366082 9052 366088 9064
rect 366140 9052 366146 9104
rect 303154 8984 303160 9036
rect 303212 9024 303218 9036
rect 364518 9024 364524 9036
rect 303212 8996 364524 9024
rect 303212 8984 303218 8996
rect 364518 8984 364524 8996
rect 364576 8984 364582 9036
rect 304350 8916 304356 8968
rect 304408 8956 304414 8968
rect 365990 8956 365996 8968
rect 304408 8928 365996 8956
rect 304408 8916 304414 8928
rect 365990 8916 365996 8928
rect 366048 8916 366054 8968
rect 330386 6808 330392 6860
rect 330444 6848 330450 6860
rect 363322 6848 363328 6860
rect 330444 6820 363328 6848
rect 330444 6808 330450 6820
rect 363322 6808 363328 6820
rect 363380 6808 363386 6860
rect 326798 6740 326804 6792
rect 326856 6780 326862 6792
rect 360194 6780 360200 6792
rect 326856 6752 360200 6780
rect 326856 6740 326862 6752
rect 360194 6740 360200 6752
rect 360252 6740 360258 6792
rect 315022 6672 315028 6724
rect 315080 6712 315086 6724
rect 361942 6712 361948 6724
rect 315080 6684 361948 6712
rect 315080 6672 315086 6684
rect 361942 6672 361948 6684
rect 362000 6672 362006 6724
rect 313826 6604 313832 6656
rect 313884 6644 313890 6656
rect 360930 6644 360936 6656
rect 313884 6616 360936 6644
rect 313884 6604 313890 6616
rect 360930 6604 360936 6616
rect 360988 6604 360994 6656
rect 318518 6536 318524 6588
rect 318576 6576 318582 6588
rect 365898 6576 365904 6588
rect 318576 6548 365904 6576
rect 318576 6536 318582 6548
rect 365898 6536 365904 6548
rect 365956 6536 365962 6588
rect 317322 6468 317328 6520
rect 317380 6508 317386 6520
rect 364794 6508 364800 6520
rect 317380 6480 364800 6508
rect 317380 6468 317386 6480
rect 364794 6468 364800 6480
rect 364852 6468 364858 6520
rect 311434 6400 311440 6452
rect 311492 6440 311498 6452
rect 359458 6440 359464 6452
rect 311492 6412 359464 6440
rect 311492 6400 311498 6412
rect 359458 6400 359464 6412
rect 359516 6400 359522 6452
rect 310238 6332 310244 6384
rect 310296 6372 310302 6384
rect 358170 6372 358176 6384
rect 310296 6344 358176 6372
rect 310296 6332 310302 6344
rect 358170 6332 358176 6344
rect 358228 6332 358234 6384
rect 307938 6264 307944 6316
rect 307996 6304 308002 6316
rect 369854 6304 369860 6316
rect 307996 6276 369860 6304
rect 307996 6264 308002 6276
rect 369854 6264 369860 6276
rect 369912 6264 369918 6316
rect 306742 6196 306748 6248
rect 306800 6236 306806 6248
rect 368474 6236 368480 6248
rect 306800 6208 368480 6236
rect 306800 6196 306806 6208
rect 368474 6196 368480 6208
rect 368532 6196 368538 6248
rect 309042 6128 309048 6180
rect 309100 6168 309106 6180
rect 372706 6168 372712 6180
rect 309100 6140 372712 6168
rect 309100 6128 309106 6140
rect 372706 6128 372712 6140
rect 372764 6128 372770 6180
rect 333882 6060 333888 6112
rect 333940 6100 333946 6112
rect 364702 6100 364708 6112
rect 333940 6072 364708 6100
rect 333940 6060 333946 6072
rect 364702 6060 364708 6072
rect 364760 6060 364766 6112
rect 337470 5992 337476 6044
rect 337528 6032 337534 6044
rect 363230 6032 363236 6044
rect 337528 6004 363236 6032
rect 337528 5992 337534 6004
rect 363230 5992 363236 6004
rect 363288 5992 363294 6044
rect 340966 5924 340972 5976
rect 341024 5964 341030 5976
rect 364610 5964 364616 5976
rect 341024 5936 364616 5964
rect 341024 5924 341030 5936
rect 364610 5924 364616 5936
rect 364668 5924 364674 5976
rect 180242 4088 180248 4140
rect 180300 4128 180306 4140
rect 181438 4128 181444 4140
rect 180300 4100 181444 4128
rect 180300 4088 180306 4100
rect 181438 4088 181444 4100
rect 181496 4088 181502 4140
rect 208578 4088 208584 4140
rect 208636 4128 208642 4140
rect 211798 4128 211804 4140
rect 208636 4100 211804 4128
rect 208636 4088 208642 4100
rect 211798 4088 211804 4100
rect 211856 4088 211862 4140
rect 212350 4088 212356 4140
rect 212408 4128 212414 4140
rect 245194 4128 245200 4140
rect 212408 4100 245200 4128
rect 212408 4088 212414 4100
rect 245194 4088 245200 4100
rect 245252 4088 245258 4140
rect 336274 4088 336280 4140
rect 336332 4128 336338 4140
rect 362954 4128 362960 4140
rect 336332 4100 362960 4128
rect 336332 4088 336338 4100
rect 362954 4088 362960 4100
rect 363012 4088 363018 4140
rect 460198 4088 460204 4140
rect 460256 4128 460262 4140
rect 462774 4128 462780 4140
rect 460256 4100 462780 4128
rect 460256 4088 460262 4100
rect 462774 4088 462780 4100
rect 462832 4088 462838 4140
rect 468478 4088 468484 4140
rect 468536 4128 468542 4140
rect 471054 4128 471060 4140
rect 468536 4100 471060 4128
rect 468536 4088 468542 4100
rect 471054 4088 471060 4100
rect 471112 4088 471118 4140
rect 51350 4020 51356 4072
rect 51408 4060 51414 4072
rect 57238 4060 57244 4072
rect 51408 4032 57244 4060
rect 51408 4020 51414 4032
rect 57238 4020 57244 4032
rect 57296 4020 57302 4072
rect 213822 4020 213828 4072
rect 213880 4060 213886 4072
rect 258258 4060 258264 4072
rect 213880 4032 258264 4060
rect 213880 4020 213886 4032
rect 258258 4020 258264 4032
rect 258316 4020 258322 4072
rect 332686 4020 332692 4072
rect 332744 4060 332750 4072
rect 364334 4060 364340 4072
rect 332744 4032 364340 4060
rect 332744 4020 332750 4032
rect 364334 4020 364340 4032
rect 364392 4020 364398 4072
rect 213730 3952 213736 4004
rect 213788 3992 213794 4004
rect 260650 3992 260656 4004
rect 213788 3964 260656 3992
rect 213788 3952 213794 3964
rect 260650 3952 260656 3964
rect 260708 3952 260714 4004
rect 329190 3952 329196 4004
rect 329248 3992 329254 4004
rect 363046 3992 363052 4004
rect 329248 3964 363052 3992
rect 329248 3952 329254 3964
rect 363046 3952 363052 3964
rect 363104 3952 363110 4004
rect 219342 3884 219348 3936
rect 219400 3924 219406 3936
rect 266538 3924 266544 3936
rect 219400 3896 266544 3924
rect 219400 3884 219406 3896
rect 266538 3884 266544 3896
rect 266596 3884 266602 3936
rect 322106 3884 322112 3936
rect 322164 3924 322170 3936
rect 356698 3924 356704 3936
rect 322164 3896 356704 3924
rect 322164 3884 322170 3896
rect 356698 3884 356704 3896
rect 356756 3884 356762 3936
rect 371878 3884 371884 3936
rect 371936 3924 371942 3936
rect 375282 3924 375288 3936
rect 371936 3896 375288 3924
rect 371936 3884 371942 3896
rect 375282 3884 375288 3896
rect 375340 3884 375346 3936
rect 4062 3816 4068 3868
rect 4120 3856 4126 3868
rect 7558 3856 7564 3868
rect 4120 3828 7564 3856
rect 4120 3816 4126 3828
rect 7558 3816 7564 3828
rect 7616 3816 7622 3868
rect 214926 3816 214932 3868
rect 214984 3856 214990 3868
rect 262950 3856 262956 3868
rect 214984 3828 262956 3856
rect 214984 3816 214990 3828
rect 262950 3816 262956 3828
rect 263008 3816 263014 3868
rect 298462 3816 298468 3868
rect 298520 3856 298526 3868
rect 345750 3856 345756 3868
rect 298520 3828 345756 3856
rect 298520 3816 298526 3828
rect 345750 3816 345756 3828
rect 345808 3816 345814 3868
rect 516778 3816 516784 3868
rect 516836 3856 516842 3868
rect 519538 3856 519544 3868
rect 516836 3828 519544 3856
rect 516836 3816 516842 3828
rect 519538 3816 519544 3828
rect 519596 3816 519602 3868
rect 566458 3816 566464 3868
rect 566516 3856 566522 3868
rect 569126 3856 569132 3868
rect 566516 3828 569132 3856
rect 566516 3816 566522 3828
rect 569126 3816 569132 3828
rect 569184 3816 569190 3868
rect 69106 3748 69112 3800
rect 69164 3788 69170 3800
rect 71038 3788 71044 3800
rect 69164 3760 71044 3788
rect 69164 3748 69170 3760
rect 71038 3748 71044 3760
rect 71096 3748 71102 3800
rect 135254 3748 135260 3800
rect 135312 3788 135318 3800
rect 136450 3788 136456 3800
rect 135312 3760 136456 3788
rect 135312 3748 135318 3760
rect 136450 3748 136456 3760
rect 136508 3748 136514 3800
rect 195974 3748 195980 3800
rect 196032 3788 196038 3800
rect 196618 3788 196624 3800
rect 196032 3760 196624 3788
rect 196032 3748 196038 3760
rect 196618 3748 196624 3760
rect 196676 3748 196682 3800
rect 218698 3748 218704 3800
rect 218756 3788 218762 3800
rect 277118 3788 277124 3800
rect 218756 3760 277124 3788
rect 218756 3748 218762 3760
rect 277118 3748 277124 3760
rect 277176 3748 277182 3800
rect 300762 3748 300768 3800
rect 300820 3788 300826 3800
rect 354122 3788 354128 3800
rect 300820 3760 354128 3788
rect 300820 3748 300826 3760
rect 354122 3748 354128 3760
rect 354180 3748 354186 3800
rect 355134 3748 355140 3800
rect 355192 3788 355198 3800
rect 361574 3788 361580 3800
rect 355192 3760 361580 3788
rect 355192 3748 355198 3760
rect 361574 3748 361580 3760
rect 361632 3748 361638 3800
rect 30098 3680 30104 3732
rect 30156 3720 30162 3732
rect 39390 3720 39396 3732
rect 30156 3692 39396 3720
rect 30156 3680 30162 3692
rect 39390 3680 39396 3692
rect 39448 3680 39454 3732
rect 44266 3680 44272 3732
rect 44324 3720 44330 3732
rect 46198 3720 46204 3732
rect 44324 3692 46204 3720
rect 44324 3680 44330 3692
rect 46198 3680 46204 3692
rect 46256 3680 46262 3732
rect 46658 3680 46664 3732
rect 46716 3720 46722 3732
rect 170490 3720 170496 3732
rect 46716 3692 170496 3720
rect 46716 3680 46722 3692
rect 170490 3680 170496 3692
rect 170548 3680 170554 3732
rect 211062 3680 211068 3732
rect 211120 3720 211126 3732
rect 268838 3720 268844 3732
rect 211120 3692 268844 3720
rect 211120 3680 211126 3692
rect 268838 3680 268844 3692
rect 268896 3680 268902 3732
rect 292574 3680 292580 3732
rect 292632 3720 292638 3732
rect 348418 3720 348424 3732
rect 292632 3692 348424 3720
rect 292632 3680 292638 3692
rect 348418 3680 348424 3692
rect 348476 3680 348482 3732
rect 352834 3680 352840 3732
rect 352892 3720 352898 3732
rect 361022 3720 361028 3732
rect 352892 3692 361028 3720
rect 352892 3680 352898 3692
rect 361022 3680 361028 3692
rect 361080 3680 361086 3732
rect 489178 3680 489184 3732
rect 489236 3720 489242 3732
rect 491110 3720 491116 3732
rect 489236 3692 491116 3720
rect 489236 3680 489242 3692
rect 491110 3680 491116 3692
rect 491168 3680 491174 3732
rect 6454 3612 6460 3664
rect 6512 3652 6518 3664
rect 18598 3652 18604 3664
rect 6512 3624 18604 3652
rect 6512 3612 6518 3624
rect 18598 3612 18604 3624
rect 18656 3612 18662 3664
rect 25314 3612 25320 3664
rect 25372 3652 25378 3664
rect 171778 3652 171784 3664
rect 25372 3624 171784 3652
rect 25372 3612 25378 3624
rect 171778 3612 171784 3624
rect 171836 3612 171842 3664
rect 183738 3612 183744 3664
rect 183796 3652 183802 3664
rect 188338 3652 188344 3664
rect 183796 3624 188344 3652
rect 183796 3612 183802 3624
rect 188338 3612 188344 3624
rect 188396 3612 188402 3664
rect 209774 3612 209780 3664
rect 209832 3652 209838 3664
rect 210970 3652 210976 3664
rect 209832 3624 210976 3652
rect 209832 3612 209838 3624
rect 210970 3612 210976 3624
rect 211028 3612 211034 3664
rect 217318 3612 217324 3664
rect 217376 3652 217382 3664
rect 276014 3652 276020 3664
rect 217376 3624 276020 3652
rect 217376 3612 217382 3624
rect 276014 3612 276020 3624
rect 276072 3612 276078 3664
rect 290182 3612 290188 3664
rect 290240 3652 290246 3664
rect 351178 3652 351184 3664
rect 290240 3624 351184 3652
rect 290240 3612 290246 3624
rect 351178 3612 351184 3624
rect 351236 3612 351242 3664
rect 354030 3612 354036 3664
rect 354088 3652 354094 3664
rect 365254 3652 365260 3664
rect 354088 3624 365260 3652
rect 354088 3612 354094 3624
rect 365254 3612 365260 3624
rect 365312 3612 365318 3664
rect 371326 3652 371332 3664
rect 367848 3624 371332 3652
rect 1670 3544 1676 3596
rect 1728 3584 1734 3596
rect 32398 3584 32404 3596
rect 1728 3556 32404 3584
rect 1728 3544 1734 3556
rect 32398 3544 32404 3556
rect 32456 3544 32462 3596
rect 33594 3544 33600 3596
rect 33652 3584 33658 3596
rect 35158 3584 35164 3596
rect 33652 3556 35164 3584
rect 33652 3544 33658 3556
rect 35158 3544 35164 3556
rect 35216 3544 35222 3596
rect 38378 3544 38384 3596
rect 38436 3584 38442 3596
rect 39298 3584 39304 3596
rect 38436 3556 39304 3584
rect 38436 3544 38442 3556
rect 39298 3544 39304 3556
rect 39356 3544 39362 3596
rect 52454 3544 52460 3596
rect 52512 3584 52518 3596
rect 53374 3584 53380 3596
rect 52512 3556 53380 3584
rect 52512 3544 52518 3556
rect 53374 3544 53380 3556
rect 53432 3544 53438 3596
rect 56042 3544 56048 3596
rect 56100 3584 56106 3596
rect 57330 3584 57336 3596
rect 56100 3556 57336 3584
rect 56100 3544 56106 3556
rect 57330 3544 57336 3556
rect 57388 3544 57394 3596
rect 59630 3544 59636 3596
rect 59688 3584 59694 3596
rect 211890 3584 211896 3596
rect 59688 3556 211896 3584
rect 59688 3544 59694 3556
rect 211890 3544 211896 3556
rect 211948 3544 211954 3596
rect 212442 3544 212448 3596
rect 212500 3584 212506 3596
rect 272426 3584 272432 3596
rect 212500 3556 272432 3584
rect 212500 3544 212506 3556
rect 272426 3544 272432 3556
rect 272484 3544 272490 3596
rect 285398 3544 285404 3596
rect 285456 3584 285462 3596
rect 345658 3584 345664 3596
rect 285456 3556 345664 3584
rect 285456 3544 285462 3556
rect 345658 3544 345664 3556
rect 345716 3544 345722 3596
rect 349246 3544 349252 3596
rect 349304 3584 349310 3596
rect 355134 3584 355140 3596
rect 349304 3556 355140 3584
rect 349304 3544 349310 3556
rect 355134 3544 355140 3556
rect 355192 3544 355198 3596
rect 355226 3544 355232 3596
rect 355284 3584 355290 3596
rect 355284 3556 358216 3584
rect 355284 3544 355290 3556
rect 12342 3476 12348 3528
rect 12400 3516 12406 3528
rect 13078 3516 13084 3528
rect 12400 3488 13084 3516
rect 12400 3476 12406 3488
rect 13078 3476 13084 3488
rect 13136 3476 13142 3528
rect 15930 3476 15936 3528
rect 15988 3516 15994 3528
rect 170398 3516 170404 3528
rect 15988 3488 170404 3516
rect 15988 3476 15994 3488
rect 170398 3476 170404 3488
rect 170456 3476 170462 3528
rect 187326 3476 187332 3528
rect 187384 3516 187390 3528
rect 195974 3516 195980 3528
rect 187384 3488 195980 3516
rect 187384 3476 187390 3488
rect 195974 3476 195980 3488
rect 196032 3476 196038 3528
rect 209682 3476 209688 3528
rect 209740 3516 209746 3528
rect 218054 3516 218060 3528
rect 209740 3488 218060 3516
rect 209740 3476 209746 3488
rect 218054 3476 218060 3488
rect 218112 3476 218118 3528
rect 219158 3476 219164 3528
rect 219216 3516 219222 3528
rect 280706 3516 280712 3528
rect 219216 3488 280712 3516
rect 219216 3476 219222 3488
rect 280706 3476 280712 3488
rect 280764 3476 280770 3528
rect 281902 3476 281908 3528
rect 281960 3516 281966 3528
rect 353938 3516 353944 3528
rect 281960 3488 353944 3516
rect 281960 3476 281966 3488
rect 353938 3476 353944 3488
rect 353996 3476 354002 3528
rect 356330 3476 356336 3528
rect 356388 3516 356394 3528
rect 358078 3516 358084 3528
rect 356388 3488 358084 3516
rect 356388 3476 356394 3488
rect 358078 3476 358084 3488
rect 358136 3476 358142 3528
rect 358188 3516 358216 3556
rect 362310 3544 362316 3596
rect 362368 3584 362374 3596
rect 367848 3584 367876 3624
rect 371326 3612 371332 3624
rect 371384 3612 371390 3664
rect 377398 3612 377404 3664
rect 377456 3652 377462 3664
rect 411898 3652 411904 3664
rect 377456 3624 411904 3652
rect 377456 3612 377462 3624
rect 411898 3612 411904 3624
rect 411956 3612 411962 3664
rect 362368 3556 367876 3584
rect 362368 3544 362374 3556
rect 369394 3544 369400 3596
rect 369452 3584 369458 3596
rect 372798 3584 372804 3596
rect 369452 3556 372804 3584
rect 369452 3544 369458 3556
rect 372798 3544 372804 3556
rect 372856 3544 372862 3596
rect 381538 3544 381544 3596
rect 381596 3584 381602 3596
rect 384758 3584 384764 3596
rect 381596 3556 384764 3584
rect 381596 3544 381602 3556
rect 384758 3544 384764 3556
rect 384816 3544 384822 3596
rect 398834 3544 398840 3596
rect 398892 3584 398898 3596
rect 400122 3584 400128 3596
rect 398892 3556 400128 3584
rect 398892 3544 398898 3556
rect 400122 3544 400128 3556
rect 400180 3544 400186 3596
rect 407206 3544 407212 3596
rect 407264 3584 407270 3596
rect 408402 3584 408408 3596
rect 407264 3556 408408 3584
rect 407264 3544 407270 3556
rect 408402 3544 408408 3556
rect 408460 3544 408466 3596
rect 421558 3544 421564 3596
rect 421616 3584 421622 3596
rect 427262 3584 427268 3596
rect 421616 3556 427268 3584
rect 421616 3544 421622 3556
rect 427262 3544 427268 3556
rect 427320 3544 427326 3596
rect 442258 3544 442264 3596
rect 442316 3584 442322 3596
rect 445018 3584 445024 3596
rect 442316 3556 445024 3584
rect 442316 3544 442322 3556
rect 445018 3544 445024 3556
rect 445076 3544 445082 3596
rect 445110 3544 445116 3596
rect 445168 3584 445174 3596
rect 458082 3584 458088 3596
rect 445168 3556 458088 3584
rect 445168 3544 445174 3556
rect 458082 3544 458088 3556
rect 458140 3544 458146 3596
rect 458818 3544 458824 3596
rect 458876 3584 458882 3596
rect 465166 3584 465172 3596
rect 458876 3556 465172 3584
rect 458876 3544 458882 3556
rect 465166 3544 465172 3556
rect 465224 3544 465230 3596
rect 467098 3544 467104 3596
rect 467156 3584 467162 3596
rect 469858 3584 469864 3596
rect 467156 3556 469864 3584
rect 467156 3544 467162 3556
rect 469858 3544 469864 3556
rect 469916 3544 469922 3596
rect 470566 3556 475240 3584
rect 365714 3516 365720 3528
rect 358188 3488 365720 3516
rect 365714 3476 365720 3488
rect 365772 3476 365778 3528
rect 381630 3476 381636 3528
rect 381688 3516 381694 3528
rect 381688 3488 423628 3516
rect 381688 3476 381694 3488
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 171134 3448 171140 3460
rect 624 3420 171140 3448
rect 624 3408 630 3420
rect 171134 3408 171140 3420
rect 171192 3408 171198 3460
rect 190822 3408 190828 3460
rect 190880 3448 190886 3460
rect 203518 3448 203524 3460
rect 190880 3420 203524 3448
rect 190880 3408 190886 3420
rect 203518 3408 203524 3420
rect 203576 3408 203582 3460
rect 216582 3408 216588 3460
rect 216640 3448 216646 3460
rect 284294 3448 284300 3460
rect 216640 3420 284300 3448
rect 216640 3408 216646 3420
rect 284294 3408 284300 3420
rect 284352 3408 284358 3460
rect 286594 3408 286600 3460
rect 286652 3448 286658 3460
rect 367094 3448 367100 3460
rect 286652 3420 367100 3448
rect 286652 3408 286658 3420
rect 367094 3408 367100 3420
rect 367152 3408 367158 3460
rect 382366 3408 382372 3460
rect 382424 3448 382430 3460
rect 383562 3448 383568 3460
rect 382424 3420 383568 3448
rect 382424 3408 382430 3420
rect 383562 3408 383568 3420
rect 383620 3408 383626 3460
rect 387058 3408 387064 3460
rect 387116 3448 387122 3460
rect 388254 3448 388260 3460
rect 387116 3420 388260 3448
rect 387116 3408 387122 3420
rect 388254 3408 388260 3420
rect 388312 3408 388318 3460
rect 390554 3408 390560 3460
rect 390612 3448 390618 3460
rect 391842 3448 391848 3460
rect 390612 3420 391848 3448
rect 390612 3408 390618 3420
rect 391842 3408 391848 3420
rect 391900 3408 391906 3460
rect 393286 3420 412634 3448
rect 37182 3340 37188 3392
rect 37240 3380 37246 3392
rect 43438 3380 43444 3392
rect 37240 3352 43444 3380
rect 37240 3340 37246 3352
rect 43438 3340 43444 3352
rect 43496 3340 43502 3392
rect 57238 3340 57244 3392
rect 57296 3380 57302 3392
rect 58618 3380 58624 3392
rect 57296 3352 58624 3380
rect 57296 3340 57302 3352
rect 58618 3340 58624 3352
rect 58676 3340 58682 3392
rect 118694 3340 118700 3392
rect 118752 3380 118758 3392
rect 119890 3380 119896 3392
rect 118752 3352 119896 3380
rect 118752 3340 118758 3352
rect 119890 3340 119896 3352
rect 119948 3340 119954 3392
rect 215018 3340 215024 3392
rect 215076 3380 215082 3392
rect 240502 3380 240508 3392
rect 215076 3352 240508 3380
rect 215076 3340 215082 3352
rect 240502 3340 240508 3352
rect 240560 3340 240566 3392
rect 339862 3340 339868 3392
rect 339920 3380 339926 3392
rect 364426 3380 364432 3392
rect 339920 3352 364432 3380
rect 339920 3340 339926 3352
rect 364426 3340 364432 3352
rect 364484 3340 364490 3392
rect 388438 3340 388444 3392
rect 388496 3380 388502 3392
rect 393286 3380 393314 3420
rect 388496 3352 393314 3380
rect 388496 3340 388502 3352
rect 215110 3272 215116 3324
rect 215168 3312 215174 3324
rect 226334 3312 226340 3324
rect 215168 3284 226340 3312
rect 215168 3272 215174 3284
rect 226334 3272 226340 3284
rect 226392 3272 226398 3324
rect 338666 3272 338672 3324
rect 338724 3312 338730 3324
rect 361666 3312 361672 3324
rect 338724 3284 361672 3312
rect 338724 3272 338730 3284
rect 361666 3272 361672 3284
rect 361724 3272 361730 3324
rect 412606 3312 412634 3420
rect 414658 3408 414664 3460
rect 414716 3448 414722 3460
rect 416682 3448 416688 3460
rect 414716 3420 416688 3448
rect 414716 3408 414722 3420
rect 416682 3408 416688 3420
rect 416740 3408 416746 3460
rect 423600 3380 423628 3488
rect 423766 3476 423772 3528
rect 423824 3516 423830 3528
rect 424962 3516 424968 3528
rect 423824 3488 424968 3516
rect 423824 3476 423830 3488
rect 424962 3476 424968 3488
rect 425020 3476 425026 3528
rect 429654 3516 429660 3528
rect 425072 3488 429660 3516
rect 425072 3380 425100 3488
rect 429654 3476 429660 3488
rect 429712 3476 429718 3528
rect 431954 3476 431960 3528
rect 432012 3516 432018 3528
rect 433242 3516 433248 3528
rect 432012 3488 433248 3516
rect 432012 3476 432018 3488
rect 433242 3476 433248 3488
rect 433300 3476 433306 3528
rect 440326 3476 440332 3528
rect 440384 3516 440390 3528
rect 441522 3516 441528 3528
rect 440384 3488 441528 3516
rect 440384 3476 440390 3488
rect 441522 3476 441528 3488
rect 441580 3476 441586 3528
rect 443638 3476 443644 3528
rect 443696 3516 443702 3528
rect 447410 3516 447416 3528
rect 443696 3488 447416 3516
rect 443696 3476 443702 3488
rect 447410 3476 447416 3488
rect 447468 3476 447474 3528
rect 448514 3476 448520 3528
rect 448572 3516 448578 3528
rect 449802 3516 449808 3528
rect 448572 3488 449808 3516
rect 448572 3476 448578 3488
rect 449802 3476 449808 3488
rect 449860 3476 449866 3528
rect 454678 3476 454684 3528
rect 454736 3516 454742 3528
rect 456886 3516 456892 3528
rect 454736 3488 456892 3516
rect 454736 3476 454742 3488
rect 456886 3476 456892 3488
rect 456944 3476 456950 3528
rect 462958 3476 462964 3528
rect 463016 3516 463022 3528
rect 470566 3516 470594 3556
rect 463016 3488 470594 3516
rect 463016 3476 463022 3488
rect 471238 3476 471244 3528
rect 471296 3516 471302 3528
rect 473446 3516 473452 3528
rect 471296 3488 473452 3516
rect 471296 3476 471302 3488
rect 473446 3476 473452 3488
rect 473504 3476 473510 3528
rect 475212 3516 475240 3556
rect 475378 3544 475384 3596
rect 475436 3584 475442 3596
rect 476942 3584 476948 3596
rect 475436 3556 476948 3584
rect 475436 3544 475442 3556
rect 476942 3544 476948 3556
rect 477000 3544 477006 3596
rect 500218 3544 500224 3596
rect 500276 3584 500282 3596
rect 501782 3584 501788 3596
rect 500276 3556 501788 3584
rect 500276 3544 500282 3556
rect 501782 3544 501788 3556
rect 501840 3544 501846 3596
rect 511258 3544 511264 3596
rect 511316 3584 511322 3596
rect 513558 3584 513564 3596
rect 511316 3556 513564 3584
rect 511316 3544 511322 3556
rect 513558 3544 513564 3556
rect 513616 3544 513622 3596
rect 518158 3544 518164 3596
rect 518216 3584 518222 3596
rect 521838 3584 521844 3596
rect 518216 3556 521844 3584
rect 518216 3544 518222 3556
rect 521838 3544 521844 3556
rect 521896 3544 521902 3596
rect 525058 3544 525064 3596
rect 525116 3584 525122 3596
rect 527726 3584 527732 3596
rect 525116 3556 527732 3584
rect 525116 3544 525122 3556
rect 527726 3544 527732 3556
rect 527784 3544 527790 3596
rect 533706 3584 533712 3596
rect 528526 3556 533712 3584
rect 479334 3516 479340 3528
rect 475212 3488 479340 3516
rect 479334 3476 479340 3488
rect 479392 3476 479398 3528
rect 481634 3476 481640 3528
rect 481692 3516 481698 3528
rect 482462 3516 482468 3528
rect 481692 3488 482468 3516
rect 481692 3476 481698 3488
rect 482462 3476 482468 3488
rect 482520 3476 482526 3528
rect 496078 3476 496084 3528
rect 496136 3516 496142 3528
rect 497090 3516 497096 3528
rect 496136 3488 497096 3516
rect 496136 3476 496142 3488
rect 497090 3476 497096 3488
rect 497148 3476 497154 3528
rect 506474 3476 506480 3528
rect 506532 3516 506538 3528
rect 507302 3516 507308 3528
rect 506532 3488 507308 3516
rect 506532 3476 506538 3488
rect 507302 3476 507308 3488
rect 507360 3476 507366 3528
rect 520918 3476 520924 3528
rect 520976 3516 520982 3528
rect 523034 3516 523040 3528
rect 520976 3488 523040 3516
rect 520976 3476 520982 3488
rect 523034 3476 523040 3488
rect 523092 3476 523098 3528
rect 527818 3476 527824 3528
rect 527876 3516 527882 3528
rect 528526 3516 528554 3556
rect 533706 3544 533712 3556
rect 533764 3544 533770 3596
rect 549898 3544 549904 3596
rect 549956 3584 549962 3596
rect 551462 3584 551468 3596
rect 549956 3556 551468 3584
rect 549956 3544 549962 3556
rect 551462 3544 551468 3556
rect 551520 3544 551526 3596
rect 567838 3544 567844 3596
rect 567896 3584 567902 3596
rect 571518 3584 571524 3596
rect 567896 3556 571524 3584
rect 567896 3544 567902 3556
rect 571518 3544 571524 3556
rect 571576 3544 571582 3596
rect 527876 3488 528554 3516
rect 527876 3476 527882 3488
rect 531314 3476 531320 3528
rect 531372 3516 531378 3528
rect 532142 3516 532148 3528
rect 531372 3488 532148 3516
rect 531372 3476 531378 3488
rect 532142 3476 532148 3488
rect 532200 3476 532206 3528
rect 545758 3476 545764 3528
rect 545816 3516 545822 3528
rect 546678 3516 546684 3528
rect 545816 3488 546684 3516
rect 545816 3476 545822 3488
rect 546678 3476 546684 3488
rect 546736 3476 546742 3528
rect 556154 3476 556160 3528
rect 556212 3516 556218 3528
rect 556982 3516 556988 3528
rect 556212 3488 556988 3516
rect 556212 3476 556218 3488
rect 556982 3476 556988 3488
rect 557040 3476 557046 3528
rect 570598 3476 570604 3528
rect 570656 3516 570662 3528
rect 572714 3516 572720 3528
rect 570656 3488 572720 3516
rect 570656 3476 570662 3488
rect 572714 3476 572720 3488
rect 572772 3476 572778 3528
rect 580994 3448 581000 3460
rect 423600 3352 425100 3380
rect 425164 3420 581000 3448
rect 425164 3312 425192 3420
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 493318 3340 493324 3392
rect 493376 3380 493382 3392
rect 499390 3380 499396 3392
rect 493376 3352 499396 3380
rect 493376 3340 493382 3352
rect 499390 3340 499396 3352
rect 499448 3340 499454 3392
rect 542998 3340 543004 3392
rect 543056 3380 543062 3392
rect 549070 3380 549076 3392
rect 543056 3352 549076 3380
rect 543056 3340 543062 3352
rect 549070 3340 549076 3352
rect 549128 3340 549134 3392
rect 412606 3284 425192 3312
rect 428550 3272 428556 3324
rect 428608 3312 428614 3324
rect 434438 3312 434444 3324
rect 428608 3284 434444 3312
rect 428608 3272 428614 3284
rect 434438 3272 434444 3284
rect 434496 3272 434502 3324
rect 509878 3272 509884 3324
rect 509936 3312 509942 3324
rect 514754 3312 514760 3324
rect 509936 3284 514760 3312
rect 509936 3272 509942 3284
rect 514754 3272 514760 3284
rect 514812 3272 514818 3324
rect 342162 3204 342168 3256
rect 342220 3244 342226 3256
rect 361758 3244 361764 3256
rect 342220 3216 361764 3244
rect 342220 3204 342226 3216
rect 361758 3204 361764 3216
rect 361816 3204 361822 3256
rect 446398 3204 446404 3256
rect 446456 3244 446462 3256
rect 452102 3244 452108 3256
rect 446456 3216 452108 3244
rect 446456 3204 446462 3216
rect 452102 3204 452108 3216
rect 452160 3204 452166 3256
rect 216490 3136 216496 3188
rect 216548 3176 216554 3188
rect 227530 3176 227536 3188
rect 216548 3148 227536 3176
rect 216548 3136 216554 3148
rect 227530 3136 227536 3148
rect 227588 3136 227594 3188
rect 345750 3136 345756 3188
rect 345808 3176 345814 3188
rect 361850 3176 361856 3188
rect 345808 3148 361856 3176
rect 345808 3136 345814 3148
rect 361850 3136 361856 3148
rect 361908 3136 361914 3188
rect 485038 3136 485044 3188
rect 485096 3176 485102 3188
rect 487614 3176 487620 3188
rect 485096 3148 487620 3176
rect 485096 3136 485102 3148
rect 487614 3136 487620 3148
rect 487672 3136 487678 3188
rect 534718 3136 534724 3188
rect 534776 3176 534782 3188
rect 537202 3176 537208 3188
rect 534776 3148 537208 3176
rect 534776 3136 534782 3148
rect 537202 3136 537208 3148
rect 537260 3136 537266 3188
rect 560938 3136 560944 3188
rect 560996 3176 561002 3188
rect 563238 3176 563244 3188
rect 560996 3148 563244 3176
rect 560996 3136 561002 3148
rect 563238 3136 563244 3148
rect 563296 3136 563302 3188
rect 19426 3000 19432 3052
rect 19484 3040 19490 3052
rect 25590 3040 25596 3052
rect 19484 3012 25596 3040
rect 19484 3000 19490 3012
rect 25590 3000 25596 3012
rect 25648 3000 25654 3052
rect 195606 3000 195612 3052
rect 195664 3040 195670 3052
rect 198090 3040 198096 3052
rect 195664 3012 198096 3040
rect 195664 3000 195670 3012
rect 198090 3000 198096 3012
rect 198148 3000 198154 3052
rect 374638 3000 374644 3052
rect 374696 3040 374702 3052
rect 376478 3040 376484 3052
rect 374696 3012 376484 3040
rect 374696 3000 374702 3012
rect 376478 3000 376484 3012
rect 376536 3000 376542 3052
rect 413278 3000 413284 3052
rect 413336 3040 413342 3052
rect 415486 3040 415492 3052
rect 413336 3012 415492 3040
rect 413336 3000 413342 3012
rect 415486 3000 415492 3012
rect 415544 3000 415550 3052
rect 417510 3000 417516 3052
rect 417568 3040 417574 3052
rect 420178 3040 420184 3052
rect 417568 3012 420184 3040
rect 417568 3000 417574 3012
rect 420178 3000 420184 3012
rect 420236 3000 420242 3052
rect 464338 3000 464344 3052
rect 464396 3040 464402 3052
rect 466270 3040 466276 3052
rect 464396 3012 466276 3040
rect 464396 3000 464402 3012
rect 466270 3000 466276 3012
rect 466328 3000 466334 3052
rect 486510 3000 486516 3052
rect 486568 3040 486574 3052
rect 488810 3040 488816 3052
rect 486568 3012 488816 3040
rect 486568 3000 486574 3012
rect 488810 3000 488816 3012
rect 488868 3000 488874 3052
rect 514018 3000 514024 3052
rect 514076 3040 514082 3052
rect 515950 3040 515956 3052
rect 514076 3012 515956 3040
rect 514076 3000 514082 3012
rect 515950 3000 515956 3012
rect 516008 3000 516014 3052
rect 522298 3000 522304 3052
rect 522356 3040 522362 3052
rect 524230 3040 524236 3052
rect 522356 3012 524236 3040
rect 522356 3000 522362 3012
rect 524230 3000 524236 3012
rect 524288 3000 524294 3052
rect 538858 3000 538864 3052
rect 538916 3040 538922 3052
rect 540790 3040 540796 3052
rect 538916 3012 540796 3040
rect 538916 3000 538922 3012
rect 540790 3000 540796 3012
rect 540848 3000 540854 3052
rect 563698 3000 563704 3052
rect 563756 3040 563762 3052
rect 565630 3040 565636 3052
rect 563756 3012 565636 3040
rect 563756 3000 563762 3012
rect 565630 3000 565636 3012
rect 565688 3000 565694 3052
rect 571978 3000 571984 3052
rect 572036 3040 572042 3052
rect 573910 3040 573916 3052
rect 572036 3012 573916 3040
rect 572036 3000 572042 3012
rect 573910 3000 573916 3012
rect 573968 3000 573974 3052
rect 378778 2932 378784 2984
rect 378836 2972 378842 2984
rect 381170 2972 381176 2984
rect 378836 2944 381176 2972
rect 378836 2932 378842 2944
rect 381170 2932 381176 2944
rect 381228 2932 381234 2984
rect 396718 2932 396724 2984
rect 396776 2972 396782 2984
rect 402514 2972 402520 2984
rect 396776 2944 402520 2972
rect 396776 2932 396782 2944
rect 402514 2932 402520 2944
rect 402572 2932 402578 2984
rect 457438 2932 457444 2984
rect 457496 2972 457502 2984
rect 459186 2972 459192 2984
rect 457496 2944 459192 2972
rect 457496 2932 457502 2944
rect 459186 2932 459192 2944
rect 459244 2932 459250 2984
rect 552750 2932 552756 2984
rect 552808 2972 552814 2984
rect 554958 2972 554964 2984
rect 552808 2944 554964 2972
rect 552808 2932 552814 2944
rect 554958 2932 554964 2944
rect 555016 2932 555022 2984
rect 13538 2864 13544 2916
rect 13596 2904 13602 2916
rect 14458 2904 14464 2916
rect 13596 2876 14464 2904
rect 13596 2864 13602 2876
rect 14458 2864 14464 2876
rect 14516 2864 14522 2916
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 219348 700408 219400 700460
rect 267648 700408 267700 700460
rect 137836 700340 137888 700392
rect 138664 700340 138716 700392
rect 217968 700340 218020 700392
rect 283840 700340 283892 700392
rect 348792 700340 348844 700392
rect 358820 700340 358872 700392
rect 24308 700272 24360 700324
rect 215944 700272 215996 700324
rect 217876 700272 217928 700324
rect 300124 700272 300176 700324
rect 332508 700272 332560 700324
rect 357440 700272 357492 700324
rect 359464 700272 359516 700324
rect 429844 700272 429896 700324
rect 442264 700272 442316 700324
rect 559656 700272 559708 700324
rect 105452 699728 105504 699780
rect 108304 699728 108356 699780
rect 8116 699660 8168 699712
rect 10324 699660 10376 699712
rect 396724 699660 396776 699712
rect 397460 699660 397512 699712
rect 391204 696940 391256 696992
rect 580172 696940 580224 696992
rect 3424 683136 3476 683188
rect 21364 683136 21416 683188
rect 378784 683136 378836 683188
rect 580172 683136 580224 683188
rect 3516 670692 3568 670744
rect 214564 670692 214616 670744
rect 377404 670692 377456 670744
rect 580172 670692 580224 670744
rect 3424 656888 3476 656940
rect 28264 656888 28316 656940
rect 373264 643084 373316 643136
rect 580172 643084 580224 643136
rect 2780 632068 2832 632120
rect 4804 632068 4856 632120
rect 3148 618264 3200 618316
rect 211804 618264 211856 618316
rect 363604 616836 363656 616888
rect 580172 616836 580224 616888
rect 3424 606024 3476 606076
rect 7564 606024 7616 606076
rect 374644 590656 374696 590708
rect 580172 590656 580224 590708
rect 3332 579640 3384 579692
rect 57244 579640 57296 579692
rect 3424 565836 3476 565888
rect 210424 565836 210476 565888
rect 217784 565088 217836 565140
rect 234620 565088 234672 565140
rect 360844 563048 360896 563100
rect 579896 563048 579948 563100
rect 3424 553664 3476 553716
rect 8944 553664 8996 553716
rect 369124 536800 369176 536852
rect 580172 536800 580224 536852
rect 3424 527144 3476 527196
rect 35164 527144 35216 527196
rect 371884 524424 371936 524476
rect 580172 524424 580224 524476
rect 3424 514768 3476 514820
rect 207664 514768 207716 514820
rect 358084 510620 358136 510672
rect 580172 510620 580224 510672
rect 3056 500964 3108 501016
rect 13084 500964 13136 501016
rect 367744 484372 367796 484424
rect 580172 484372 580224 484424
rect 217876 478592 217928 478644
rect 269948 478592 270000 478644
rect 217968 478524 218020 478576
rect 271236 478524 271288 478576
rect 268660 478456 268712 478508
rect 357440 478456 357492 478508
rect 269304 478388 269356 478440
rect 358820 478388 358872 478440
rect 217416 478320 217468 478372
rect 308588 478320 308640 478372
rect 218980 478252 219032 478304
rect 314476 478252 314528 478304
rect 256884 478184 256936 478236
rect 374644 478184 374696 478236
rect 7564 478116 7616 478168
rect 282368 478116 282420 478168
rect 241428 476824 241480 476876
rect 238484 476756 238536 476808
rect 237288 476688 237340 476740
rect 239404 476688 239456 476740
rect 316408 476756 316460 476808
rect 311256 476688 311308 476740
rect 242808 476620 242860 476672
rect 319076 476620 319128 476672
rect 271788 476552 271840 476604
rect 330208 476552 330260 476604
rect 266268 476484 266320 476536
rect 326896 476484 326948 476536
rect 256608 476416 256660 476468
rect 318432 476416 318484 476468
rect 318708 476416 318760 476468
rect 336004 476416 336056 476468
rect 262128 476348 262180 476400
rect 323032 476348 323084 476400
rect 326988 476348 327040 476400
rect 338764 476348 338816 476400
rect 309048 476280 309100 476332
rect 329104 476280 329156 476332
rect 311808 476212 311860 476264
rect 331864 476212 331916 476264
rect 315948 476144 316000 476196
rect 334624 476144 334676 476196
rect 240048 476076 240100 476128
rect 313832 476076 313884 476128
rect 314568 476076 314620 476128
rect 333244 476076 333296 476128
rect 274548 475464 274600 475516
rect 331496 475464 331548 475516
rect 219072 475396 219124 475448
rect 321652 475396 321704 475448
rect 324228 475396 324280 475448
rect 352564 475396 352616 475448
rect 255596 475328 255648 475380
rect 371884 475328 371936 475380
rect 3424 474716 3476 474768
rect 287612 474716 287664 474768
rect 253756 474172 253808 474224
rect 329564 474172 329616 474224
rect 217508 474104 217560 474156
rect 323676 474104 323728 474156
rect 254860 474036 254912 474088
rect 369124 474036 369176 474088
rect 8944 473968 8996 474020
rect 284392 473968 284444 474020
rect 321468 473968 321520 474020
rect 356428 473968 356480 474020
rect 259276 472812 259328 472864
rect 294604 472812 294656 472864
rect 219164 472744 219216 472796
rect 319720 472744 319772 472796
rect 252928 472676 252980 472728
rect 367744 472676 367796 472728
rect 153200 472608 153252 472660
rect 275192 472608 275244 472660
rect 275928 472608 275980 472660
rect 354404 472608 354456 472660
rect 264796 471384 264848 471436
rect 295984 471384 296036 471436
rect 217600 471316 217652 471368
rect 327540 471316 327592 471368
rect 13084 471248 13136 471300
rect 286324 471248 286376 471300
rect 286508 471248 286560 471300
rect 338028 471248 338080 471300
rect 253204 470568 253256 470620
rect 580172 470568 580224 470620
rect 253848 470024 253900 470076
rect 315764 470024 315816 470076
rect 255228 469956 255280 470008
rect 330852 469956 330904 470008
rect 261484 469888 261536 469940
rect 378784 469888 378836 469940
rect 35164 469820 35216 469872
rect 285680 469820 285732 469872
rect 288348 469820 288400 469872
rect 339408 469820 339460 469872
rect 248236 468664 248288 468716
rect 320364 468664 320416 468716
rect 219256 468596 219308 468648
rect 317144 468596 317196 468648
rect 264704 468528 264756 468580
rect 462320 468528 462372 468580
rect 57244 468460 57296 468512
rect 283748 468460 283800 468512
rect 296628 468460 296680 468512
rect 343272 468460 343324 468512
rect 252376 467304 252428 467356
rect 326252 467304 326304 467356
rect 217692 467236 217744 467288
rect 325608 467236 325660 467288
rect 262772 467168 262824 467220
rect 527180 467168 527232 467220
rect 4804 467100 4856 467152
rect 281724 467100 281776 467152
rect 306288 467100 306340 467152
rect 348516 467100 348568 467152
rect 268936 465944 268988 465996
rect 291844 465944 291896 465996
rect 277216 465876 277268 465928
rect 355692 465876 355744 465928
rect 218888 465808 218940 465860
rect 307300 465808 307352 465860
rect 258816 465740 258868 465792
rect 373264 465740 373316 465792
rect 21364 465672 21416 465724
rect 279792 465672 279844 465724
rect 299388 465672 299440 465724
rect 344560 465672 344612 465724
rect 246948 464448 247000 464500
rect 317788 464448 317840 464500
rect 218060 464380 218112 464432
rect 273260 464380 273312 464432
rect 274456 464380 274508 464432
rect 351828 464380 351880 464432
rect 266728 464312 266780 464364
rect 396724 464312 396776 464364
rect 293868 463156 293920 463208
rect 341984 463156 342036 463208
rect 244188 463088 244240 463140
rect 309876 463088 309928 463140
rect 249708 463020 249760 463072
rect 322296 463020 322348 463072
rect 260840 462952 260892 463004
rect 391204 462952 391256 463004
rect 3240 462340 3292 462392
rect 288992 462340 289044 462392
rect 210424 461796 210476 461848
rect 285036 461796 285088 461848
rect 262036 461728 262088 461780
rect 338672 461728 338724 461780
rect 268016 461660 268068 461712
rect 364340 461660 364392 461712
rect 71780 461592 71832 461644
rect 276480 461592 276532 461644
rect 291108 461592 291160 461644
rect 340696 461592 340748 461644
rect 250996 460368 251048 460420
rect 313188 460368 313240 460420
rect 239404 460300 239456 460352
rect 309232 460300 309284 460352
rect 265992 460232 266044 460284
rect 359464 460232 359516 460284
rect 10324 460164 10376 460216
rect 278504 460164 278556 460216
rect 278596 460164 278648 460216
rect 357072 460164 357124 460216
rect 214564 459008 214616 459060
rect 281080 459008 281132 459060
rect 259368 458940 259420 458992
rect 334808 458940 334860 458992
rect 138664 458872 138716 458924
rect 274548 458872 274600 458924
rect 281448 458872 281500 458924
rect 335452 458872 335504 458924
rect 264060 458804 264112 458856
rect 494060 458804 494112 458856
rect 251088 457580 251140 457632
rect 324320 457580 324372 457632
rect 256516 457512 256568 457564
rect 332140 457512 332192 457564
rect 28264 457444 28316 457496
rect 280436 457444 280488 457496
rect 252284 456764 252336 456816
rect 580172 456764 580224 456816
rect 215944 456220 215996 456272
rect 279148 456220 279200 456272
rect 201500 456152 201552 456204
rect 272616 456152 272668 456204
rect 278688 456152 278740 456204
rect 334164 456152 334216 456204
rect 260656 456084 260708 456136
rect 336096 456084 336148 456136
rect 262128 456016 262180 456068
rect 442264 456016 442316 456068
rect 237196 454792 237248 454844
rect 311900 454792 311952 454844
rect 260104 454724 260156 454776
rect 377404 454724 377456 454776
rect 40040 454656 40092 454708
rect 277860 454656 277912 454708
rect 280068 454656 280120 454708
rect 358360 454656 358412 454708
rect 248328 453568 248380 453620
rect 310520 453568 310572 453620
rect 211804 453500 211856 453552
rect 283012 453500 283064 453552
rect 271696 453432 271748 453484
rect 349160 453432 349212 453484
rect 169760 453364 169812 453416
rect 273904 453364 273956 453416
rect 302148 453364 302200 453416
rect 345940 453364 345992 453416
rect 258172 453296 258224 453348
rect 363604 453296 363656 453348
rect 273168 452072 273220 452124
rect 350540 452072 350592 452124
rect 207664 452004 207716 452056
rect 286968 452004 287020 452056
rect 256240 451936 256292 451988
rect 360844 451936 360896 451988
rect 108304 451868 108356 451920
rect 275836 451868 275888 451920
rect 284208 451868 284260 451920
rect 336740 451868 336792 451920
rect 260748 450644 260800 450696
rect 337384 450644 337436 450696
rect 254216 450576 254268 450628
rect 358084 450576 358136 450628
rect 88340 450508 88392 450560
rect 277124 450508 277176 450560
rect 277308 450508 277360 450560
rect 332784 450508 332836 450560
rect 245568 449692 245620 449744
rect 312544 449692 312596 449744
rect 245476 449624 245528 449676
rect 315120 449624 315172 449676
rect 266176 449556 266228 449608
rect 342628 449556 342680 449608
rect 264888 449488 264940 449540
rect 341340 449488 341392 449540
rect 267648 449420 267700 449472
rect 343916 449420 343968 449472
rect 263508 449352 263560 449404
rect 340052 449352 340104 449404
rect 269028 449284 269080 449336
rect 346584 449284 346636 449336
rect 270408 449216 270460 449268
rect 347872 449216 347924 449268
rect 267556 449148 267608 449200
rect 345296 449148 345348 449200
rect 257988 447992 258040 448044
rect 333428 447992 333480 448044
rect 252468 447924 252520 447976
rect 328276 447924 328328 447976
rect 274364 447856 274416 447908
rect 353116 447856 353168 447908
rect 217324 447788 217376 447840
rect 307944 447788 307996 447840
rect 267372 446700 267424 446752
rect 412640 446700 412692 446752
rect 265348 446632 265400 446684
rect 477500 446632 477552 446684
rect 263416 446564 263468 446616
rect 542360 446564 542412 446616
rect 4160 446496 4212 446548
rect 288256 446496 288308 446548
rect 259460 446428 259512 446480
rect 580264 446428 580316 446480
rect 257528 446360 257580 446412
rect 580356 446360 580408 446412
rect 206284 446020 206336 446072
rect 300124 446020 300176 446072
rect 203616 445952 203668 446004
rect 298100 445952 298152 446004
rect 192484 445884 192536 445936
rect 302700 445884 302752 445936
rect 235908 445816 235960 445868
rect 373264 445816 373316 445868
rect 8944 445748 8996 445800
rect 296812 445748 296864 445800
rect 231124 444864 231176 444916
rect 290280 444864 290332 444916
rect 225604 444796 225656 444848
rect 295524 444796 295576 444848
rect 199384 444728 199436 444780
rect 303988 444728 304040 444780
rect 249708 444660 249760 444712
rect 378784 444660 378836 444712
rect 100024 444592 100076 444644
rect 291568 444592 291620 444644
rect 98644 444524 98696 444576
rect 293500 444524 293552 444576
rect 7564 444456 7616 444508
rect 289636 444456 289688 444508
rect 244464 444388 244516 444440
rect 578884 444388 578936 444440
rect 245752 444116 245804 444168
rect 362224 444116 362276 444168
rect 336004 444048 336056 444100
rect 355048 444048 355100 444100
rect 334624 443980 334676 444032
rect 353760 443980 353812 444032
rect 252560 443912 252612 443964
rect 301412 443912 301464 443964
rect 331864 443912 331916 443964
rect 351184 443912 351236 443964
rect 239220 443844 239272 443896
rect 282920 443844 282972 443896
rect 294604 443844 294656 443896
rect 321008 443844 321060 443896
rect 333244 443844 333296 443896
rect 352472 443844 352524 443896
rect 94504 443776 94556 443828
rect 294880 443776 294932 443828
rect 295984 443776 296036 443828
rect 324964 443776 325016 443828
rect 338764 443776 338816 443828
rect 359004 443776 359056 443828
rect 219348 443708 219400 443760
rect 270592 443708 270644 443760
rect 291844 443708 291896 443760
rect 328920 443708 328972 443760
rect 329104 443708 329156 443760
rect 349804 443708 349856 443760
rect 217784 443640 217836 443692
rect 271972 443640 272024 443692
rect 303528 443640 303580 443692
rect 347228 443640 347280 443692
rect 352564 443640 352616 443692
rect 357716 443640 357768 443692
rect 246396 443572 246448 443624
rect 277400 443572 277452 443624
rect 241152 443504 241204 443556
rect 274732 443504 274784 443556
rect 245108 443436 245160 443488
rect 288348 443436 288400 443488
rect 248328 443368 248380 443420
rect 276112 443368 276164 443420
rect 279516 443368 279568 443420
rect 296168 443368 296220 443420
rect 229744 443300 229796 443352
rect 253204 443300 253256 443352
rect 253572 443300 253624 443352
rect 224224 443232 224276 443284
rect 292856 443232 292908 443284
rect 196716 443164 196768 443216
rect 298744 443164 298796 443216
rect 359648 443164 359700 443216
rect 388444 443164 388496 443216
rect 140780 443096 140832 443148
rect 250352 443096 250404 443148
rect 362500 443096 362552 443148
rect 233976 443028 234028 443080
rect 246948 443028 247000 443080
rect 269028 443028 269080 443080
rect 292212 443028 292264 443080
rect 360292 443028 360344 443080
rect 581092 443028 581144 443080
rect 250996 442960 251048 443012
rect 268568 442960 268620 443012
rect 274640 442960 274692 443012
rect 294144 442960 294196 443012
rect 360936 442960 360988 443012
rect 582380 442960 582432 443012
rect 231216 442484 231268 442536
rect 290924 442484 290976 442536
rect 3608 442416 3660 442468
rect 274640 442416 274692 442468
rect 288348 442416 288400 442468
rect 580816 442416 580868 442468
rect 3516 442348 3568 442400
rect 279516 442348 279568 442400
rect 282920 442348 282972 442400
rect 580632 442348 580684 442400
rect 3700 442212 3752 442264
rect 269028 442280 269080 442332
rect 274732 442280 274784 442332
rect 580724 442280 580776 442332
rect 268568 442212 268620 442264
rect 580080 442212 580132 442264
rect 200764 442144 200816 442196
rect 302056 442144 302108 442196
rect 198004 442076 198056 442128
rect 300768 442076 300820 442128
rect 248972 442008 249024 442060
rect 362408 442008 362460 442060
rect 247040 441940 247092 441992
rect 362316 441940 362368 441992
rect 241796 441872 241848 441924
rect 374736 441872 374788 441924
rect 64144 441804 64196 441856
rect 306656 441804 306708 441856
rect 242440 441736 242492 441788
rect 577596 441736 577648 441788
rect 237196 441668 237248 441720
rect 580448 441668 580500 441720
rect 233332 441600 233384 441652
rect 577504 441600 577556 441652
rect 290004 441396 290056 441448
rect 294604 441396 294656 441448
rect 3424 440852 3476 440904
rect 252560 441124 252612 441176
rect 290740 441124 290792 441176
rect 207664 440580 207716 440632
rect 240784 440988 240836 441040
rect 247960 440988 248012 441040
rect 252008 440988 252060 441040
rect 276112 440988 276164 441040
rect 277400 440988 277452 441040
rect 289820 440988 289872 441040
rect 290004 440988 290056 441040
rect 293592 441260 293644 441312
rect 293408 441192 293460 441244
rect 294604 441192 294656 441244
rect 293408 440988 293460 441040
rect 25504 440308 25556 440360
rect 293592 440988 293644 441040
rect 293684 440988 293736 441040
rect 293776 440988 293828 441040
rect 303068 440988 303120 441040
rect 304356 440988 304408 441040
rect 580908 440920 580960 440972
rect 580172 440852 580224 440904
rect 363604 440512 363656 440564
rect 377404 440444 377456 440496
rect 371976 440376 372028 440428
rect 3332 423580 3384 423632
rect 7564 423580 7616 423632
rect 363604 419432 363656 419484
rect 579988 419432 580040 419484
rect 2964 411204 3016 411256
rect 231216 411204 231268 411256
rect 362500 405628 362552 405680
rect 579804 405628 579856 405680
rect 3056 398760 3108 398812
rect 231124 398760 231176 398812
rect 362408 379448 362460 379500
rect 580080 379448 580132 379500
rect 3792 378768 3844 378820
rect 224224 378768 224276 378820
rect 97816 377408 97868 377460
rect 229744 377408 229796 377460
rect 154764 374824 154816 374876
rect 173164 374824 173216 374876
rect 110972 374756 111024 374808
rect 228364 374756 228416 374808
rect 100668 374688 100720 374740
rect 229836 374688 229888 374740
rect 126428 374620 126480 374672
rect 170588 374620 170640 374672
rect 121276 374552 121328 374604
rect 170956 374552 171008 374604
rect 165528 374484 165580 374536
rect 227076 374484 227128 374536
rect 105820 374416 105872 374468
rect 171784 374416 171836 374468
rect 157340 374348 157392 374400
rect 228548 374348 228600 374400
rect 108396 374280 108448 374332
rect 180064 374280 180116 374332
rect 152188 374212 152240 374264
rect 231216 374212 231268 374264
rect 147036 374144 147088 374196
rect 229744 374144 229796 374196
rect 139308 374008 139360 374060
rect 155868 374008 155920 374060
rect 162492 374008 162544 374060
rect 170404 374008 170456 374060
rect 32404 373124 32456 373176
rect 165068 373124 165120 373176
rect 165528 373124 165580 373176
rect 123852 373056 123904 373108
rect 174544 373056 174596 373108
rect 118700 372988 118752 373040
rect 173256 372988 173308 373040
rect 103244 372920 103296 372972
rect 173440 372920 173492 372972
rect 134156 372852 134208 372904
rect 226984 372852 227036 372904
rect 131580 372784 131632 372836
rect 231124 372784 231176 372836
rect 129004 372716 129056 372768
rect 228456 372716 228508 372768
rect 113548 372648 113600 372700
rect 229928 372648 229980 372700
rect 149612 372580 149664 372632
rect 170496 372580 170548 372632
rect 3148 372512 3200 372564
rect 100024 372512 100076 372564
rect 124772 371832 124824 371884
rect 116400 371628 116452 371680
rect 125692 371764 125744 371816
rect 128268 371832 128320 371884
rect 97724 371560 97776 371612
rect 128268 371696 128320 371748
rect 124680 371560 124732 371612
rect 124772 371560 124824 371612
rect 97632 371492 97684 371544
rect 99840 371424 99892 371476
rect 97908 371356 97960 371408
rect 125692 371560 125744 371612
rect 137008 371832 137060 371884
rect 138480 371832 138532 371884
rect 138020 371764 138072 371816
rect 144000 371764 144052 371816
rect 167920 371696 167972 371748
rect 170772 371696 170824 371748
rect 135214 371560 135266 371612
rect 137928 371560 137980 371612
rect 138020 371560 138072 371612
rect 138480 371560 138532 371612
rect 144000 371560 144052 371612
rect 144184 371560 144236 371612
rect 144736 371628 144788 371680
rect 174636 371628 174688 371680
rect 228640 371560 228692 371612
rect 230020 371492 230072 371544
rect 231308 371424 231360 371476
rect 231492 371356 231544 371408
rect 231400 371288 231452 371340
rect 231584 371220 231636 371272
rect 172336 368500 172388 368552
rect 232228 368500 232280 368552
rect 169944 367888 169996 367940
rect 170680 367888 170732 367940
rect 172428 365712 172480 365764
rect 231676 365712 231728 365764
rect 378784 365644 378836 365696
rect 580080 365644 580132 365696
rect 172336 362924 172388 362976
rect 230112 362924 230164 362976
rect 171692 357416 171744 357468
rect 228732 357416 228784 357468
rect 172428 351908 172480 351960
rect 224224 351908 224276 351960
rect 172428 346400 172480 346452
rect 220084 346400 220136 346452
rect 171140 345040 171192 345092
rect 178684 345040 178736 345092
rect 172428 336744 172480 336796
rect 225696 336744 225748 336796
rect 172428 333956 172480 334008
rect 225788 333956 225840 334008
rect 172428 331236 172480 331288
rect 230204 331236 230256 331288
rect 172428 325660 172480 325712
rect 232228 325660 232280 325712
rect 362316 325592 362368 325644
rect 580172 325592 580224 325644
rect 171324 322940 171376 322992
rect 231768 322940 231820 322992
rect 171508 320152 171560 320204
rect 231032 320152 231084 320204
rect 2964 320084 3016 320136
rect 98644 320084 98696 320136
rect 171508 317432 171560 317484
rect 231860 317432 231912 317484
rect 172428 314644 172480 314696
rect 230388 314644 230440 314696
rect 377404 313216 377456 313268
rect 580172 313216 580224 313268
rect 172428 311856 172480 311908
rect 232044 311856 232096 311908
rect 172336 311380 172388 311432
rect 230848 311380 230900 311432
rect 171876 311244 171928 311296
rect 232228 311244 232280 311296
rect 172244 311176 172296 311228
rect 230940 311176 230992 311228
rect 178684 311108 178736 311160
rect 232228 311108 232280 311160
rect 230388 310700 230440 310752
rect 172152 310564 172204 310616
rect 230756 310564 230808 310616
rect 227076 310496 227128 310548
rect 235448 310496 235500 310548
rect 255412 310496 255464 310548
rect 255596 310496 255648 310548
rect 273536 310496 273588 310548
rect 273720 310496 273772 310548
rect 315028 310496 315080 310548
rect 315396 310496 315448 310548
rect 232596 310428 232648 310480
rect 231952 310360 232004 310412
rect 230112 310292 230164 310344
rect 233240 310292 233292 310344
rect 244464 310292 244516 310344
rect 230940 310224 230992 310276
rect 231952 310224 232004 310276
rect 232044 310224 232096 310276
rect 236276 310224 236328 310276
rect 231860 310156 231912 310208
rect 241796 310156 241848 310208
rect 230848 310088 230900 310140
rect 232044 310088 232096 310140
rect 171968 310020 172020 310072
rect 237472 310020 237524 310072
rect 225696 309952 225748 310004
rect 238944 309952 238996 310004
rect 286968 309952 287020 310004
rect 287612 309952 287664 310004
rect 231768 309884 231820 309936
rect 239496 309884 239548 309936
rect 230204 309748 230256 309800
rect 241704 309748 241756 309800
rect 228732 309544 228784 309596
rect 242992 309544 243044 309596
rect 232136 309476 232188 309528
rect 249064 309476 249116 309528
rect 231676 309408 231728 309460
rect 247500 309408 247552 309460
rect 241796 309340 241848 309392
rect 249616 309340 249668 309392
rect 231032 309272 231084 309324
rect 249800 309272 249852 309324
rect 170680 309204 170732 309256
rect 234160 309204 234212 309256
rect 172244 309136 172296 309188
rect 235908 309136 235960 309188
rect 237472 309136 237524 309188
rect 230020 309068 230072 309120
rect 233608 309068 233660 309120
rect 234068 309068 234120 309120
rect 238576 309068 238628 309120
rect 238760 309068 238812 309120
rect 347688 309068 347740 309120
rect 229928 309000 229980 309052
rect 235356 309000 235408 309052
rect 239772 309000 239824 309052
rect 246764 309000 246816 309052
rect 326160 309000 326212 309052
rect 340144 309000 340196 309052
rect 348976 309000 349028 309052
rect 350908 309000 350960 309052
rect 231400 308932 231452 308984
rect 237012 308932 237064 308984
rect 237104 308932 237156 308984
rect 247132 308932 247184 308984
rect 310336 308932 310388 308984
rect 230756 308864 230808 308916
rect 252836 308864 252888 308916
rect 226984 308796 227036 308848
rect 243360 308796 243412 308848
rect 251088 308796 251140 308848
rect 257804 308796 257856 308848
rect 228456 308728 228508 308780
rect 242164 308728 242216 308780
rect 247960 308728 248012 308780
rect 254400 308728 254452 308780
rect 231124 308660 231176 308712
rect 237104 308660 237156 308712
rect 237288 308660 237340 308712
rect 241612 308660 241664 308712
rect 246304 308660 246356 308712
rect 255964 308660 256016 308712
rect 170496 308592 170548 308644
rect 239772 308592 239824 308644
rect 174544 308524 174596 308576
rect 242348 308592 242400 308644
rect 250904 308592 250956 308644
rect 259552 308796 259604 308848
rect 333980 308932 334032 308984
rect 334256 308932 334308 308984
rect 336740 308932 336792 308984
rect 337384 308932 337436 308984
rect 350632 308932 350684 308984
rect 351368 308932 351420 308984
rect 354220 309068 354272 309120
rect 367560 309068 367612 309120
rect 354588 309000 354640 309052
rect 367836 309000 367888 309052
rect 366180 308932 366232 308984
rect 312176 308864 312228 308916
rect 355232 308864 355284 308916
rect 355324 308864 355376 308916
rect 367376 308864 367428 308916
rect 356888 308796 356940 308848
rect 358820 308796 358872 308848
rect 359188 308796 359240 308848
rect 258172 308728 258224 308780
rect 258816 308728 258868 308780
rect 267096 308728 267148 308780
rect 281264 308728 281316 308780
rect 303804 308728 303856 308780
rect 355600 308728 355652 308780
rect 356060 308728 356112 308780
rect 363512 308728 363564 308780
rect 232412 308456 232464 308508
rect 237288 308456 237340 308508
rect 237932 308456 237984 308508
rect 241980 308524 242032 308576
rect 242808 308524 242860 308576
rect 252468 308524 252520 308576
rect 253204 308524 253256 308576
rect 267188 308660 267240 308712
rect 287244 308660 287296 308712
rect 287520 308660 287572 308712
rect 302700 308660 302752 308712
rect 355416 308660 355468 308712
rect 356520 308660 356572 308712
rect 367284 308660 367336 308712
rect 260564 308592 260616 308644
rect 268752 308592 268804 308644
rect 287152 308592 287204 308644
rect 258816 308524 258868 308576
rect 271604 308524 271656 308576
rect 240140 308456 240192 308508
rect 241060 308456 241112 308508
rect 271144 308456 271196 308508
rect 273444 308456 273496 308508
rect 236184 308388 236236 308440
rect 236828 308388 236880 308440
rect 238852 308388 238904 308440
rect 239312 308388 239364 308440
rect 240232 308388 240284 308440
rect 240692 308388 240744 308440
rect 242992 308388 243044 308440
rect 243544 308388 243596 308440
rect 174636 308320 174688 308372
rect 238208 308320 238260 308372
rect 238944 308320 238996 308372
rect 239864 308320 239916 308372
rect 240324 308320 240376 308372
rect 240876 308320 240928 308372
rect 236092 308252 236144 308304
rect 236368 308252 236420 308304
rect 237564 308252 237616 308304
rect 237840 308252 237892 308304
rect 246396 308320 246448 308372
rect 231584 308184 231636 308236
rect 243176 308252 243228 308304
rect 244096 308252 244148 308304
rect 236092 308116 236144 308168
rect 236644 308116 236696 308168
rect 232044 308048 232096 308100
rect 237932 308048 237984 308100
rect 231952 307980 232004 308032
rect 245844 307980 245896 308032
rect 251088 307912 251140 307964
rect 252192 307912 252244 307964
rect 272708 308388 272760 308440
rect 284300 308388 284352 308440
rect 285128 308388 285180 308440
rect 286140 308388 286192 308440
rect 286416 308388 286468 308440
rect 288532 308592 288584 308644
rect 302332 308592 302384 308644
rect 355692 308592 355744 308644
rect 356980 308592 357032 308644
rect 369952 308592 370004 308644
rect 287796 308456 287848 308508
rect 287980 308456 288032 308508
rect 287336 308252 287388 308304
rect 287428 308252 287480 308304
rect 287244 308184 287296 308236
rect 301688 308524 301740 308576
rect 355048 308524 355100 308576
rect 357256 308524 357308 308576
rect 370504 308524 370556 308576
rect 289820 308456 289872 308508
rect 290280 308456 290332 308508
rect 291292 308456 291344 308508
rect 291660 308456 291712 308508
rect 300768 308456 300820 308508
rect 356796 308456 356848 308508
rect 288808 308388 288860 308440
rect 289728 308388 289780 308440
rect 291476 308388 291528 308440
rect 292396 308388 292448 308440
rect 299664 308388 299716 308440
rect 354680 308388 354732 308440
rect 354864 308388 354916 308440
rect 355876 308388 355928 308440
rect 359280 308388 359332 308440
rect 359924 308388 359976 308440
rect 288532 308320 288584 308372
rect 291660 308320 291712 308372
rect 292212 308320 292264 308372
rect 331220 308320 331272 308372
rect 332232 308320 332284 308372
rect 333060 308320 333112 308372
rect 333612 308320 333664 308372
rect 334440 308320 334492 308372
rect 334900 308320 334952 308372
rect 335820 308320 335872 308372
rect 336464 308320 336516 308372
rect 338488 308320 338540 308372
rect 339316 308320 339368 308372
rect 352104 308320 352156 308372
rect 352472 308320 352524 308372
rect 353392 308320 353444 308372
rect 354036 308320 354088 308372
rect 288624 308252 288676 308304
rect 289084 308252 289136 308304
rect 290280 308252 290332 308304
rect 291016 308252 291068 308304
rect 291200 308252 291252 308304
rect 291752 308252 291804 308304
rect 331312 308252 331364 308304
rect 331772 308252 331824 308304
rect 332692 308252 332744 308304
rect 333428 308252 333480 308304
rect 334532 308252 334584 308304
rect 335084 308252 335136 308304
rect 335544 308252 335596 308304
rect 336280 308252 336332 308304
rect 336832 308252 336884 308304
rect 337108 308252 337160 308304
rect 338212 308252 338264 308304
rect 338672 308252 338724 308304
rect 339868 308252 339920 308304
rect 340236 308252 340288 308304
rect 350540 308252 350592 308304
rect 351000 308252 351052 308304
rect 351184 308252 351236 308304
rect 352012 308252 352064 308304
rect 352196 308252 352248 308304
rect 352656 308252 352708 308304
rect 353300 308252 353352 308304
rect 354404 308252 354456 308304
rect 288716 308184 288768 308236
rect 289544 308184 289596 308236
rect 332600 308184 332652 308236
rect 333796 308184 333848 308236
rect 334072 308184 334124 308236
rect 334716 308184 334768 308236
rect 335360 308184 335412 308236
rect 336096 308184 336148 308236
rect 338120 308184 338172 308236
rect 338948 308184 339000 308236
rect 339684 308184 339736 308236
rect 340052 308184 340104 308236
rect 350908 308184 350960 308236
rect 351736 308184 351788 308236
rect 352840 308184 352892 308236
rect 353024 308184 353076 308236
rect 353852 308184 353904 308236
rect 367652 308320 367704 308372
rect 284668 308116 284720 308168
rect 285496 308116 285548 308168
rect 285864 308116 285916 308168
rect 286048 308116 286100 308168
rect 291200 308116 291252 308168
rect 292028 308116 292080 308168
rect 331312 308116 331364 308168
rect 332048 308116 332100 308168
rect 332508 308116 332560 308168
rect 332876 308116 332928 308168
rect 334164 308116 334216 308168
rect 335268 308116 335320 308168
rect 335452 308116 335504 308168
rect 336648 308116 336700 308168
rect 336924 308116 336976 308168
rect 337292 308116 337344 308168
rect 338212 308116 338264 308168
rect 339132 308116 339184 308168
rect 352012 308116 352064 308168
rect 365076 308252 365128 308304
rect 357348 308184 357400 308236
rect 357808 308184 357860 308236
rect 359096 308184 359148 308236
rect 359740 308184 359792 308236
rect 355784 308116 355836 308168
rect 284760 308048 284812 308100
rect 285312 308048 285364 308100
rect 354680 308048 354732 308100
rect 356980 308048 357032 308100
rect 357624 308048 357676 308100
rect 357992 308048 358044 308100
rect 359188 308116 359240 308168
rect 360108 308116 360160 308168
rect 366364 308048 366416 308100
rect 351920 307980 351972 308032
rect 352564 307980 352616 308032
rect 353484 307980 353536 308032
rect 364892 307980 364944 308032
rect 256240 307912 256292 307964
rect 262404 307912 262456 307964
rect 356704 307912 356756 307964
rect 359556 307912 359608 307964
rect 250444 307844 250496 307896
rect 250536 307844 250588 307896
rect 250904 307844 250956 307896
rect 252008 307844 252060 307896
rect 258816 307844 258868 307896
rect 261760 307844 261812 307896
rect 269856 307844 269908 307896
rect 282920 307844 282972 307896
rect 283288 307844 283340 307896
rect 283380 307844 283432 307896
rect 284024 307844 284076 307896
rect 285680 307844 285732 307896
rect 285956 307844 286008 307896
rect 289820 307844 289872 307896
rect 290648 307844 290700 307896
rect 336924 307844 336976 307896
rect 337752 307844 337804 307896
rect 354956 307844 355008 307896
rect 367468 307844 367520 307896
rect 247776 307776 247828 307828
rect 248512 307776 248564 307828
rect 250628 307776 250680 307828
rect 251364 307776 251416 307828
rect 257712 307776 257764 307828
rect 259000 307776 259052 307828
rect 264428 307776 264480 307828
rect 267004 307776 267056 307828
rect 284392 307776 284444 307828
rect 284852 307776 284904 307828
rect 285864 307776 285916 307828
rect 286876 307776 286928 307828
rect 317328 307776 317380 307828
rect 318064 307776 318116 307828
rect 336832 307776 336884 307828
rect 337936 307776 337988 307828
rect 348424 307776 348476 307828
rect 350356 307776 350408 307828
rect 228364 307708 228416 307760
rect 246580 307708 246632 307760
rect 282920 307708 282972 307760
rect 283748 307708 283800 307760
rect 285680 307708 285732 307760
rect 286508 307708 286560 307760
rect 354956 307708 355008 307760
rect 355140 307708 355192 307760
rect 171416 307640 171468 307692
rect 246948 307640 247000 307692
rect 331588 307640 331640 307692
rect 332416 307640 332468 307692
rect 171784 307572 171836 307624
rect 244280 307572 244332 307624
rect 354772 307572 354824 307624
rect 355508 307572 355560 307624
rect 229744 307504 229796 307556
rect 250260 307504 250312 307556
rect 180064 307436 180116 307488
rect 244832 307436 244884 307488
rect 220084 307368 220136 307420
rect 242532 307368 242584 307420
rect 229836 307300 229888 307352
rect 252284 307300 252336 307352
rect 332968 307300 333020 307352
rect 333244 307300 333296 307352
rect 224224 307232 224276 307284
rect 243728 307232 243780 307284
rect 339592 307232 339644 307284
rect 340604 307232 340656 307284
rect 170404 307164 170456 307216
rect 249984 307164 250036 307216
rect 314108 307164 314160 307216
rect 378784 307164 378836 307216
rect 170588 307096 170640 307148
rect 238392 307096 238444 307148
rect 243084 307096 243136 307148
rect 243912 307096 243964 307148
rect 200120 307028 200172 307080
rect 284944 307096 284996 307148
rect 317788 307096 317840 307148
rect 402980 307096 403032 307148
rect 283104 307028 283156 307080
rect 283932 307028 283984 307080
rect 340420 307028 340472 307080
rect 543740 307028 543792 307080
rect 173164 306960 173216 307012
rect 239680 306960 239732 307012
rect 253020 306960 253072 307012
rect 281724 306960 281776 307012
rect 282000 306960 282052 307012
rect 297180 306960 297232 307012
rect 321836 306960 321888 307012
rect 322112 306960 322164 307012
rect 252836 306756 252888 306808
rect 297088 306756 297140 306808
rect 330116 306824 330168 306876
rect 356060 306824 356112 306876
rect 357072 306824 357124 306876
rect 357532 306824 357584 306876
rect 358360 306824 358412 306876
rect 267924 306688 267976 306740
rect 295616 306688 295668 306740
rect 300860 306688 300912 306740
rect 301136 306688 301188 306740
rect 252744 306484 252796 306536
rect 253112 306484 253164 306536
rect 256608 306484 256660 306536
rect 257252 306484 257304 306536
rect 342720 306688 342772 306740
rect 360660 306688 360712 306740
rect 328644 306620 328696 306672
rect 328920 306620 328972 306672
rect 330116 306620 330168 306672
rect 309324 306552 309376 306604
rect 316224 306552 316276 306604
rect 316868 306552 316920 306604
rect 317696 306552 317748 306604
rect 318248 306552 318300 306604
rect 252652 306416 252704 306468
rect 253480 306416 253532 306468
rect 256792 306416 256844 306468
rect 257436 306416 257488 306468
rect 267924 306416 267976 306468
rect 269212 306416 269264 306468
rect 269672 306416 269724 306468
rect 270684 306416 270736 306468
rect 270960 306416 271012 306468
rect 277400 306416 277452 306468
rect 277860 306416 277912 306468
rect 278780 306416 278832 306468
rect 279792 306416 279844 306468
rect 280344 306416 280396 306468
rect 280804 306416 280856 306468
rect 295616 306416 295668 306468
rect 305092 306416 305144 306468
rect 305736 306416 305788 306468
rect 248512 306348 248564 306400
rect 249248 306348 249300 306400
rect 264980 306348 265032 306400
rect 265900 306348 265952 306400
rect 266636 306348 266688 306400
rect 267004 306348 267056 306400
rect 272156 306348 272208 306400
rect 272340 306348 272392 306400
rect 273720 306348 273772 306400
rect 274456 306348 274508 306400
rect 279056 306348 279108 306400
rect 279424 306348 279476 306400
rect 294144 306348 294196 306400
rect 294880 306348 294932 306400
rect 295432 306348 295484 306400
rect 296168 306348 296220 306400
rect 299572 306348 299624 306400
rect 300584 306348 300636 306400
rect 301044 306348 301096 306400
rect 302056 306348 302108 306400
rect 3332 306280 3384 306332
rect 94504 306280 94556 306332
rect 169852 306280 169904 306332
rect 243268 306280 243320 306332
rect 247132 306280 247184 306332
rect 247868 306280 247920 306332
rect 248604 306280 248656 306332
rect 249432 306280 249484 306332
rect 251732 306280 251784 306332
rect 252100 306280 252152 306332
rect 253112 306280 253164 306332
rect 253664 306280 253716 306332
rect 253940 306280 253992 306332
rect 255136 306280 255188 306332
rect 255320 306280 255372 306332
rect 255596 306280 255648 306332
rect 258540 306280 258592 306332
rect 259368 306280 259420 306332
rect 259644 306280 259696 306332
rect 260656 306280 260708 306332
rect 262404 306280 262456 306332
rect 263140 306280 263192 306332
rect 265348 306280 265400 306332
rect 266268 306280 266320 306332
rect 266544 306280 266596 306332
rect 267372 306280 267424 306332
rect 267740 306280 267792 306332
rect 268016 306280 268068 306332
rect 272064 306280 272116 306332
rect 272524 306280 272576 306332
rect 273628 306280 273680 306332
rect 274088 306280 274140 306332
rect 276204 306280 276256 306332
rect 276756 306280 276808 306332
rect 277584 306280 277636 306332
rect 278228 306280 278280 306332
rect 278872 306280 278924 306332
rect 279148 306280 279200 306332
rect 294328 306280 294380 306332
rect 295064 306280 295116 306332
rect 295524 306280 295576 306332
rect 295984 306280 296036 306332
rect 296812 306280 296864 306332
rect 297548 306280 297600 306332
rect 298560 306280 298612 306332
rect 299204 306280 299256 306332
rect 299480 306280 299532 306332
rect 300400 306280 300452 306332
rect 301136 306280 301188 306332
rect 301504 306280 301556 306332
rect 302240 306280 302292 306332
rect 303252 306280 303304 306332
rect 303804 306280 303856 306332
rect 304356 306280 304408 306332
rect 305460 306280 305512 306332
rect 307300 306416 307352 306468
rect 307944 306416 307996 306468
rect 308404 306416 308456 306468
rect 308128 306280 308180 306332
rect 308588 306280 308640 306332
rect 215208 306212 215260 306264
rect 288532 306212 288584 306264
rect 294236 306212 294288 306264
rect 295248 306212 295300 306264
rect 303988 306212 304040 306264
rect 304632 306212 304684 306264
rect 305184 306212 305236 306264
rect 306564 306212 306616 306264
rect 308220 306212 308272 306264
rect 308772 306212 308824 306264
rect 310612 306416 310664 306468
rect 310888 306416 310940 306468
rect 311900 306416 311952 306468
rect 312452 306416 312504 306468
rect 319076 306416 319128 306468
rect 319352 306416 319404 306468
rect 313280 306348 313332 306400
rect 313924 306348 313976 306400
rect 316040 306348 316092 306400
rect 316224 306348 316276 306400
rect 317696 306348 317748 306400
rect 318708 306348 318760 306400
rect 318800 306348 318852 306400
rect 319444 306348 319496 306400
rect 320364 306348 320416 306400
rect 320640 306348 320692 306400
rect 310980 306280 311032 306332
rect 311624 306280 311676 306332
rect 313556 306280 313608 306332
rect 313832 306280 313884 306332
rect 314752 306280 314804 306332
rect 315488 306280 315540 306332
rect 317604 306280 317656 306332
rect 318340 306280 318392 306332
rect 319168 306280 319220 306332
rect 319812 306280 319864 306332
rect 320180 306280 320232 306332
rect 321192 306280 321244 306332
rect 321836 306280 321888 306332
rect 322664 306280 322716 306332
rect 323308 306552 323360 306604
rect 325792 306552 325844 306604
rect 326436 306552 326488 306604
rect 328460 306552 328512 306604
rect 329104 306552 329156 306604
rect 324412 306484 324464 306536
rect 325240 306484 325292 306536
rect 340880 306484 340932 306536
rect 341708 306484 341760 306536
rect 323216 306280 323268 306332
rect 323492 306280 323544 306332
rect 324780 306416 324832 306468
rect 342720 306416 342772 306468
rect 360660 306416 360712 306468
rect 325792 306348 325844 306400
rect 326896 306348 326948 306400
rect 340880 306348 340932 306400
rect 341432 306348 341484 306400
rect 347780 306348 347832 306400
rect 349068 306348 349120 306400
rect 325884 306280 325936 306332
rect 326528 306280 326580 306332
rect 327448 306280 327500 306332
rect 327632 306280 327684 306332
rect 328552 306280 328604 306332
rect 329748 306280 329800 306332
rect 329840 306280 329892 306332
rect 330392 306280 330444 306332
rect 341156 306280 341208 306332
rect 342168 306280 342220 306332
rect 342628 306280 342680 306332
rect 343272 306280 343324 306332
rect 343824 306280 343876 306332
rect 344652 306280 344704 306332
rect 345020 306280 345072 306332
rect 345756 306280 345808 306332
rect 347872 306280 347924 306332
rect 348240 306280 348292 306332
rect 354864 306280 354916 306332
rect 370412 306280 370464 306332
rect 309508 306212 309560 306264
rect 310704 306212 310756 306264
rect 311256 306212 311308 306264
rect 317420 306212 317472 306264
rect 318524 306212 318576 306264
rect 321560 306212 321612 306264
rect 322020 306212 322072 306264
rect 322940 306212 322992 306264
rect 323400 306212 323452 306264
rect 324044 306212 324096 306264
rect 324412 306212 324464 306264
rect 324504 306212 324556 306264
rect 325332 306212 325384 306264
rect 327080 306212 327132 306264
rect 328276 306212 328328 306264
rect 328736 306212 328788 306264
rect 329380 306212 329432 306264
rect 330024 306212 330076 306264
rect 331128 306212 331180 306264
rect 340972 306212 341024 306264
rect 341800 306212 341852 306264
rect 342352 306212 342404 306264
rect 342904 306212 342956 306264
rect 343732 306212 343784 306264
rect 344284 306212 344336 306264
rect 345204 306212 345256 306264
rect 345388 306212 345440 306264
rect 352380 306212 352432 306264
rect 360200 306212 360252 306264
rect 360292 306212 360344 306264
rect 360844 306212 360896 306264
rect 218980 306144 219032 306196
rect 293500 306144 293552 306196
rect 295616 306144 295668 306196
rect 296352 306144 296404 306196
rect 309140 306144 309192 306196
rect 310152 306144 310204 306196
rect 310796 306144 310848 306196
rect 311808 306144 311860 306196
rect 311992 306144 312044 306196
rect 313188 306144 313240 306196
rect 313556 306144 313608 306196
rect 314292 306144 314344 306196
rect 314936 306144 314988 306196
rect 315856 306144 315908 306196
rect 316408 306144 316460 306196
rect 317144 306144 317196 306196
rect 317788 306144 317840 306196
rect 318156 306144 318208 306196
rect 318984 306144 319036 306196
rect 319628 306144 319680 306196
rect 321744 306144 321796 306196
rect 322480 306144 322532 306196
rect 323032 306144 323084 306196
rect 323860 306144 323912 306196
rect 324596 306144 324648 306196
rect 325608 306144 325660 306196
rect 328828 306144 328880 306196
rect 329564 306144 329616 306196
rect 341248 306144 341300 306196
rect 341616 306144 341668 306196
rect 352196 306144 352248 306196
rect 368664 306144 368716 306196
rect 216404 306076 216456 306128
rect 291476 306076 291528 306128
rect 305000 306076 305052 306128
rect 305368 306076 305420 306128
rect 305460 306076 305512 306128
rect 306288 306076 306340 306128
rect 307944 306076 307996 306128
rect 308956 306076 309008 306128
rect 313372 306076 313424 306128
rect 314476 306076 314528 306128
rect 314660 306076 314712 306128
rect 315120 306076 315172 306128
rect 318892 306076 318944 306128
rect 319996 306076 320048 306128
rect 320272 306076 320324 306128
rect 320640 306076 320692 306128
rect 321560 306076 321612 306128
rect 322296 306076 322348 306128
rect 328644 306076 328696 306128
rect 329196 306076 329248 306128
rect 341064 306076 341116 306128
rect 341432 306076 341484 306128
rect 345204 306076 345256 306128
rect 346216 306076 346268 306128
rect 354772 306076 354824 306128
rect 371424 306076 371476 306128
rect 216312 306008 216364 306060
rect 292948 306008 293000 306060
rect 320456 306008 320508 306060
rect 321008 306008 321060 306060
rect 343916 306008 343968 306060
rect 354956 306008 355008 306060
rect 371700 306008 371752 306060
rect 213644 305940 213696 305992
rect 294052 305940 294104 305992
rect 305000 305940 305052 305992
rect 306104 305940 306156 305992
rect 306840 305940 306892 305992
rect 307668 305940 307720 305992
rect 320272 305940 320324 305992
rect 321376 305940 321428 305992
rect 327356 305940 327408 305992
rect 327816 305940 327868 305992
rect 341064 305940 341116 305992
rect 341984 305940 342036 305992
rect 216588 305872 216640 305924
rect 298468 305872 298520 305924
rect 327448 305872 327500 305924
rect 327724 305872 327776 305924
rect 170404 305804 170456 305856
rect 253940 305804 253992 305856
rect 254032 305804 254084 305856
rect 254216 305804 254268 305856
rect 255688 305804 255740 305856
rect 255872 305804 255924 305856
rect 257160 305804 257212 305856
rect 257436 305804 257488 305856
rect 258080 305804 258132 305856
rect 258356 305804 258408 305856
rect 258448 305804 258500 305856
rect 259184 305804 259236 305856
rect 262588 305804 262640 305856
rect 263324 305804 263376 305856
rect 263600 305804 263652 305856
rect 263784 305804 263836 305856
rect 264060 305804 264112 305856
rect 264888 305804 264940 305856
rect 265072 305804 265124 305856
rect 265256 305804 265308 305856
rect 266728 305804 266780 305856
rect 267556 305804 267608 305856
rect 269120 305804 269172 305856
rect 269488 305804 269540 305856
rect 269580 305804 269632 305856
rect 270040 305804 270092 305856
rect 270592 305804 270644 305856
rect 271052 305804 271104 305856
rect 272248 305804 272300 305856
rect 273076 305804 273128 305856
rect 273352 305804 273404 305856
rect 274272 305804 274324 305856
rect 274640 305804 274692 305856
rect 275744 305804 275796 305856
rect 276296 305804 276348 305856
rect 276848 305804 276900 305856
rect 277492 305804 277544 305856
rect 277860 305804 277912 305856
rect 279240 305804 279292 305856
rect 279976 305804 280028 305856
rect 280436 305804 280488 305856
rect 281080 305804 281132 305856
rect 281816 305804 281868 305856
rect 282276 305804 282328 305856
rect 293040 305804 293092 305856
rect 293684 305804 293736 305856
rect 306380 305804 306432 305856
rect 306932 305804 306984 305856
rect 354680 305940 354732 305992
rect 371516 305940 371568 305992
rect 352288 305872 352340 305924
rect 370320 305872 370372 305924
rect 344100 305804 344152 305856
rect 350816 305804 350868 305856
rect 360292 305804 360344 305856
rect 360568 305804 360620 305856
rect 361212 305804 361264 305856
rect 210976 305736 211028 305788
rect 195980 305668 196032 305720
rect 284852 305668 284904 305720
rect 292948 305736 293000 305788
rect 293868 305736 293920 305788
rect 342260 305736 342312 305788
rect 343088 305736 343140 305788
rect 353392 305736 353444 305788
rect 371608 305736 371660 305788
rect 295892 305668 295944 305720
rect 306380 305668 306432 305720
rect 307208 305668 307260 305720
rect 347136 305668 347188 305720
rect 364984 305668 365036 305720
rect 178040 305600 178092 305652
rect 275836 305600 275888 305652
rect 276296 305600 276348 305652
rect 277124 305600 277176 305652
rect 277492 305600 277544 305652
rect 278412 305600 278464 305652
rect 278872 305600 278924 305652
rect 279608 305600 279660 305652
rect 280252 305600 280304 305652
rect 280896 305600 280948 305652
rect 281724 305600 281776 305652
rect 282828 305600 282880 305652
rect 353300 305600 353352 305652
rect 371792 305600 371844 305652
rect 219072 305532 219124 305584
rect 291292 305532 291344 305584
rect 353576 305532 353628 305584
rect 368940 305532 368992 305584
rect 218888 305464 218940 305516
rect 289820 305464 289872 305516
rect 356152 305464 356204 305516
rect 367744 305464 367796 305516
rect 171692 305396 171744 305448
rect 234988 305396 235040 305448
rect 251364 305396 251416 305448
rect 251640 305396 251692 305448
rect 253020 305396 253072 305448
rect 253848 305396 253900 305448
rect 254032 305396 254084 305448
rect 254768 305396 254820 305448
rect 255688 305396 255740 305448
rect 256332 305396 256384 305448
rect 257160 305396 257212 305448
rect 257988 305396 258040 305448
rect 260840 305396 260892 305448
rect 261300 305396 261352 305448
rect 263784 305396 263836 305448
rect 264520 305396 264572 305448
rect 265072 305396 265124 305448
rect 265624 305396 265676 305448
rect 269672 305396 269724 305448
rect 270224 305396 270276 305448
rect 270776 305396 270828 305448
rect 271420 305396 271472 305448
rect 276204 305396 276256 305448
rect 277308 305396 277360 305448
rect 280160 305396 280212 305448
rect 280528 305396 280580 305448
rect 350908 305396 350960 305448
rect 362040 305396 362092 305448
rect 255504 305328 255556 305380
rect 256516 305328 256568 305380
rect 261116 305328 261168 305380
rect 262036 305328 262088 305380
rect 269304 305328 269356 305380
rect 270408 305328 270460 305380
rect 270592 305328 270644 305380
rect 271788 305328 271840 305380
rect 275836 305328 275888 305380
rect 281540 305328 281592 305380
rect 360292 305328 360344 305380
rect 368848 305328 368900 305380
rect 260840 305260 260892 305312
rect 261852 305260 261904 305312
rect 360200 305260 360252 305312
rect 368756 305260 368808 305312
rect 97264 305056 97316 305108
rect 97540 305056 97592 305108
rect 97540 304920 97592 304972
rect 97908 304920 97960 304972
rect 172336 304920 172388 304972
rect 245200 304920 245252 304972
rect 314660 304648 314712 304700
rect 315672 304648 315724 304700
rect 170036 304580 170088 304632
rect 240048 304580 240100 304632
rect 171968 304512 172020 304564
rect 245476 304512 245528 304564
rect 172244 304444 172296 304496
rect 248880 304444 248932 304496
rect 207020 304376 207072 304428
rect 285772 304376 285824 304428
rect 326436 304376 326488 304428
rect 452660 304376 452712 304428
rect 171784 304308 171836 304360
rect 256700 304308 256752 304360
rect 256884 304308 256936 304360
rect 257068 304308 257120 304360
rect 263508 304308 263560 304360
rect 263692 304308 263744 304360
rect 331772 304308 331824 304360
rect 485044 304308 485096 304360
rect 189080 304240 189132 304292
rect 283012 304240 283064 304292
rect 335912 304240 335964 304292
rect 514024 304240 514076 304292
rect 256608 304172 256660 304224
rect 256976 304172 257028 304224
rect 274824 303968 274876 304020
rect 275928 303968 275980 304020
rect 302516 303968 302568 304020
rect 303436 303968 303488 304020
rect 300952 303696 301004 303748
rect 301872 303696 301924 303748
rect 342444 303696 342496 303748
rect 343364 303696 343416 303748
rect 214656 303560 214708 303612
rect 288440 303560 288492 303612
rect 344008 303560 344060 303612
rect 344468 303560 344520 303612
rect 356060 303560 356112 303612
rect 373448 303560 373500 303612
rect 215944 303492 215996 303544
rect 290832 303492 290884 303544
rect 316132 303492 316184 303544
rect 316960 303492 317012 303544
rect 350724 303492 350776 303544
rect 370688 303492 370740 303544
rect 169944 303424 169996 303476
rect 246028 303424 246080 303476
rect 352012 303424 352064 303476
rect 372988 303424 373040 303476
rect 217968 303356 218020 303408
rect 293224 303356 293276 303408
rect 352104 303356 352156 303408
rect 373080 303356 373132 303408
rect 214748 303288 214800 303340
rect 289912 303288 289964 303340
rect 348700 303288 348752 303340
rect 370228 303288 370280 303340
rect 216036 303220 216088 303272
rect 291200 303220 291252 303272
rect 350632 303220 350684 303272
rect 372896 303220 372948 303272
rect 215024 303152 215076 303204
rect 291384 303152 291436 303204
rect 349620 303152 349672 303204
rect 373172 303152 373224 303204
rect 214564 303084 214616 303136
rect 292580 303084 292632 303136
rect 347964 303084 348016 303136
rect 372068 303084 372120 303136
rect 219164 303016 219216 303068
rect 299020 303016 299072 303068
rect 348884 303016 348936 303068
rect 373356 303016 373408 303068
rect 169760 302948 169812 303000
rect 251548 302948 251600 303000
rect 301228 302948 301280 303000
rect 363604 302948 363656 303000
rect 212172 302880 212224 302932
rect 294512 302880 294564 302932
rect 299388 302880 299440 302932
rect 365168 302880 365220 302932
rect 215116 302812 215168 302864
rect 288624 302812 288676 302864
rect 303712 302812 303764 302864
rect 304540 302812 304592 302864
rect 327172 302812 327224 302864
rect 327908 302812 327960 302864
rect 349436 302812 349488 302864
rect 366548 302812 366600 302864
rect 215852 302744 215904 302796
rect 288808 302744 288860 302796
rect 352564 302744 352616 302796
rect 369124 302744 369176 302796
rect 216496 302676 216548 302728
rect 289176 302676 289228 302728
rect 350172 302676 350224 302728
rect 363696 302676 363748 302728
rect 247684 302608 247736 302660
rect 247960 302608 248012 302660
rect 329932 302608 329984 302660
rect 330300 302608 330352 302660
rect 297180 302472 297232 302524
rect 297916 302472 297968 302524
rect 345112 302336 345164 302388
rect 345848 302336 345900 302388
rect 262312 302268 262364 302320
rect 262772 302200 262824 302252
rect 172428 302132 172480 302184
rect 240416 302132 240468 302184
rect 216220 302064 216272 302116
rect 293132 302064 293184 302116
rect 216128 301996 216180 302048
rect 296812 301996 296864 302048
rect 212448 301928 212500 301980
rect 296536 301928 296588 301980
rect 212264 301860 212316 301912
rect 296720 301860 296772 301912
rect 211068 301792 211120 301844
rect 295524 301792 295576 301844
rect 210792 301724 210844 301776
rect 295432 301724 295484 301776
rect 312268 301724 312320 301776
rect 374092 301724 374144 301776
rect 218428 301656 218480 301708
rect 349804 301656 349856 301708
rect 211712 301588 211764 301640
rect 347964 301588 348016 301640
rect 210884 301520 210936 301572
rect 295616 301520 295668 301572
rect 331588 301520 331640 301572
rect 494060 301520 494112 301572
rect 193220 301452 193272 301504
rect 282920 301452 282972 301504
rect 338672 301452 338724 301504
rect 529940 301452 529992 301504
rect 97356 300772 97408 300824
rect 249892 300772 249944 300824
rect 98644 300704 98696 300756
rect 251364 300704 251416 300756
rect 97724 300636 97776 300688
rect 246212 300636 246264 300688
rect 97816 300568 97868 300620
rect 242808 300568 242860 300620
rect 296996 300568 297048 300620
rect 297364 300568 297416 300620
rect 99104 300500 99156 300552
rect 243084 300500 243136 300552
rect 97632 300432 97684 300484
rect 242716 300432 242768 300484
rect 300216 300432 300268 300484
rect 362316 300432 362368 300484
rect 99380 300364 99432 300416
rect 240324 300364 240376 300416
rect 313832 300364 313884 300416
rect 376760 300364 376812 300416
rect 99564 300296 99616 300348
rect 240140 300296 240192 300348
rect 301228 300296 301280 300348
rect 370596 300296 370648 300348
rect 99840 300228 99892 300280
rect 238944 300228 238996 300280
rect 327632 300228 327684 300280
rect 463700 300228 463752 300280
rect 99196 300160 99248 300212
rect 237748 300160 237800 300212
rect 333152 300160 333204 300212
rect 498292 300160 498344 300212
rect 99472 300092 99524 300144
rect 236184 300092 236236 300144
rect 339960 300092 340012 300144
rect 538864 300092 538916 300144
rect 210608 300024 210660 300076
rect 347872 300024 347924 300076
rect 99012 299956 99064 300008
rect 233332 299956 233384 300008
rect 217784 299888 217836 299940
rect 348976 299888 349028 299940
rect 305552 299684 305604 299736
rect 305920 299684 305972 299736
rect 98828 299412 98880 299464
rect 247316 299412 247368 299464
rect 97908 299344 97960 299396
rect 242992 299344 243044 299396
rect 99748 299276 99800 299328
rect 240232 299276 240284 299328
rect 98920 299208 98972 299260
rect 238024 299208 238076 299260
rect 114836 299140 114888 299192
rect 244464 299140 244516 299192
rect 119988 299072 120040 299124
rect 247132 299072 247184 299124
rect 130292 299004 130344 299056
rect 249984 299004 250036 299056
rect 313648 299004 313700 299056
rect 378140 299004 378192 299056
rect 125140 298936 125192 298988
rect 238852 298936 238904 298988
rect 315120 298936 315172 298988
rect 381544 298936 381596 298988
rect 140596 298868 140648 298920
rect 250628 298868 250680 298920
rect 333060 298868 333112 298920
rect 500224 298868 500276 298920
rect 143448 298800 143500 298852
rect 248512 298800 248564 298852
rect 341432 298800 341484 298852
rect 547972 298800 548024 298852
rect 133788 298732 133840 298784
rect 243176 298732 243228 298784
rect 344836 298732 344888 298784
rect 567844 298732 567896 298784
rect 156052 298664 156104 298716
rect 251732 298664 251784 298716
rect 161204 298596 161256 298648
rect 247776 298596 247828 298648
rect 163780 298528 163832 298580
rect 234712 298528 234764 298580
rect 107108 298052 107160 298104
rect 111156 298052 111208 298104
rect 166356 298052 166408 298104
rect 170588 298052 170640 298104
rect 117412 297984 117464 298036
rect 133788 297984 133840 298036
rect 158628 297984 158680 298036
rect 169852 297984 169904 298036
rect 122564 297916 122616 297968
rect 237656 297916 237708 297968
rect 138020 297848 138072 297900
rect 239036 297848 239088 297900
rect 127716 297780 127768 297832
rect 143448 297780 143500 297832
rect 148324 297780 148376 297832
rect 236368 297780 236420 297832
rect 100024 297712 100076 297764
rect 169944 297712 169996 297764
rect 213460 297712 213512 297764
rect 293040 297712 293092 297764
rect 109684 297644 109736 297696
rect 135444 297576 135496 297628
rect 214472 297644 214524 297696
rect 294144 297644 294196 297696
rect 322204 297644 322256 297696
rect 381636 297644 381688 297696
rect 143172 297508 143224 297560
rect 172244 297576 172296 297628
rect 213828 297576 213880 297628
rect 294420 297576 294472 297628
rect 319260 297576 319312 297628
rect 412640 297576 412692 297628
rect 150900 297440 150952 297492
rect 171968 297508 172020 297560
rect 213184 297508 213236 297560
rect 346584 297508 346636 297560
rect 213736 297440 213788 297492
rect 294696 297440 294748 297492
rect 342812 297440 342864 297492
rect 556160 297440 556212 297492
rect 171692 297372 171744 297424
rect 210700 297372 210752 297424
rect 292948 297372 293000 297424
rect 342720 297372 342772 297424
rect 557540 297372 557592 297424
rect 170036 297304 170088 297356
rect 212356 297304 212408 297356
rect 291660 297304 291712 297356
rect 217876 297236 217928 297288
rect 295800 297236 295852 297288
rect 218796 297168 218848 297220
rect 294236 297168 294288 297220
rect 112260 297100 112312 297152
rect 235908 297100 235960 297152
rect 132868 297032 132920 297084
rect 251456 297032 251508 297084
rect 98736 296624 98788 296676
rect 240508 296624 240560 296676
rect 103520 296556 103572 296608
rect 234804 296556 234856 296608
rect 111156 296488 111208 296540
rect 236460 296488 236512 296540
rect 153200 296420 153252 296472
rect 248696 296420 248748 296472
rect 312176 296216 312228 296268
rect 372620 296216 372672 296268
rect 322020 296148 322072 296200
rect 421564 296148 421616 296200
rect 209780 296080 209832 296132
rect 285680 296080 285732 296132
rect 320732 296080 320784 296132
rect 422300 296080 422352 296132
rect 129740 296012 129792 296064
rect 273812 296012 273864 296064
rect 335820 296012 335872 296064
rect 516784 296012 516836 296064
rect 125600 295944 125652 295996
rect 272432 295944 272484 295996
rect 344100 295944 344152 295996
rect 563704 295944 563756 295996
rect 219348 295128 219400 295180
rect 295708 295128 295760 295180
rect 209688 295060 209740 295112
rect 287428 295060 287480 295112
rect 214932 294992 214984 295044
rect 294328 294992 294380 295044
rect 215760 294924 215812 294976
rect 296996 294924 297048 294976
rect 214380 294856 214432 294908
rect 297088 294856 297140 294908
rect 213276 294788 213328 294840
rect 296904 294788 296956 294840
rect 168380 294720 168432 294772
rect 278780 294720 278832 294772
rect 315028 294720 315080 294772
rect 387064 294720 387116 294772
rect 135260 294652 135312 294704
rect 274732 294652 274784 294704
rect 326068 294652 326120 294704
rect 457444 294652 457496 294704
rect 43444 294584 43496 294636
rect 258632 294584 258684 294636
rect 337200 294584 337252 294636
rect 525800 294584 525852 294636
rect 202880 293360 202932 293412
rect 284668 293360 284720 293412
rect 329104 293360 329156 293412
rect 467104 293360 467156 293412
rect 58624 293292 58676 293344
rect 260840 293292 260892 293344
rect 335728 293292 335780 293344
rect 509884 293292 509936 293344
rect 13084 293224 13136 293276
rect 254308 293224 254360 293276
rect 338580 293224 338632 293276
rect 527824 293224 527876 293276
rect 161480 292000 161532 292052
rect 279148 292000 279200 292052
rect 128360 291932 128412 291984
rect 271144 291932 271196 291984
rect 71044 291864 71096 291916
rect 263600 291864 263652 291916
rect 317788 291864 317840 291916
rect 405740 291864 405792 291916
rect 27620 291796 27672 291848
rect 257436 291796 257488 291848
rect 338488 291796 338540 291848
rect 534724 291796 534776 291848
rect 187700 290640 187752 290692
rect 283288 290640 283340 290692
rect 317696 290640 317748 290692
rect 408500 290640 408552 290692
rect 143540 290572 143592 290624
rect 274640 290572 274692 290624
rect 320640 290572 320692 290624
rect 418160 290572 418212 290624
rect 57244 290504 57296 290556
rect 261300 290504 261352 290556
rect 341340 290504 341392 290556
rect 543004 290504 543056 290556
rect 8300 290436 8352 290488
rect 254216 290436 254268 290488
rect 341248 290436 341300 290488
rect 549904 290436 549956 290488
rect 205640 289280 205692 289332
rect 286048 289280 286100 289332
rect 132500 289212 132552 289264
rect 273628 289212 273680 289264
rect 321928 289212 321980 289264
rect 430580 289212 430632 289264
rect 103520 289144 103572 289196
rect 269764 289144 269816 289196
rect 331496 289144 331548 289196
rect 490012 289144 490064 289196
rect 9680 289076 9732 289128
rect 254124 289076 254176 289128
rect 341156 289076 341208 289128
rect 552664 289076 552716 289128
rect 313556 287920 313608 287972
rect 382280 287920 382332 287972
rect 181444 287852 181496 287904
rect 281908 287852 281960 287904
rect 327540 287852 327592 287904
rect 460204 287852 460256 287904
rect 217692 287784 217744 287836
rect 351184 287784 351236 287836
rect 139400 287716 139452 287768
rect 275100 287716 275152 287768
rect 337108 287716 337160 287768
rect 518164 287716 518216 287768
rect 22100 287648 22152 287700
rect 255688 287648 255740 287700
rect 342628 287648 342680 287700
rect 561680 287648 561732 287700
rect 203524 286560 203576 286612
rect 283196 286560 283248 286612
rect 146300 286492 146352 286544
rect 276572 286492 276624 286544
rect 46940 286424 46992 286476
rect 259828 286424 259880 286476
rect 325976 286424 326028 286476
rect 454684 286424 454736 286476
rect 40040 286356 40092 286408
rect 258448 286356 258500 286408
rect 327448 286356 327500 286408
rect 458824 286356 458876 286408
rect 18604 286288 18656 286340
rect 252928 286288 252980 286340
rect 344008 286288 344060 286340
rect 566464 286288 566516 286340
rect 150440 285132 150492 285184
rect 276480 285132 276532 285184
rect 81440 285064 81492 285116
rect 265532 285064 265584 285116
rect 311992 285064 312044 285116
rect 371884 285064 371936 285116
rect 26240 284996 26292 285048
rect 257068 284996 257120 285048
rect 329012 284996 329064 285048
rect 471244 284996 471296 285048
rect 2780 284928 2832 284980
rect 252836 284928 252888 284980
rect 345480 284928 345532 284980
rect 575480 284928 575532 284980
rect 211160 283772 211212 283824
rect 285864 283772 285916 283824
rect 314936 283772 314988 283824
rect 390560 283772 390612 283824
rect 153200 283704 153252 283756
rect 277860 283704 277912 283756
rect 324872 283704 324924 283756
rect 442264 283704 442316 283756
rect 138020 283636 138072 283688
rect 275008 283636 275060 283688
rect 337016 283636 337068 283688
rect 522304 283636 522356 283688
rect 16580 283568 16632 283620
rect 255596 283568 255648 283620
rect 338396 283568 338448 283620
rect 531320 283568 531372 283620
rect 157340 282344 157392 282396
rect 277768 282344 277820 282396
rect 313464 282344 313516 282396
rect 374644 282344 374696 282396
rect 131120 282276 131172 282328
rect 273536 282276 273588 282328
rect 319168 282276 319220 282328
rect 414664 282276 414716 282328
rect 114560 282208 114612 282260
rect 270960 282208 271012 282260
rect 327356 282208 327408 282260
rect 464344 282208 464396 282260
rect 44180 282140 44232 282192
rect 259736 282140 259788 282192
rect 342536 282140 342588 282192
rect 556252 282140 556304 282192
rect 198740 280984 198792 281036
rect 284576 280984 284628 281036
rect 126980 280916 127032 280968
rect 272248 280916 272300 280968
rect 107660 280848 107712 280900
rect 269580 280848 269632 280900
rect 320548 280848 320600 280900
rect 417424 280848 417476 280900
rect 34520 280780 34572 280832
rect 258356 280780 258408 280832
rect 345388 280780 345440 280832
rect 571984 280780 572036 280832
rect 165620 279624 165672 279676
rect 279056 279624 279108 279676
rect 98000 279556 98052 279608
rect 268200 279556 268252 279608
rect 317604 279556 317656 279608
rect 407120 279556 407172 279608
rect 71780 279488 71832 279540
rect 264152 279488 264204 279540
rect 320456 279488 320508 279540
rect 423680 279488 423732 279540
rect 38660 279420 38712 279472
rect 257344 279420 257396 279472
rect 332968 279420 333020 279472
rect 493324 279420 493376 279472
rect 188344 278264 188396 278316
rect 281816 278264 281868 278316
rect 147680 278196 147732 278248
rect 276388 278196 276440 278248
rect 102140 278128 102192 278180
rect 269488 278128 269540 278180
rect 319076 278128 319128 278180
rect 409880 278128 409932 278180
rect 78680 278060 78732 278112
rect 265440 278060 265492 278112
rect 321836 278060 321888 278112
rect 428464 278060 428516 278112
rect 35900 277992 35952 278044
rect 258264 277992 258316 278044
rect 341064 277992 341116 278044
rect 553400 277992 553452 278044
rect 196624 276836 196676 276888
rect 281724 276836 281776 276888
rect 136640 276768 136692 276820
rect 274916 276768 274968 276820
rect 325884 276768 325936 276820
rect 445024 276768 445076 276820
rect 111800 276700 111852 276752
rect 270868 276700 270920 276752
rect 324780 276700 324832 276752
rect 448520 276700 448572 276752
rect 27712 276632 27764 276684
rect 256976 276632 257028 276684
rect 335636 276632 335688 276684
rect 511264 276632 511316 276684
rect 193312 275544 193364 275596
rect 283104 275544 283156 275596
rect 127072 275476 127124 275528
rect 273444 275476 273496 275528
rect 317512 275476 317564 275528
rect 404360 275476 404412 275528
rect 115940 275408 115992 275460
rect 270776 275408 270828 275460
rect 324688 275408 324740 275460
rect 448612 275408 448664 275460
rect 96620 275340 96672 275392
rect 268108 275340 268160 275392
rect 328920 275340 328972 275392
rect 468484 275340 468536 275392
rect 42800 275272 42852 275324
rect 250536 275272 250588 275324
rect 336924 275272 336976 275324
rect 525064 275272 525116 275324
rect 197360 274184 197412 274236
rect 284484 274184 284536 274236
rect 162860 274116 162912 274168
rect 278964 274116 279016 274168
rect 324596 274116 324648 274168
rect 446404 274116 446456 274168
rect 113180 274048 113232 274100
rect 270684 274048 270736 274100
rect 327264 274048 327316 274100
rect 460940 274048 460992 274100
rect 93860 273980 93912 274032
rect 268016 273980 268068 274032
rect 325792 273980 325844 274032
rect 459560 273980 459612 274032
rect 14464 273912 14516 273964
rect 254032 273912 254084 273964
rect 338304 273912 338356 273964
rect 531412 273912 531464 273964
rect 201500 272756 201552 272808
rect 284392 272756 284444 272808
rect 180800 272688 180852 272740
rect 281632 272688 281684 272740
rect 99380 272620 99432 272672
rect 260104 272620 260156 272672
rect 84200 272552 84252 272604
rect 265348 272552 265400 272604
rect 53840 272484 53892 272536
rect 261208 272484 261260 272536
rect 328828 272484 328880 272536
rect 475384 272484 475436 272536
rect 211804 271328 211856 271380
rect 286232 271328 286284 271380
rect 167000 271260 167052 271312
rect 278872 271260 278924 271312
rect 102232 271192 102284 271244
rect 269396 271192 269448 271244
rect 314844 271192 314896 271244
rect 386420 271192 386472 271244
rect 57980 271124 58032 271176
rect 261116 271124 261168 271176
rect 335544 271124 335596 271176
rect 517520 271124 517572 271176
rect 151820 269968 151872 270020
rect 276296 269968 276348 270020
rect 318064 269968 318116 270020
rect 400220 269968 400272 270020
rect 110420 269900 110472 269952
rect 269304 269900 269356 269952
rect 320364 269900 320416 269952
rect 420920 269900 420972 269952
rect 93952 269832 94004 269884
rect 267924 269832 267976 269884
rect 331404 269832 331456 269884
rect 486424 269832 486476 269884
rect 75920 269764 75972 269816
rect 264060 269764 264112 269816
rect 340972 269764 341024 269816
rect 552020 269764 552072 269816
rect 151912 268472 151964 268524
rect 276204 268472 276256 268524
rect 143632 268404 143684 268456
rect 274824 268404 274876 268456
rect 328644 268404 328696 268456
rect 473452 268404 473504 268456
rect 77300 268336 77352 268388
rect 265256 268336 265308 268388
rect 328736 268336 328788 268388
rect 474740 268336 474792 268388
rect 2964 267656 3016 267708
rect 225604 267656 225656 267708
rect 317420 267248 317472 267300
rect 407212 267248 407264 267300
rect 217324 267180 217376 267232
rect 351092 267180 351144 267232
rect 332876 267112 332928 267164
rect 495440 267112 495492 267164
rect 340880 267044 340932 267096
rect 549260 267044 549312 267096
rect 70400 266976 70452 267028
rect 263968 266976 264020 267028
rect 343916 266976 343968 267028
rect 565820 266976 565872 267028
rect 191840 265888 191892 265940
rect 283472 265888 283524 265940
rect 133880 265820 133932 265872
rect 273352 265820 273404 265872
rect 313372 265820 313424 265872
rect 382372 265820 382424 265872
rect 121460 265752 121512 265804
rect 272156 265752 272208 265804
rect 331312 265752 331364 265804
rect 491300 265752 491352 265804
rect 39304 265684 39356 265736
rect 258172 265684 258224 265736
rect 338212 265684 338264 265736
rect 535460 265684 535512 265736
rect 11060 265616 11112 265668
rect 247684 265616 247736 265668
rect 342444 265616 342496 265668
rect 560944 265616 560996 265668
rect 314752 264392 314804 264444
rect 389180 264392 389232 264444
rect 154580 264324 154632 264376
rect 277676 264324 277728 264376
rect 323492 264324 323544 264376
rect 440240 264324 440292 264376
rect 149060 264256 149112 264308
rect 276112 264256 276164 264308
rect 323584 264256 323636 264308
rect 443000 264256 443052 264308
rect 69020 264188 69072 264240
rect 263876 264188 263928 264240
rect 345296 264188 345348 264240
rect 574100 264188 574152 264240
rect 316592 263100 316644 263152
rect 393320 263100 393372 263152
rect 316500 263032 316552 263084
rect 397460 263032 397512 263084
rect 142160 262964 142212 263016
rect 275284 262964 275336 263016
rect 323308 262964 323360 263016
rect 436100 262964 436152 263016
rect 52460 262896 52512 262948
rect 261024 262896 261076 262948
rect 323400 262896 323452 262948
rect 441620 262896 441672 262948
rect 7564 262828 7616 262880
rect 252744 262828 252796 262880
rect 324504 262828 324556 262880
rect 449900 262828 449952 262880
rect 314660 261808 314712 261860
rect 390652 261808 390704 261860
rect 212540 261740 212592 261792
rect 287336 261740 287388 261792
rect 316408 261740 316460 261792
rect 398840 261740 398892 261792
rect 158720 261672 158772 261724
rect 277584 261672 277636 261724
rect 323216 261672 323268 261724
rect 438860 261672 438912 261724
rect 144920 261604 144972 261656
rect 276020 261604 276072 261656
rect 334624 261604 334676 261656
rect 506480 261604 506532 261656
rect 73160 261536 73212 261588
rect 263784 261536 263836 261588
rect 334532 261536 334584 261588
rect 510620 261536 510672 261588
rect 13820 261468 13872 261520
rect 254400 261468 254452 261520
rect 343824 261468 343876 261520
rect 569960 261468 570012 261520
rect 124220 260380 124272 260432
rect 251916 260380 251968 260432
rect 63500 260312 63552 260364
rect 262680 260312 262732 260364
rect 316224 260312 316276 260364
rect 391940 260312 391992 260364
rect 39396 260244 39448 260296
rect 256884 260244 256936 260296
rect 316316 260244 316368 260296
rect 396080 260244 396132 260296
rect 30380 260176 30432 260228
rect 257252 260176 257304 260228
rect 339868 260176 339920 260228
rect 542360 260176 542412 260228
rect 19340 260108 19392 260160
rect 246304 260108 246356 260160
rect 342352 260108 342404 260160
rect 558920 260108 558972 260160
rect 362224 259360 362276 259412
rect 579804 259360 579856 259412
rect 176660 258816 176712 258868
rect 267004 258816 267056 258868
rect 323124 258816 323176 258868
rect 434720 258816 434772 258868
rect 217600 258748 217652 258800
rect 346492 258748 346544 258800
rect 173900 258680 173952 258732
rect 280620 258680 280672 258732
rect 339776 258680 339828 258732
rect 539692 258680 539744 258732
rect 218612 257592 218664 257644
rect 287244 257592 287296 257644
rect 117320 257524 117372 257576
rect 251824 257524 251876 257576
rect 106280 257456 106332 257508
rect 261484 257456 261536 257508
rect 334440 257456 334492 257508
rect 509240 257456 509292 257508
rect 25596 257388 25648 257440
rect 255412 257388 255464 257440
rect 339684 257388 339736 257440
rect 540980 257388 541032 257440
rect 23480 257320 23532 257372
rect 255504 257320 255556 257372
rect 339592 257320 339644 257372
rect 545120 257320 545172 257372
rect 318984 256368 319036 256420
rect 413284 256368 413336 256420
rect 217140 256300 217192 256352
rect 348424 256300 348476 256352
rect 122840 256232 122892 256284
rect 272064 256232 272116 256284
rect 320272 256232 320324 256284
rect 425060 256232 425112 256284
rect 118700 256164 118752 256216
rect 271972 256164 272024 256216
rect 321744 256164 321796 256216
rect 431960 256164 432012 256216
rect 92480 256096 92532 256148
rect 266728 256096 266780 256148
rect 323032 256096 323084 256148
rect 440332 256096 440384 256148
rect 77392 256028 77444 256080
rect 265164 256028 265216 256080
rect 325700 256028 325752 256080
rect 454040 256028 454092 256080
rect 17960 255960 18012 256012
rect 255872 255960 255924 256012
rect 334348 255960 334400 256012
rect 506572 255960 506624 256012
rect 169760 254872 169812 254924
rect 280528 254872 280580 254924
rect 217416 254804 217468 254856
rect 345204 254804 345256 254856
rect 3332 254736 3384 254788
rect 8944 254736 8996 254788
rect 95240 254736 95292 254788
rect 267832 254736 267884 254788
rect 316132 254736 316184 254788
rect 398932 254736 398984 254788
rect 91100 254668 91152 254720
rect 266544 254668 266596 254720
rect 324412 254668 324464 254720
rect 443644 254668 443696 254720
rect 88340 254600 88392 254652
rect 264244 254600 264296 254652
rect 343640 254600 343692 254652
rect 564532 254600 564584 254652
rect 86960 254532 87012 254584
rect 266636 254532 266688 254584
rect 343732 254532 343784 254584
rect 567200 254532 567252 254584
rect 302608 253784 302660 253836
rect 360292 253784 360344 253836
rect 304080 253716 304132 253768
rect 367192 253716 367244 253768
rect 301136 253648 301188 253700
rect 364524 253648 364576 253700
rect 301044 253580 301096 253632
rect 368480 253580 368532 253632
rect 176752 253512 176804 253564
rect 280436 253512 280488 253564
rect 316040 253512 316092 253564
rect 394700 253512 394752 253564
rect 218520 253444 218572 253496
rect 347780 253444 347832 253496
rect 118792 253376 118844 253428
rect 270592 253376 270644 253428
rect 322940 253376 322992 253428
rect 437480 253376 437532 253428
rect 110512 253308 110564 253360
rect 271052 253308 271104 253360
rect 332784 253308 332836 253360
rect 496084 253308 496136 253360
rect 85580 253240 85632 253292
rect 266452 253240 266504 253292
rect 332692 253240 332744 253292
rect 499580 253240 499632 253292
rect 80060 253172 80112 253224
rect 265072 253172 265124 253224
rect 336832 253172 336884 253224
rect 528560 253172 528612 253224
rect 172520 252084 172572 252136
rect 280344 252084 280396 252136
rect 321652 252084 321704 252136
rect 427820 252084 427872 252136
rect 160192 252016 160244 252068
rect 277492 252016 277544 252068
rect 321560 252016 321612 252068
rect 432052 252016 432104 252068
rect 155960 251948 156012 252000
rect 277400 251948 277452 252000
rect 327172 251948 327224 252000
rect 466460 251948 466512 252000
rect 49700 251880 49752 251932
rect 259644 251880 259696 251932
rect 339500 251880 339552 251932
rect 538220 251880 538272 251932
rect 46204 251812 46256 251864
rect 259552 251812 259604 251864
rect 345112 251812 345164 251864
rect 578240 251812 578292 251864
rect 309508 251132 309560 251184
rect 365812 251132 365864 251184
rect 306748 251064 306800 251116
rect 363236 251064 363288 251116
rect 306840 250996 306892 251048
rect 364616 250996 364668 251048
rect 306932 250928 306984 250980
rect 364708 250928 364760 250980
rect 305552 250860 305604 250912
rect 363328 250860 363380 250912
rect 209872 250792 209924 250844
rect 286140 250792 286192 250844
rect 311900 250792 311952 250844
rect 371240 250792 371292 250844
rect 135352 250724 135404 250776
rect 273720 250724 273772 250776
rect 303896 250724 303948 250776
rect 365904 250724 365956 250776
rect 60740 250656 60792 250708
rect 255964 250656 256016 250708
rect 318892 250656 318944 250708
rect 416780 250656 416832 250708
rect 67640 250588 67692 250640
rect 263692 250588 263744 250640
rect 330300 250588 330352 250640
rect 484400 250588 484452 250640
rect 66260 250520 66312 250572
rect 262588 250520 262640 250572
rect 334256 250520 334308 250572
rect 503720 250520 503772 250572
rect 52552 250452 52604 250504
rect 260932 250452 260984 250504
rect 345020 250452 345072 250504
rect 576860 250452 576912 250504
rect 309600 250384 309652 250436
rect 365720 250384 365772 250436
rect 305644 250316 305696 250368
rect 360200 250316 360252 250368
rect 318800 249432 318852 249484
rect 414020 249432 414072 249484
rect 185032 249364 185084 249416
rect 282184 249364 282236 249416
rect 340144 249364 340196 249416
rect 455420 249364 455472 249416
rect 217232 249296 217284 249348
rect 346400 249296 346452 249348
rect 82820 249228 82872 249280
rect 264980 249228 265032 249280
rect 327080 249228 327132 249280
rect 467840 249228 467892 249280
rect 74540 249160 74592 249212
rect 264336 249160 264388 249212
rect 328552 249160 328604 249212
rect 477500 249160 477552 249212
rect 62120 249092 62172 249144
rect 262496 249092 262548 249144
rect 334164 249092 334216 249144
rect 512000 249092 512052 249144
rect 57336 249024 57388 249076
rect 261392 249024 261444 249076
rect 335452 249024 335504 249076
rect 520280 249024 520332 249076
rect 306656 248344 306708 248396
rect 362960 248344 363012 248396
rect 302424 248276 302476 248328
rect 359464 248276 359516 248328
rect 306564 248208 306616 248260
rect 364432 248208 364484 248260
rect 305092 248140 305144 248192
rect 363052 248140 363104 248192
rect 305460 248072 305512 248124
rect 364340 248072 364392 248124
rect 201592 248004 201644 248056
rect 284760 248004 284812 248056
rect 302516 248004 302568 248056
rect 361948 248004 362000 248056
rect 140780 247936 140832 247988
rect 275192 247936 275244 247988
rect 302332 247936 302384 247988
rect 372712 247936 372764 247988
rect 89720 247868 89772 247920
rect 253204 247868 253256 247920
rect 320180 247868 320232 247920
rect 423772 247868 423824 247920
rect 41420 247800 41472 247852
rect 258540 247800 258592 247852
rect 332600 247800 332652 247852
rect 502340 247800 502392 247852
rect 35164 247732 35216 247784
rect 257160 247732 257212 247784
rect 333980 247732 334032 247784
rect 505100 247732 505152 247784
rect 4160 247664 4212 247716
rect 252652 247664 252704 247716
rect 334072 247664 334124 247716
rect 507860 247664 507912 247716
rect 308036 247596 308088 247648
rect 363144 247596 363196 247648
rect 303712 247528 303764 247580
rect 356704 247528 356756 247580
rect 355692 247460 355744 247512
rect 369860 247460 369912 247512
rect 211896 246780 211948 246832
rect 262312 246780 262364 246832
rect 175280 246712 175332 246764
rect 280252 246712 280304 246764
rect 120080 246644 120132 246696
rect 272340 246644 272392 246696
rect 328460 246644 328512 246696
rect 471980 246644 472032 246696
rect 104900 246576 104952 246628
rect 269212 246576 269264 246628
rect 330116 246576 330168 246628
rect 480260 246576 480312 246628
rect 85672 246508 85724 246560
rect 266820 246508 266872 246560
rect 330208 246508 330260 246560
rect 483020 246508 483072 246560
rect 64880 246440 64932 246492
rect 262404 246440 262456 246492
rect 330024 246440 330076 246492
rect 485780 246440 485832 246492
rect 48320 246372 48372 246424
rect 260012 246372 260064 246424
rect 331220 246372 331272 246424
rect 492680 246372 492732 246424
rect 6920 246304 6972 246356
rect 253020 246304 253072 246356
rect 335360 246304 335412 246356
rect 516140 246304 516192 246356
rect 355416 245556 355468 245608
rect 372804 245556 372856 245608
rect 307944 245488 307996 245540
rect 361580 245488 361632 245540
rect 307760 245420 307812 245472
rect 361764 245420 361816 245472
rect 307852 245352 307904 245404
rect 361856 245352 361908 245404
rect 198096 245284 198148 245336
rect 283380 245284 283432 245336
rect 306380 245284 306432 245336
rect 361672 245284 361724 245336
rect 171232 245216 171284 245268
rect 280712 245216 280764 245268
rect 302240 245216 302292 245268
rect 360936 245216 360988 245268
rect 168472 245148 168524 245200
rect 279240 245148 279292 245200
rect 324320 245148 324372 245200
rect 445760 245148 445812 245200
rect 109040 245080 109092 245132
rect 269672 245080 269724 245132
rect 329932 245080 329984 245132
rect 481732 245080 481784 245132
rect 100760 245012 100812 245064
rect 268292 245012 268344 245064
rect 329840 245012 329892 245064
rect 481640 245012 481692 245064
rect 60832 244944 60884 244996
rect 262772 244944 262824 244996
rect 338120 244944 338172 244996
rect 534080 244944 534132 244996
rect 31760 244876 31812 244928
rect 250444 244876 250496 244928
rect 342260 244876 342312 244928
rect 560300 244876 560352 244928
rect 355324 244808 355376 244860
rect 365996 244808 366048 244860
rect 355600 244740 355652 244792
rect 364800 244740 364852 244792
rect 355508 244604 355560 244656
rect 358176 244604 358228 244656
rect 356980 243924 357032 243976
rect 367928 243924 367980 243976
rect 299664 243856 299716 243908
rect 362408 243856 362460 243908
rect 299480 243788 299532 243840
rect 362224 243788 362276 243840
rect 298560 243720 298612 243772
rect 361028 243720 361080 243772
rect 300860 243652 300912 243704
rect 363788 243652 363840 243704
rect 219256 243584 219308 243636
rect 297180 243584 297232 243636
rect 300952 243584 301004 243636
rect 366088 243584 366140 243636
rect 217508 243516 217560 243568
rect 297272 243516 297324 243568
rect 299572 243516 299624 243568
rect 369308 243516 369360 243568
rect 356796 242156 356848 242208
rect 369216 242156 369268 242208
rect 577596 206932 577648 206984
rect 579620 206932 579672 206984
rect 3056 202784 3108 202836
rect 196716 202784 196768 202836
rect 214380 195644 214432 195696
rect 217324 195644 217376 195696
rect 215760 193128 215812 193180
rect 218704 193128 218756 193180
rect 3516 188980 3568 189032
rect 203616 188980 203668 189032
rect 210608 188980 210660 189032
rect 216680 188980 216732 189032
rect 374736 179324 374788 179376
rect 580172 179324 580224 179376
rect 371976 166948 372028 167000
rect 579620 166948 579672 167000
rect 213644 159604 213696 159656
rect 256700 159604 256752 159656
rect 214472 159536 214524 159588
rect 260840 159536 260892 159588
rect 322940 159536 322992 159588
rect 358084 159536 358136 159588
rect 217876 159468 217928 159520
rect 264980 159468 265032 159520
rect 320088 159468 320140 159520
rect 357992 159468 358044 159520
rect 212172 159400 212224 159452
rect 259460 159400 259512 159452
rect 314660 159400 314712 159452
rect 357900 159400 357952 159452
rect 214840 159332 214892 159384
rect 282920 159332 282972 159384
rect 310428 159332 310480 159384
rect 357716 159332 357768 159384
rect 300952 159264 301004 159316
rect 357808 159264 357860 159316
rect 279240 159196 279292 159248
rect 360752 159196 360804 159248
rect 278136 159128 278188 159180
rect 360660 159128 360712 159180
rect 275836 159060 275888 159112
rect 359280 159060 359332 159112
rect 277032 158992 277084 159044
rect 360844 158992 360896 159044
rect 274456 158924 274508 158976
rect 359372 158924 359424 158976
rect 267648 158856 267700 158908
rect 370504 158856 370556 158908
rect 262864 158788 262916 158840
rect 366364 158788 366416 158840
rect 211712 158720 211764 158772
rect 239588 158720 239640 158772
rect 258540 158720 258592 158772
rect 363696 158720 363748 158772
rect 213184 158652 213236 158704
rect 238116 158652 238168 158704
rect 308680 158652 308732 158704
rect 320088 158652 320140 158704
rect 211988 158584 212040 158636
rect 230480 158584 230532 158636
rect 306104 158584 306156 158636
rect 314660 158584 314712 158636
rect 215944 158516 215996 158568
rect 236000 158516 236052 158568
rect 259552 158516 259604 158568
rect 367836 158516 367888 158568
rect 213368 158448 213420 158500
rect 234712 158448 234764 158500
rect 265992 158448 266044 158500
rect 369124 158448 369176 158500
rect 219072 158380 219124 158432
rect 242992 158380 243044 158432
rect 268752 158380 268804 158432
rect 357440 158380 357492 158432
rect 216036 158312 216088 158364
rect 242900 158312 242952 158364
rect 270224 158312 270276 158364
rect 357624 158312 357676 158364
rect 216404 158244 216456 158296
rect 245660 158244 245712 158296
rect 271144 158244 271196 158296
rect 357532 158244 357584 158296
rect 214564 158176 214616 158228
rect 247040 158176 247092 158228
rect 298928 158176 298980 158228
rect 373448 158176 373500 158228
rect 217968 158108 218020 158160
rect 251180 158108 251232 158160
rect 303528 158108 303580 158160
rect 310428 158108 310480 158160
rect 321192 158108 321244 158160
rect 360384 158108 360436 158160
rect 216312 158040 216364 158092
rect 249800 158040 249852 158092
rect 313464 158040 313516 158092
rect 359004 158040 359056 158092
rect 218980 157972 219032 158024
rect 252560 157972 252612 158024
rect 315856 157972 315908 158024
rect 359096 157972 359148 158024
rect 214748 157904 214800 157956
rect 233240 157904 233292 157956
rect 318616 157904 318668 157956
rect 359188 157904 359240 157956
rect 218888 157836 218940 157888
rect 234620 157836 234672 157888
rect 272248 157836 272300 157888
rect 322940 157836 322992 157888
rect 323400 157836 323452 157888
rect 360476 157836 360528 157888
rect 215852 157768 215904 157820
rect 229100 157768 229152 157820
rect 325976 157768 326028 157820
rect 360568 157768 360620 157820
rect 240692 157700 240744 157752
rect 373356 157700 373408 157752
rect 256608 157632 256660 157684
rect 366548 157632 366600 157684
rect 261760 157360 261812 157412
rect 317052 157360 317104 157412
rect 250168 157292 250220 157344
rect 368848 157292 368900 157344
rect 248328 157224 248380 157276
rect 364984 157224 365036 157276
rect 257160 157156 257212 157208
rect 367652 157156 367704 157208
rect 255964 157088 256016 157140
rect 364892 157088 364944 157140
rect 258632 157020 258684 157072
rect 367560 157020 367612 157072
rect 260656 156952 260708 157004
rect 367468 156952 367520 157004
rect 276112 156884 276164 156936
rect 368940 156884 368992 156936
rect 281356 156816 281408 156868
rect 371792 156816 371844 156868
rect 286232 156748 286284 156800
rect 371700 156748 371752 156800
rect 273352 156680 273404 156732
rect 358820 156680 358872 156732
rect 291016 156612 291068 156664
rect 370412 156612 370464 156664
rect 296260 156544 296312 156596
rect 359556 156544 359608 156596
rect 317052 156476 317104 156528
rect 370688 156476 370740 156528
rect 311256 156408 311308 156460
rect 358912 156408 358964 156460
rect 245384 155864 245436 155916
rect 366180 155864 366232 155916
rect 212080 155796 212132 155848
rect 237380 155796 237432 155848
rect 253572 155796 253624 155848
rect 368664 155796 368716 155848
rect 213552 155728 213604 155780
rect 241520 155728 241572 155780
rect 252100 155728 252152 155780
rect 362040 155728 362092 155780
rect 216220 155660 216272 155712
rect 248420 155660 248472 155712
rect 261944 155660 261996 155712
rect 367376 155660 367428 155712
rect 210976 155592 211028 155644
rect 267832 155592 267884 155644
rect 268936 155592 268988 155644
rect 373080 155592 373132 155644
rect 213460 155524 213512 155576
rect 253940 155524 253992 155576
rect 266728 155524 266780 155576
rect 369952 155524 370004 155576
rect 210884 155456 210936 155508
rect 270500 155456 270552 155508
rect 271052 155456 271104 155508
rect 372988 155456 373040 155508
rect 210700 155388 210752 155440
rect 255320 155388 255372 155440
rect 265992 155388 266044 155440
rect 367284 155388 367336 155440
rect 218796 155320 218848 155372
rect 263600 155320 263652 155372
rect 264428 155320 264480 155372
rect 363512 155320 363564 155372
rect 212264 155252 212316 155304
rect 273260 155252 273312 155304
rect 274456 155252 274508 155304
rect 368756 155252 368808 155304
rect 213276 155184 213328 155236
rect 274640 155184 274692 155236
rect 278688 155184 278740 155236
rect 371608 155184 371660 155236
rect 217508 155116 217560 155168
rect 278780 155116 278832 155168
rect 284116 155116 284168 155168
rect 371516 155116 371568 155168
rect 219164 155048 219216 155100
rect 287060 155048 287112 155100
rect 288256 155048 288308 155100
rect 371424 155048 371476 155100
rect 216128 154980 216180 155032
rect 277400 154980 277452 155032
rect 293592 154980 293644 155032
rect 367744 154980 367796 155032
rect 253664 154504 253716 154556
rect 370228 154504 370280 154556
rect 263968 154436 264020 154488
rect 372896 154436 372948 154488
rect 299480 153960 299532 154012
rect 363604 153960 363656 154012
rect 295340 153892 295392 153944
rect 362224 153892 362276 153944
rect 288440 153824 288492 153876
rect 361028 153824 361080 153876
rect 345756 152532 345808 152584
rect 369216 152532 369268 152584
rect 300860 152464 300912 152516
rect 370596 152464 370648 152516
rect 3516 150356 3568 150408
rect 198004 150356 198056 150408
rect 3516 137912 3568 137964
rect 206284 137912 206336 137964
rect 3424 97928 3476 97980
rect 192484 97928 192536 97980
rect 3148 85484 3200 85536
rect 200764 85484 200816 85536
rect 3424 71680 3476 71732
rect 207664 71680 207716 71732
rect 373264 60664 373316 60716
rect 580172 60664 580224 60716
rect 3056 59304 3108 59356
rect 25504 59304 25556 59356
rect 3424 45500 3476 45552
rect 199384 45500 199436 45552
rect 3516 33056 3568 33108
rect 95884 33056 95936 33108
rect 577504 33056 577556 33108
rect 579620 33056 579672 33108
rect 3424 20612 3476 20664
rect 64144 20612 64196 20664
rect 160100 11704 160152 11756
rect 161296 11704 161348 11756
rect 176660 11704 176712 11756
rect 177856 11704 177908 11756
rect 184940 11704 184992 11756
rect 186136 11704 186188 11756
rect 234620 11704 234672 11756
rect 235816 11704 235868 11756
rect 242900 11704 242952 11756
rect 244096 11704 244148 11756
rect 316224 9256 316276 9308
rect 363420 9256 363472 9308
rect 319720 9188 319772 9240
rect 367192 9188 367244 9240
rect 312636 9120 312688 9172
rect 360292 9120 360344 9172
rect 305552 9052 305604 9104
rect 366088 9052 366140 9104
rect 303160 8984 303212 9036
rect 364524 8984 364576 9036
rect 304356 8916 304408 8968
rect 365996 8916 366048 8968
rect 330392 6808 330444 6860
rect 363328 6808 363380 6860
rect 326804 6740 326856 6792
rect 360200 6740 360252 6792
rect 315028 6672 315080 6724
rect 361948 6672 362000 6724
rect 313832 6604 313884 6656
rect 360936 6604 360988 6656
rect 318524 6536 318576 6588
rect 365904 6536 365956 6588
rect 317328 6468 317380 6520
rect 364800 6468 364852 6520
rect 311440 6400 311492 6452
rect 359464 6400 359516 6452
rect 310244 6332 310296 6384
rect 358176 6332 358228 6384
rect 307944 6264 307996 6316
rect 369860 6264 369912 6316
rect 306748 6196 306800 6248
rect 368480 6196 368532 6248
rect 309048 6128 309100 6180
rect 372712 6128 372764 6180
rect 333888 6060 333940 6112
rect 364708 6060 364760 6112
rect 337476 5992 337528 6044
rect 363236 5992 363288 6044
rect 340972 5924 341024 5976
rect 364616 5924 364668 5976
rect 180248 4088 180300 4140
rect 181444 4088 181496 4140
rect 208584 4088 208636 4140
rect 211804 4088 211856 4140
rect 212356 4088 212408 4140
rect 245200 4088 245252 4140
rect 336280 4088 336332 4140
rect 362960 4088 363012 4140
rect 460204 4088 460256 4140
rect 462780 4088 462832 4140
rect 468484 4088 468536 4140
rect 471060 4088 471112 4140
rect 51356 4020 51408 4072
rect 57244 4020 57296 4072
rect 213828 4020 213880 4072
rect 258264 4020 258316 4072
rect 332692 4020 332744 4072
rect 364340 4020 364392 4072
rect 213736 3952 213788 4004
rect 260656 3952 260708 4004
rect 329196 3952 329248 4004
rect 363052 3952 363104 4004
rect 219348 3884 219400 3936
rect 266544 3884 266596 3936
rect 322112 3884 322164 3936
rect 356704 3884 356756 3936
rect 371884 3884 371936 3936
rect 375288 3884 375340 3936
rect 4068 3816 4120 3868
rect 7564 3816 7616 3868
rect 214932 3816 214984 3868
rect 262956 3816 263008 3868
rect 298468 3816 298520 3868
rect 345756 3816 345808 3868
rect 516784 3816 516836 3868
rect 519544 3816 519596 3868
rect 566464 3816 566516 3868
rect 569132 3816 569184 3868
rect 69112 3748 69164 3800
rect 71044 3748 71096 3800
rect 135260 3748 135312 3800
rect 136456 3748 136508 3800
rect 195980 3748 196032 3800
rect 196624 3748 196676 3800
rect 218704 3748 218756 3800
rect 277124 3748 277176 3800
rect 300768 3748 300820 3800
rect 354128 3748 354180 3800
rect 355140 3748 355192 3800
rect 361580 3748 361632 3800
rect 30104 3680 30156 3732
rect 39396 3680 39448 3732
rect 44272 3680 44324 3732
rect 46204 3680 46256 3732
rect 46664 3680 46716 3732
rect 170496 3680 170548 3732
rect 211068 3680 211120 3732
rect 268844 3680 268896 3732
rect 292580 3680 292632 3732
rect 348424 3680 348476 3732
rect 352840 3680 352892 3732
rect 361028 3680 361080 3732
rect 489184 3680 489236 3732
rect 491116 3680 491168 3732
rect 6460 3612 6512 3664
rect 18604 3612 18656 3664
rect 25320 3612 25372 3664
rect 171784 3612 171836 3664
rect 183744 3612 183796 3664
rect 188344 3612 188396 3664
rect 209780 3612 209832 3664
rect 210976 3612 211028 3664
rect 217324 3612 217376 3664
rect 276020 3612 276072 3664
rect 290188 3612 290240 3664
rect 351184 3612 351236 3664
rect 354036 3612 354088 3664
rect 365260 3612 365312 3664
rect 1676 3544 1728 3596
rect 32404 3544 32456 3596
rect 33600 3544 33652 3596
rect 35164 3544 35216 3596
rect 38384 3544 38436 3596
rect 39304 3544 39356 3596
rect 52460 3544 52512 3596
rect 53380 3544 53432 3596
rect 56048 3544 56100 3596
rect 57336 3544 57388 3596
rect 59636 3544 59688 3596
rect 211896 3544 211948 3596
rect 212448 3544 212500 3596
rect 272432 3544 272484 3596
rect 285404 3544 285456 3596
rect 345664 3544 345716 3596
rect 349252 3544 349304 3596
rect 355140 3544 355192 3596
rect 355232 3544 355284 3596
rect 12348 3476 12400 3528
rect 13084 3476 13136 3528
rect 15936 3476 15988 3528
rect 170404 3476 170456 3528
rect 187332 3476 187384 3528
rect 195980 3476 196032 3528
rect 209688 3476 209740 3528
rect 218060 3476 218112 3528
rect 219164 3476 219216 3528
rect 280712 3476 280764 3528
rect 281908 3476 281960 3528
rect 353944 3476 353996 3528
rect 356336 3476 356388 3528
rect 358084 3476 358136 3528
rect 362316 3544 362368 3596
rect 371332 3612 371384 3664
rect 377404 3612 377456 3664
rect 411904 3612 411956 3664
rect 369400 3544 369452 3596
rect 372804 3544 372856 3596
rect 381544 3544 381596 3596
rect 384764 3544 384816 3596
rect 398840 3544 398892 3596
rect 400128 3544 400180 3596
rect 407212 3544 407264 3596
rect 408408 3544 408460 3596
rect 421564 3544 421616 3596
rect 427268 3544 427320 3596
rect 442264 3544 442316 3596
rect 445024 3544 445076 3596
rect 445116 3544 445168 3596
rect 458088 3544 458140 3596
rect 458824 3544 458876 3596
rect 465172 3544 465224 3596
rect 467104 3544 467156 3596
rect 469864 3544 469916 3596
rect 365720 3476 365772 3528
rect 381636 3476 381688 3528
rect 572 3408 624 3460
rect 171140 3408 171192 3460
rect 190828 3408 190880 3460
rect 203524 3408 203576 3460
rect 216588 3408 216640 3460
rect 284300 3408 284352 3460
rect 286600 3408 286652 3460
rect 367100 3408 367152 3460
rect 382372 3408 382424 3460
rect 383568 3408 383620 3460
rect 387064 3408 387116 3460
rect 388260 3408 388312 3460
rect 390560 3408 390612 3460
rect 391848 3408 391900 3460
rect 37188 3340 37240 3392
rect 43444 3340 43496 3392
rect 57244 3340 57296 3392
rect 58624 3340 58676 3392
rect 118700 3340 118752 3392
rect 119896 3340 119948 3392
rect 215024 3340 215076 3392
rect 240508 3340 240560 3392
rect 339868 3340 339920 3392
rect 364432 3340 364484 3392
rect 388444 3340 388496 3392
rect 215116 3272 215168 3324
rect 226340 3272 226392 3324
rect 338672 3272 338724 3324
rect 361672 3272 361724 3324
rect 414664 3408 414716 3460
rect 416688 3408 416740 3460
rect 423772 3476 423824 3528
rect 424968 3476 425020 3528
rect 429660 3476 429712 3528
rect 431960 3476 432012 3528
rect 433248 3476 433300 3528
rect 440332 3476 440384 3528
rect 441528 3476 441580 3528
rect 443644 3476 443696 3528
rect 447416 3476 447468 3528
rect 448520 3476 448572 3528
rect 449808 3476 449860 3528
rect 454684 3476 454736 3528
rect 456892 3476 456944 3528
rect 462964 3476 463016 3528
rect 471244 3476 471296 3528
rect 473452 3476 473504 3528
rect 475384 3544 475436 3596
rect 476948 3544 477000 3596
rect 500224 3544 500276 3596
rect 501788 3544 501840 3596
rect 511264 3544 511316 3596
rect 513564 3544 513616 3596
rect 518164 3544 518216 3596
rect 521844 3544 521896 3596
rect 525064 3544 525116 3596
rect 527732 3544 527784 3596
rect 479340 3476 479392 3528
rect 481640 3476 481692 3528
rect 482468 3476 482520 3528
rect 496084 3476 496136 3528
rect 497096 3476 497148 3528
rect 506480 3476 506532 3528
rect 507308 3476 507360 3528
rect 520924 3476 520976 3528
rect 523040 3476 523092 3528
rect 527824 3476 527876 3528
rect 533712 3544 533764 3596
rect 549904 3544 549956 3596
rect 551468 3544 551520 3596
rect 567844 3544 567896 3596
rect 571524 3544 571576 3596
rect 531320 3476 531372 3528
rect 532148 3476 532200 3528
rect 545764 3476 545816 3528
rect 546684 3476 546736 3528
rect 556160 3476 556212 3528
rect 556988 3476 557040 3528
rect 570604 3476 570656 3528
rect 572720 3476 572772 3528
rect 581000 3408 581052 3460
rect 493324 3340 493376 3392
rect 499396 3340 499448 3392
rect 543004 3340 543056 3392
rect 549076 3340 549128 3392
rect 428556 3272 428608 3324
rect 434444 3272 434496 3324
rect 509884 3272 509936 3324
rect 514760 3272 514812 3324
rect 342168 3204 342220 3256
rect 361764 3204 361816 3256
rect 446404 3204 446456 3256
rect 452108 3204 452160 3256
rect 216496 3136 216548 3188
rect 227536 3136 227588 3188
rect 345756 3136 345808 3188
rect 361856 3136 361908 3188
rect 485044 3136 485096 3188
rect 487620 3136 487672 3188
rect 534724 3136 534776 3188
rect 537208 3136 537260 3188
rect 560944 3136 560996 3188
rect 563244 3136 563296 3188
rect 19432 3000 19484 3052
rect 25596 3000 25648 3052
rect 195612 3000 195664 3052
rect 198096 3000 198148 3052
rect 374644 3000 374696 3052
rect 376484 3000 376536 3052
rect 413284 3000 413336 3052
rect 415492 3000 415544 3052
rect 417516 3000 417568 3052
rect 420184 3000 420236 3052
rect 464344 3000 464396 3052
rect 466276 3000 466328 3052
rect 486516 3000 486568 3052
rect 488816 3000 488868 3052
rect 514024 3000 514076 3052
rect 515956 3000 516008 3052
rect 522304 3000 522356 3052
rect 524236 3000 524288 3052
rect 538864 3000 538916 3052
rect 540796 3000 540848 3052
rect 563704 3000 563756 3052
rect 565636 3000 565688 3052
rect 571984 3000 572036 3052
rect 573916 3000 573968 3052
rect 378784 2932 378836 2984
rect 381176 2932 381228 2984
rect 396724 2932 396776 2984
rect 402520 2932 402572 2984
rect 457444 2932 457496 2984
rect 459192 2932 459244 2984
rect 552756 2932 552808 2984
rect 554964 2932 555016 2984
rect 13544 2864 13596 2916
rect 14464 2864 14516 2916
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 699718 8156 703520
rect 24320 700330 24348 703520
rect 24308 700324 24360 700330
rect 24308 700266 24360 700272
rect 8116 699712 8168 699718
rect 8116 699654 8168 699660
rect 10324 699712 10376 699718
rect 10324 699654 10376 699660
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 2780 632120 2832 632126
rect 2778 632088 2780 632097
rect 4804 632120 4856 632126
rect 2832 632088 2834 632097
rect 4804 632062 4856 632068
rect 2778 632023 2834 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3422 606112 3478 606121
rect 3422 606047 3424 606056
rect 3476 606047 3478 606056
rect 3424 606018 3476 606024
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 553722 3464 553823
rect 3424 553716 3476 553722
rect 3424 553658 3476 553664
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 527202 3464 527847
rect 3424 527196 3476 527202
rect 3424 527138 3476 527144
rect 3422 514856 3478 514865
rect 3422 514791 3424 514800
rect 3476 514791 3478 514800
rect 3424 514762 3476 514768
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3436 474774 3464 475623
rect 3424 474768 3476 474774
rect 3424 474710 3476 474716
rect 4816 467158 4844 632062
rect 7564 606076 7616 606082
rect 7564 606018 7616 606024
rect 7576 478174 7604 606018
rect 8944 553716 8996 553722
rect 8944 553658 8996 553664
rect 7564 478168 7616 478174
rect 7564 478110 7616 478116
rect 8956 474026 8984 553658
rect 8944 474020 8996 474026
rect 8944 473962 8996 473968
rect 4804 467152 4856 467158
rect 4804 467094 4856 467100
rect 3238 462632 3294 462641
rect 3238 462567 3294 462576
rect 3252 462398 3280 462567
rect 3240 462392 3292 462398
rect 3240 462334 3292 462340
rect 10336 460222 10364 699654
rect 21364 683188 21416 683194
rect 21364 683130 21416 683136
rect 13084 501016 13136 501022
rect 13084 500958 13136 500964
rect 13096 471306 13124 500958
rect 13084 471300 13136 471306
rect 13084 471242 13136 471248
rect 21376 465730 21404 683130
rect 28264 656940 28316 656946
rect 28264 656882 28316 656888
rect 21364 465724 21416 465730
rect 21364 465666 21416 465672
rect 10324 460216 10376 460222
rect 10324 460158 10376 460164
rect 28276 457502 28304 656882
rect 35164 527196 35216 527202
rect 35164 527138 35216 527144
rect 35176 469878 35204 527138
rect 35164 469872 35216 469878
rect 35164 469814 35216 469820
rect 28264 457496 28316 457502
rect 28264 457438 28316 457444
rect 40052 454714 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 57244 579692 57296 579698
rect 57244 579634 57296 579640
rect 57256 468518 57284 579634
rect 57244 468512 57296 468518
rect 57244 468454 57296 468460
rect 71792 461650 71820 702986
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 71780 461644 71832 461650
rect 71780 461586 71832 461592
rect 40040 454708 40092 454714
rect 40040 454650 40092 454656
rect 88352 450566 88380 702406
rect 105464 699786 105492 703520
rect 137848 700398 137876 703520
rect 154132 702434 154160 703520
rect 170324 702434 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 153212 702406 154160 702434
rect 169772 702406 170352 702434
rect 137836 700392 137888 700398
rect 137836 700334 137888 700340
rect 138664 700392 138716 700398
rect 138664 700334 138716 700340
rect 105452 699780 105504 699786
rect 105452 699722 105504 699728
rect 108304 699780 108356 699786
rect 108304 699722 108356 699728
rect 108316 451926 108344 699722
rect 138676 458930 138704 700334
rect 153212 472666 153240 702406
rect 153200 472660 153252 472666
rect 153200 472602 153252 472608
rect 138664 458924 138716 458930
rect 138664 458866 138716 458872
rect 169772 453422 169800 702406
rect 201512 456210 201540 702986
rect 217968 700392 218020 700398
rect 217968 700334 218020 700340
rect 215944 700324 215996 700330
rect 215944 700266 215996 700272
rect 217876 700324 217928 700330
rect 217876 700266 217928 700272
rect 214564 670744 214616 670750
rect 214564 670686 214616 670692
rect 211804 618316 211856 618322
rect 211804 618258 211856 618264
rect 210424 565888 210476 565894
rect 210424 565830 210476 565836
rect 207664 514820 207716 514826
rect 207664 514762 207716 514768
rect 201500 456204 201552 456210
rect 201500 456146 201552 456152
rect 169760 453416 169812 453422
rect 169760 453358 169812 453364
rect 207676 452062 207704 514762
rect 210436 461854 210464 565830
rect 210424 461848 210476 461854
rect 210424 461790 210476 461796
rect 211816 453558 211844 618258
rect 214576 459066 214604 670686
rect 214564 459060 214616 459066
rect 214564 459002 214616 459008
rect 215956 456278 215984 700266
rect 217784 565140 217836 565146
rect 217784 565082 217836 565088
rect 217598 516896 217654 516905
rect 217598 516831 217654 516840
rect 217506 513768 217562 513777
rect 217506 513703 217562 513712
rect 217414 489968 217470 489977
rect 217414 489903 217470 489912
rect 217322 488064 217378 488073
rect 217322 487999 217378 488008
rect 215944 456272 215996 456278
rect 215944 456214 215996 456220
rect 211804 453552 211856 453558
rect 211804 453494 211856 453500
rect 207664 452056 207716 452062
rect 207664 451998 207716 452004
rect 108304 451920 108356 451926
rect 108304 451862 108356 451868
rect 88340 450560 88392 450566
rect 88340 450502 88392 450508
rect 4066 449576 4122 449585
rect 4122 449534 4200 449562
rect 4066 449511 4122 449520
rect 4172 446554 4200 449534
rect 217336 447846 217364 487999
rect 217428 478378 217456 489903
rect 217416 478372 217468 478378
rect 217416 478314 217468 478320
rect 217520 474162 217548 513703
rect 217508 474156 217560 474162
rect 217508 474098 217560 474104
rect 217612 471374 217640 516831
rect 217690 515944 217746 515953
rect 217690 515879 217746 515888
rect 217600 471368 217652 471374
rect 217600 471310 217652 471316
rect 217704 467294 217732 515879
rect 217692 467288 217744 467294
rect 217692 467230 217744 467236
rect 217324 447840 217376 447846
rect 217324 447782 217376 447788
rect 4160 446548 4212 446554
rect 4160 446490 4212 446496
rect 206284 446072 206336 446078
rect 206284 446014 206336 446020
rect 203616 446004 203668 446010
rect 203616 445946 203668 445952
rect 192484 445936 192536 445942
rect 192484 445878 192536 445884
rect 8944 445800 8996 445806
rect 8944 445742 8996 445748
rect 7564 444508 7616 444514
rect 7564 444450 7616 444456
rect 3608 442468 3660 442474
rect 3608 442410 3660 442416
rect 3516 442400 3568 442406
rect 3516 442342 3568 442348
rect 3424 440904 3476 440910
rect 3424 440846 3476 440852
rect 3332 423632 3384 423638
rect 3330 423600 3332 423609
rect 3384 423600 3386 423609
rect 3330 423535 3386 423544
rect 2964 411256 3016 411262
rect 2964 411198 3016 411204
rect 2976 410553 3004 411198
rect 2962 410544 3018 410553
rect 2962 410479 3018 410488
rect 3056 398812 3108 398818
rect 3056 398754 3108 398760
rect 3068 397497 3096 398754
rect 3054 397488 3110 397497
rect 3054 397423 3110 397432
rect 3148 372564 3200 372570
rect 3148 372506 3200 372512
rect 3160 371385 3188 372506
rect 3146 371376 3202 371385
rect 3146 371311 3202 371320
rect 2964 320136 3016 320142
rect 2964 320078 3016 320084
rect 2976 319297 3004 320078
rect 2962 319288 3018 319297
rect 2962 319223 3018 319232
rect 3332 306332 3384 306338
rect 3332 306274 3384 306280
rect 3344 306241 3372 306274
rect 3330 306232 3386 306241
rect 3330 306167 3386 306176
rect 2780 284980 2832 284986
rect 2780 284922 2832 284928
rect 2792 16574 2820 284922
rect 2964 267708 3016 267714
rect 2964 267650 3016 267656
rect 2976 267209 3004 267650
rect 2962 267200 3018 267209
rect 2962 267135 3018 267144
rect 3332 254788 3384 254794
rect 3332 254730 3384 254736
rect 3344 254153 3372 254730
rect 3330 254144 3386 254153
rect 3330 254079 3386 254088
rect 3056 202836 3108 202842
rect 3056 202778 3108 202784
rect 3068 201929 3096 202778
rect 3054 201920 3110 201929
rect 3054 201855 3110 201864
rect 3436 110673 3464 440846
rect 3528 241097 3556 442342
rect 3620 293185 3648 442410
rect 3700 442264 3752 442270
rect 3700 442206 3752 442212
rect 3712 345409 3740 442206
rect 7576 423638 7604 444450
rect 7564 423632 7616 423638
rect 7564 423574 7616 423580
rect 3792 378820 3844 378826
rect 3792 378762 3844 378768
rect 3804 358465 3832 378762
rect 3790 358456 3846 358465
rect 3790 358391 3846 358400
rect 3698 345400 3754 345409
rect 3698 345335 3754 345344
rect 3606 293176 3662 293185
rect 3606 293111 3662 293120
rect 8300 290488 8352 290494
rect 8300 290430 8352 290436
rect 7564 262880 7616 262886
rect 7564 262822 7616 262828
rect 4160 247716 4212 247722
rect 4160 247658 4212 247664
rect 3514 241088 3570 241097
rect 3514 241023 3570 241032
rect 3516 189032 3568 189038
rect 3516 188974 3568 188980
rect 3528 188873 3556 188974
rect 3514 188864 3570 188873
rect 3514 188799 3570 188808
rect 3516 150408 3568 150414
rect 3516 150350 3568 150356
rect 3528 149841 3556 150350
rect 3514 149832 3570 149841
rect 3514 149767 3570 149776
rect 3516 137964 3568 137970
rect 3516 137906 3568 137912
rect 3528 136785 3556 137906
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 3424 97980 3476 97986
rect 3424 97922 3476 97928
rect 3436 97617 3464 97922
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 4172 16574 4200 247658
rect 6920 246356 6972 246362
rect 6920 246298 6972 246304
rect 6932 16574 6960 246298
rect 2792 16546 2912 16574
rect 4172 16546 5304 16574
rect 6932 16546 7512 16574
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 1688 480 1716 3538
rect 2884 480 2912 16546
rect 4068 3868 4120 3874
rect 4068 3810 4120 3816
rect 4080 480 4108 3810
rect 5276 480 5304 16546
rect 6460 3664 6512 3670
rect 6460 3606 6512 3612
rect 6472 480 6500 3606
rect 7484 3482 7512 16546
rect 7576 3874 7604 262822
rect 8312 16574 8340 290430
rect 8956 254794 8984 445742
rect 100024 444644 100076 444650
rect 100024 444586 100076 444592
rect 98644 444576 98696 444582
rect 98644 444518 98696 444524
rect 94504 443828 94556 443834
rect 94504 443770 94556 443776
rect 64144 441856 64196 441862
rect 64144 441798 64196 441804
rect 25504 440360 25556 440366
rect 25504 440302 25556 440308
rect 20718 300112 20774 300121
rect 20718 300047 20774 300056
rect 13084 293276 13136 293282
rect 13084 293218 13136 293224
rect 9680 289128 9732 289134
rect 9680 289070 9732 289076
rect 8944 254788 8996 254794
rect 8944 254730 8996 254736
rect 8312 16546 8800 16574
rect 7564 3868 7616 3874
rect 7564 3810 7616 3816
rect 7484 3454 7696 3482
rect 7668 480 7696 3454
rect 8772 480 8800 16546
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 289070
rect 11060 265668 11112 265674
rect 11060 265610 11112 265616
rect 11072 16574 11100 265610
rect 11072 16546 11192 16574
rect 11164 480 11192 16546
rect 13096 3534 13124 293218
rect 18604 286340 18656 286346
rect 18604 286282 18656 286288
rect 16580 283620 16632 283626
rect 16580 283562 16632 283568
rect 14464 273964 14516 273970
rect 14464 273906 14516 273912
rect 13820 261520 13872 261526
rect 13820 261462 13872 261468
rect 13832 16574 13860 261462
rect 13832 16546 14320 16574
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 12360 480 12388 3470
rect 13544 2916 13596 2922
rect 13544 2858 13596 2864
rect 13556 480 13584 2858
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 14476 2922 14504 273906
rect 16592 16574 16620 283562
rect 17960 256012 18012 256018
rect 17960 255954 18012 255960
rect 16592 16546 17080 16574
rect 15936 3528 15988 3534
rect 15936 3470 15988 3476
rect 14464 2916 14516 2922
rect 14464 2858 14516 2864
rect 15948 480 15976 3470
rect 17052 480 17080 16546
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 255954
rect 18616 3670 18644 286282
rect 19340 260160 19392 260166
rect 19340 260102 19392 260108
rect 19352 16574 19380 260102
rect 20732 16574 20760 300047
rect 22100 287700 22152 287706
rect 22100 287642 22152 287648
rect 22112 16574 22140 287642
rect 23480 257372 23532 257378
rect 23480 257314 23532 257320
rect 23492 16574 23520 257314
rect 25516 59362 25544 440302
rect 32404 373176 32456 373182
rect 32404 373118 32456 373124
rect 27620 291848 27672 291854
rect 27620 291790 27672 291796
rect 26240 285048 26292 285054
rect 26240 284990 26292 284996
rect 25596 257440 25648 257446
rect 25596 257382 25648 257388
rect 25504 59356 25556 59362
rect 25504 59298 25556 59304
rect 19352 16546 20208 16574
rect 20732 16546 21864 16574
rect 22112 16546 22600 16574
rect 23492 16546 24256 16574
rect 18604 3664 18656 3670
rect 18604 3606 18656 3612
rect 19432 3052 19484 3058
rect 19432 2994 19484 3000
rect 19444 480 19472 2994
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20180 354 20208 16546
rect 21836 480 21864 16546
rect 20598 354 20710 480
rect 20180 326 20710 354
rect 20598 -960 20710 326
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 24228 480 24256 16546
rect 25320 3664 25372 3670
rect 25320 3606 25372 3612
rect 25332 480 25360 3606
rect 25608 3058 25636 257382
rect 25596 3052 25648 3058
rect 25596 2994 25648 3000
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 284990
rect 27632 6914 27660 291790
rect 27712 276684 27764 276690
rect 27712 276626 27764 276632
rect 27724 16574 27752 276626
rect 30380 260228 30432 260234
rect 30380 260170 30432 260176
rect 30392 16574 30420 260170
rect 31760 244928 31812 244934
rect 31760 244870 31812 244876
rect 31772 16574 31800 244870
rect 27724 16546 28488 16574
rect 30392 16546 30880 16574
rect 31772 16546 31984 16574
rect 27632 6886 27752 6914
rect 27724 480 27752 6886
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28460 354 28488 16546
rect 30104 3732 30156 3738
rect 30104 3674 30156 3680
rect 30116 480 30144 3674
rect 28878 354 28990 480
rect 28460 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 32416 3602 32444 373118
rect 43444 294636 43496 294642
rect 43444 294578 43496 294584
rect 40040 286408 40092 286414
rect 40040 286350 40092 286356
rect 34520 280832 34572 280838
rect 34520 280774 34572 280780
rect 32404 3596 32456 3602
rect 32404 3538 32456 3544
rect 33600 3596 33652 3602
rect 33600 3538 33652 3544
rect 33612 480 33640 3538
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 280774
rect 38660 279472 38712 279478
rect 38660 279414 38712 279420
rect 35900 278044 35952 278050
rect 35900 277986 35952 277992
rect 35164 247784 35216 247790
rect 35164 247726 35216 247732
rect 35176 3602 35204 247726
rect 35912 16574 35940 277986
rect 38672 16574 38700 279414
rect 39304 265736 39356 265742
rect 39304 265678 39356 265684
rect 35912 16546 36032 16574
rect 38672 16546 39160 16574
rect 35164 3596 35216 3602
rect 35164 3538 35216 3544
rect 36004 480 36032 16546
rect 38384 3596 38436 3602
rect 38384 3538 38436 3544
rect 37188 3392 37240 3398
rect 37188 3334 37240 3340
rect 37200 480 37228 3334
rect 38396 480 38424 3538
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 39316 3602 39344 265678
rect 39396 260296 39448 260302
rect 39396 260238 39448 260244
rect 39408 3738 39436 260238
rect 40052 16574 40080 286350
rect 42800 275324 42852 275330
rect 42800 275266 42852 275272
rect 41420 247852 41472 247858
rect 41420 247794 41472 247800
rect 41432 16574 41460 247794
rect 40052 16546 40264 16574
rect 41432 16546 41920 16574
rect 39396 3732 39448 3738
rect 39396 3674 39448 3680
rect 39304 3596 39356 3602
rect 39304 3538 39356 3544
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 41892 480 41920 16546
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 275266
rect 43456 3398 43484 294578
rect 58624 293344 58676 293350
rect 58624 293286 58676 293292
rect 57244 290556 57296 290562
rect 57244 290498 57296 290504
rect 46940 286476 46992 286482
rect 46940 286418 46992 286424
rect 44180 282192 44232 282198
rect 44180 282134 44232 282140
rect 44192 16574 44220 282134
rect 46204 251864 46256 251870
rect 46204 251806 46256 251812
rect 44192 16546 45048 16574
rect 44272 3732 44324 3738
rect 44272 3674 44324 3680
rect 43444 3392 43496 3398
rect 43444 3334 43496 3340
rect 44284 480 44312 3674
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45020 354 45048 16546
rect 46216 3738 46244 251806
rect 46952 16574 46980 286418
rect 53840 272536 53892 272542
rect 53840 272478 53892 272484
rect 52460 262948 52512 262954
rect 52460 262890 52512 262896
rect 49700 251932 49752 251938
rect 49700 251874 49752 251880
rect 48320 246424 48372 246430
rect 48320 246366 48372 246372
rect 48332 16574 48360 246366
rect 49712 16574 49740 251874
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 49712 16546 50200 16574
rect 46204 3732 46256 3738
rect 46204 3674 46256 3680
rect 46664 3732 46716 3738
rect 46664 3674 46716 3680
rect 46676 480 46704 3674
rect 45438 354 45550 480
rect 45020 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50172 480 50200 16546
rect 51356 4072 51408 4078
rect 51356 4014 51408 4020
rect 51368 480 51396 4014
rect 52472 3602 52500 262890
rect 52552 250504 52604 250510
rect 52552 250446 52604 250452
rect 52460 3596 52512 3602
rect 52460 3538 52512 3544
rect 52564 480 52592 250446
rect 53852 16574 53880 272478
rect 53852 16546 54984 16574
rect 53380 3596 53432 3602
rect 53380 3538 53432 3544
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53392 354 53420 3538
rect 54956 480 54984 16546
rect 57256 4078 57284 290498
rect 57980 271176 58032 271182
rect 57980 271118 58032 271124
rect 57336 249076 57388 249082
rect 57336 249018 57388 249024
rect 57244 4072 57296 4078
rect 57244 4014 57296 4020
rect 57348 3602 57376 249018
rect 57992 16574 58020 271118
rect 57992 16546 58480 16574
rect 56048 3596 56100 3602
rect 56048 3538 56100 3544
rect 57336 3596 57388 3602
rect 57336 3538 57388 3544
rect 56060 480 56088 3538
rect 57244 3392 57296 3398
rect 57244 3334 57296 3340
rect 57256 480 57284 3334
rect 58452 480 58480 16546
rect 58636 3398 58664 293286
rect 63500 260364 63552 260370
rect 63500 260306 63552 260312
rect 60740 250708 60792 250714
rect 60740 250650 60792 250656
rect 60752 6914 60780 250650
rect 62120 249144 62172 249150
rect 62120 249086 62172 249092
rect 60832 244996 60884 245002
rect 60832 244938 60884 244944
rect 60844 16574 60872 244938
rect 62132 16574 62160 249086
rect 63512 16574 63540 260306
rect 64156 20670 64184 441798
rect 94516 306338 94544 443770
rect 95882 440328 95938 440337
rect 95882 440263 95938 440272
rect 94504 306332 94556 306338
rect 94504 306274 94556 306280
rect 71044 291916 71096 291922
rect 71044 291858 71096 291864
rect 70400 267028 70452 267034
rect 70400 266970 70452 266976
rect 69020 264240 69072 264246
rect 69020 264182 69072 264188
rect 67640 250640 67692 250646
rect 67640 250582 67692 250588
rect 66260 250572 66312 250578
rect 66260 250514 66312 250520
rect 64880 246492 64932 246498
rect 64880 246434 64932 246440
rect 64144 20664 64196 20670
rect 64144 20606 64196 20612
rect 64892 16574 64920 246434
rect 66272 16574 66300 250514
rect 60844 16546 61608 16574
rect 62132 16546 63264 16574
rect 63512 16546 64368 16574
rect 64892 16546 65104 16574
rect 66272 16546 66760 16574
rect 60752 6886 60872 6914
rect 59636 3596 59688 3602
rect 59636 3538 59688 3544
rect 58624 3392 58676 3398
rect 58624 3334 58676 3340
rect 59648 480 59676 3538
rect 60844 480 60872 6886
rect 53718 354 53830 480
rect 53392 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61580 354 61608 16546
rect 63236 480 63264 16546
rect 64340 480 64368 16546
rect 61998 354 62110 480
rect 61580 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66732 480 66760 16546
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 250582
rect 69032 16574 69060 264182
rect 70412 16574 70440 266970
rect 69032 16546 69888 16574
rect 70412 16546 70992 16574
rect 69112 3800 69164 3806
rect 69112 3742 69164 3748
rect 69124 480 69152 3742
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 16546
rect 70964 3482 70992 16546
rect 71056 3806 71084 291858
rect 81440 285116 81492 285122
rect 81440 285058 81492 285064
rect 71780 279540 71832 279546
rect 71780 279482 71832 279488
rect 71792 16574 71820 279482
rect 78680 278112 78732 278118
rect 78680 278054 78732 278060
rect 75920 269816 75972 269822
rect 75920 269758 75972 269764
rect 73160 261588 73212 261594
rect 73160 261530 73212 261536
rect 73172 16574 73200 261530
rect 74540 249212 74592 249218
rect 74540 249154 74592 249160
rect 74552 16574 74580 249154
rect 71792 16546 72648 16574
rect 73172 16546 73384 16574
rect 74552 16546 75040 16574
rect 71044 3800 71096 3806
rect 71044 3742 71096 3748
rect 70964 3454 71544 3482
rect 71516 480 71544 3454
rect 72620 480 72648 16546
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 16546
rect 75012 480 75040 16546
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 269758
rect 77300 268388 77352 268394
rect 77300 268330 77352 268336
rect 77312 6914 77340 268330
rect 77392 256080 77444 256086
rect 77392 256022 77444 256028
rect 77404 16574 77432 256022
rect 78692 16574 78720 278054
rect 80060 253224 80112 253230
rect 80060 253166 80112 253172
rect 80072 16574 80100 253166
rect 81452 16574 81480 285058
rect 93860 274032 93912 274038
rect 93860 273974 93912 273980
rect 84200 272604 84252 272610
rect 84200 272546 84252 272552
rect 82820 249280 82872 249286
rect 82820 249222 82872 249228
rect 82832 16574 82860 249222
rect 77404 16546 78168 16574
rect 78692 16546 79272 16574
rect 80072 16546 80928 16574
rect 81452 16546 81664 16574
rect 82832 16546 83320 16574
rect 77312 6886 77432 6914
rect 77404 480 77432 6886
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78140 354 78168 16546
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 79244 354 79272 16546
rect 80900 480 80928 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83292 480 83320 16546
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 272546
rect 92480 256148 92532 256154
rect 92480 256090 92532 256096
rect 91100 254720 91152 254726
rect 91100 254662 91152 254668
rect 88340 254652 88392 254658
rect 88340 254594 88392 254600
rect 86960 254584 87012 254590
rect 86960 254526 87012 254532
rect 85580 253292 85632 253298
rect 85580 253234 85632 253240
rect 85592 6914 85620 253234
rect 85672 246560 85724 246566
rect 85672 246502 85724 246508
rect 85684 16574 85712 246502
rect 86972 16574 87000 254526
rect 88352 16574 88380 254594
rect 89720 247920 89772 247926
rect 89720 247862 89772 247868
rect 89732 16574 89760 247862
rect 91112 16574 91140 254662
rect 85684 16546 86448 16574
rect 86972 16546 87552 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 85592 6886 85712 6914
rect 85684 480 85712 6886
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86420 354 86448 16546
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 87524 354 87552 16546
rect 89180 480 89208 16546
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 256090
rect 93872 6914 93900 273974
rect 93952 269884 94004 269890
rect 93952 269826 94004 269832
rect 93964 16574 93992 269826
rect 95240 254788 95292 254794
rect 95240 254730 95292 254736
rect 95252 16574 95280 254730
rect 95896 33114 95924 440263
rect 97816 377460 97868 377466
rect 97816 377402 97868 377408
rect 97724 371612 97776 371618
rect 97724 371554 97776 371560
rect 97632 371544 97684 371550
rect 97632 371486 97684 371492
rect 97644 362001 97672 371486
rect 97736 364721 97764 371554
rect 97722 364712 97778 364721
rect 97722 364647 97778 364656
rect 97630 361992 97686 362001
rect 97630 361927 97686 361936
rect 97828 351121 97856 377402
rect 97908 371408 97960 371414
rect 97908 371350 97960 371356
rect 97920 367441 97948 371350
rect 97906 367432 97962 367441
rect 97906 367367 97962 367376
rect 97906 356552 97962 356561
rect 97906 356487 97962 356496
rect 97814 351112 97870 351121
rect 97814 351047 97870 351056
rect 97814 348392 97870 348401
rect 97814 348327 97870 348336
rect 97722 345672 97778 345681
rect 97722 345607 97778 345616
rect 97630 340232 97686 340241
rect 97630 340167 97686 340176
rect 97538 334792 97594 334801
rect 97538 334727 97594 334736
rect 97446 332072 97502 332081
rect 97446 332007 97502 332016
rect 97354 326632 97410 326641
rect 97354 326567 97410 326576
rect 97264 305108 97316 305114
rect 97264 305050 97316 305056
rect 97276 299169 97304 305050
rect 97368 300830 97396 326567
rect 97356 300824 97408 300830
rect 97356 300766 97408 300772
rect 97460 299441 97488 332007
rect 97552 305114 97580 334727
rect 97540 305108 97592 305114
rect 97540 305050 97592 305056
rect 97540 304972 97592 304978
rect 97540 304914 97592 304920
rect 97446 299432 97502 299441
rect 97446 299367 97502 299376
rect 97552 299305 97580 304914
rect 97644 300490 97672 340167
rect 97736 300694 97764 345607
rect 97724 300688 97776 300694
rect 97724 300630 97776 300636
rect 97828 300626 97856 348327
rect 97920 304978 97948 356487
rect 98656 320142 98684 444518
rect 100036 372570 100064 444586
rect 140780 443148 140832 443154
rect 140780 443090 140832 443096
rect 140792 383654 140820 443090
rect 140792 383626 141464 383654
rect 110972 374808 111024 374814
rect 110972 374750 111024 374756
rect 100668 374740 100720 374746
rect 100668 374682 100720 374688
rect 100024 372564 100076 372570
rect 100024 372506 100076 372512
rect 100680 372028 100708 374682
rect 105820 374468 105872 374474
rect 105820 374410 105872 374416
rect 103244 372972 103296 372978
rect 103244 372914 103296 372920
rect 103256 372028 103284 372914
rect 105832 372028 105860 374410
rect 108396 374332 108448 374338
rect 108396 374274 108448 374280
rect 108408 372028 108436 374274
rect 110984 372028 111012 374750
rect 126428 374672 126480 374678
rect 126428 374614 126480 374620
rect 121276 374604 121328 374610
rect 121276 374546 121328 374552
rect 118700 373040 118752 373046
rect 118700 372982 118752 372988
rect 113548 372700 113600 372706
rect 113548 372642 113600 372648
rect 113560 372028 113588 372642
rect 118712 372028 118740 372982
rect 121288 372028 121316 374546
rect 123852 373108 123904 373114
rect 123852 373050 123904 373056
rect 123864 372028 123892 373050
rect 126440 372028 126468 374614
rect 139308 374060 139360 374066
rect 139308 374002 139360 374008
rect 134156 372904 134208 372910
rect 134156 372846 134208 372852
rect 131580 372836 131632 372842
rect 131580 372778 131632 372784
rect 129004 372768 129056 372774
rect 129004 372710 129056 372716
rect 129016 372028 129044 372710
rect 131592 372028 131620 372778
rect 134168 372028 134196 372846
rect 139320 372028 139348 374002
rect 141436 372042 141464 383626
rect 154764 374876 154816 374882
rect 154764 374818 154816 374824
rect 173164 374876 173216 374882
rect 173164 374818 173216 374824
rect 152188 374264 152240 374270
rect 152188 374206 152240 374212
rect 147036 374196 147088 374202
rect 147036 374138 147088 374144
rect 141436 372014 141910 372042
rect 147048 372028 147076 374138
rect 149612 372632 149664 372638
rect 149612 372574 149664 372580
rect 149624 372028 149652 372574
rect 152200 372028 152228 374206
rect 154776 372028 154804 374818
rect 170588 374672 170640 374678
rect 170588 374614 170640 374620
rect 165528 374536 165580 374542
rect 165528 374478 165580 374484
rect 157340 374400 157392 374406
rect 157340 374342 157392 374348
rect 155868 374060 155920 374066
rect 155868 374002 155920 374008
rect 155880 373289 155908 374002
rect 155866 373280 155922 373289
rect 155866 373215 155922 373224
rect 157352 372028 157380 374342
rect 159914 374096 159970 374105
rect 159914 374031 159970 374040
rect 162492 374060 162544 374066
rect 159928 372028 159956 374031
rect 162492 374002 162544 374008
rect 162504 372028 162532 374002
rect 165540 373182 165568 374478
rect 170404 374060 170456 374066
rect 170404 374002 170456 374008
rect 165068 373176 165120 373182
rect 165068 373118 165120 373124
rect 165528 373176 165580 373182
rect 165528 373118 165580 373124
rect 165080 372028 165108 373118
rect 136758 371890 137048 371906
rect 124772 371884 124824 371890
rect 124772 371826 124824 371832
rect 128268 371884 128320 371890
rect 136758 371884 137060 371890
rect 136758 371878 137008 371884
rect 128268 371826 128320 371832
rect 137008 371826 137060 371832
rect 138480 371884 138532 371890
rect 138480 371826 138532 371832
rect 116400 371680 116452 371686
rect 116150 371628 116400 371634
rect 116150 371622 116452 371628
rect 124678 371648 124734 371657
rect 116150 371606 116440 371622
rect 124784 371618 124812 371826
rect 125692 371816 125744 371822
rect 125692 371758 125744 371764
rect 125704 371618 125732 371758
rect 128280 371754 128308 371826
rect 138020 371816 138072 371822
rect 138020 371758 138072 371764
rect 128268 371748 128320 371754
rect 128268 371690 128320 371696
rect 135074 371648 135130 371657
rect 124678 371583 124680 371592
rect 124732 371583 124734 371592
rect 124772 371612 124824 371618
rect 124680 371554 124732 371560
rect 124772 371554 124824 371560
rect 125692 371612 125744 371618
rect 137926 371648 137982 371657
rect 135130 371618 135254 371634
rect 135130 371612 135266 371618
rect 135130 371606 135214 371612
rect 135074 371583 135130 371592
rect 125692 371554 125744 371560
rect 138032 371618 138060 371758
rect 138492 371618 138520 371826
rect 144000 371816 144052 371822
rect 144000 371758 144052 371764
rect 144012 371618 144040 371758
rect 167670 371754 167960 371770
rect 167670 371748 167972 371754
rect 167670 371742 167920 371748
rect 167920 371690 167972 371696
rect 144736 371680 144788 371686
rect 144182 371648 144238 371657
rect 137926 371583 137928 371592
rect 135214 371554 135266 371560
rect 137980 371583 137982 371592
rect 138020 371612 138072 371618
rect 137928 371554 137980 371560
rect 138020 371554 138072 371560
rect 138480 371612 138532 371618
rect 138480 371554 138532 371560
rect 144000 371612 144052 371618
rect 144486 371628 144736 371634
rect 144486 371622 144788 371628
rect 144486 371606 144776 371622
rect 144182 371583 144184 371592
rect 144000 371554 144052 371560
rect 144236 371583 144238 371592
rect 144184 371554 144236 371560
rect 99840 371476 99892 371482
rect 169602 371470 169984 371498
rect 99840 371418 99892 371424
rect 99852 370705 99880 371418
rect 99838 370696 99894 370705
rect 99838 370631 99894 370640
rect 169956 367946 169984 371470
rect 169944 367940 169996 367946
rect 169944 367882 169996 367888
rect 99286 359272 99342 359281
rect 99286 359207 99342 359216
rect 99194 353832 99250 353841
rect 99194 353767 99250 353776
rect 99102 337512 99158 337521
rect 99102 337447 99158 337456
rect 99010 329352 99066 329361
rect 99010 329287 99066 329296
rect 98918 323912 98974 323921
rect 98918 323847 98974 323856
rect 98644 320136 98696 320142
rect 98644 320078 98696 320084
rect 98826 318472 98882 318481
rect 98826 318407 98882 318416
rect 98734 315752 98790 315761
rect 98734 315687 98790 315696
rect 98642 310312 98698 310321
rect 98642 310247 98698 310256
rect 97908 304972 97960 304978
rect 97908 304914 97960 304920
rect 97906 304872 97962 304881
rect 97906 304807 97962 304816
rect 97816 300620 97868 300626
rect 97816 300562 97868 300568
rect 97632 300484 97684 300490
rect 97632 300426 97684 300432
rect 97920 299402 97948 304807
rect 98656 300762 98684 310247
rect 98644 300756 98696 300762
rect 98644 300698 98696 300704
rect 97908 299396 97960 299402
rect 97908 299338 97960 299344
rect 97538 299296 97594 299305
rect 97538 299231 97594 299240
rect 97262 299160 97318 299169
rect 97262 299095 97318 299104
rect 98748 296682 98776 315687
rect 98840 299470 98868 318407
rect 98828 299464 98880 299470
rect 98828 299406 98880 299412
rect 98932 299266 98960 323847
rect 99024 300014 99052 329287
rect 99116 300558 99144 337447
rect 99104 300552 99156 300558
rect 99104 300494 99156 300500
rect 99208 300218 99236 353767
rect 99300 300801 99328 359207
rect 99378 342952 99434 342961
rect 99378 342887 99434 342896
rect 99286 300792 99342 300801
rect 99286 300727 99342 300736
rect 99392 300422 99420 342887
rect 99470 321192 99526 321201
rect 99470 321127 99526 321136
rect 99380 300416 99432 300422
rect 99380 300358 99432 300364
rect 99196 300212 99248 300218
rect 99196 300154 99248 300160
rect 99484 300150 99512 321127
rect 99562 313032 99618 313041
rect 99562 312967 99618 312976
rect 99576 300354 99604 312967
rect 99838 307592 99894 307601
rect 99838 307527 99894 307536
rect 99746 301608 99802 301617
rect 99746 301543 99802 301552
rect 99564 300348 99616 300354
rect 99564 300290 99616 300296
rect 99472 300144 99524 300150
rect 99472 300086 99524 300092
rect 99012 300008 99064 300014
rect 99012 299950 99064 299956
rect 99760 299334 99788 301543
rect 99852 300286 99880 307527
rect 170416 307222 170444 374002
rect 170496 372632 170548 372638
rect 170496 372574 170548 372580
rect 170508 308650 170536 372574
rect 170600 309369 170628 374614
rect 170956 374604 171008 374610
rect 170956 374546 171008 374552
rect 170772 371748 170824 371754
rect 170772 371690 170824 371696
rect 170680 367940 170732 367946
rect 170680 367882 170732 367888
rect 170586 309360 170642 309369
rect 170586 309295 170642 309304
rect 170692 309262 170720 367882
rect 170680 309256 170732 309262
rect 170784 309233 170812 371690
rect 170968 309505 170996 374546
rect 171784 374468 171836 374474
rect 171784 374410 171836 374416
rect 171690 358592 171746 358601
rect 171690 358527 171746 358536
rect 171704 357474 171732 358527
rect 171692 357468 171744 357474
rect 171692 357410 171744 357416
rect 171138 350432 171194 350441
rect 171138 350367 171194 350376
rect 171152 345098 171180 350367
rect 171140 345092 171192 345098
rect 171140 345034 171192 345040
rect 170954 309496 171010 309505
rect 170954 309431 171010 309440
rect 170680 309198 170732 309204
rect 170770 309224 170826 309233
rect 170770 309159 170826 309168
rect 170496 308644 170548 308650
rect 170496 308586 170548 308592
rect 170404 307216 170456 307222
rect 170404 307158 170456 307164
rect 170588 307148 170640 307154
rect 170588 307090 170640 307096
rect 169852 306332 169904 306338
rect 169852 306274 169904 306280
rect 169760 303000 169812 303006
rect 169760 302942 169812 302948
rect 169772 300642 169800 302942
rect 168958 300614 169800 300642
rect 164238 300384 164294 300393
rect 164238 300319 164294 300328
rect 99840 300280 99892 300286
rect 99840 300222 99892 300228
rect 160098 300248 160154 300257
rect 160098 300183 160154 300192
rect 99748 299328 99800 299334
rect 99748 299270 99800 299276
rect 98920 299260 98972 299266
rect 98920 299202 98972 299208
rect 100036 297770 100064 300084
rect 101968 298081 101996 300084
rect 103532 300070 104558 300098
rect 101954 298072 102010 298081
rect 101954 298007 102010 298016
rect 100024 297764 100076 297770
rect 100024 297706 100076 297712
rect 98736 296676 98788 296682
rect 98736 296618 98788 296624
rect 103532 296614 103560 300070
rect 107120 298110 107148 300084
rect 107108 298104 107160 298110
rect 107108 298046 107160 298052
rect 109696 297702 109724 300084
rect 111156 298104 111208 298110
rect 111156 298046 111208 298052
rect 109684 297696 109736 297702
rect 109684 297638 109736 297644
rect 103520 296608 103572 296614
rect 103520 296550 103572 296556
rect 111168 296546 111196 298046
rect 112272 297158 112300 300084
rect 114848 299198 114876 300084
rect 114836 299192 114888 299198
rect 114836 299134 114888 299140
rect 117424 298042 117452 300084
rect 120000 299130 120028 300084
rect 119988 299124 120040 299130
rect 119988 299066 120040 299072
rect 117412 298036 117464 298042
rect 117412 297978 117464 297984
rect 122576 297974 122604 300084
rect 125152 298994 125180 300084
rect 125140 298988 125192 298994
rect 125140 298930 125192 298936
rect 122564 297968 122616 297974
rect 122564 297910 122616 297916
rect 127728 297838 127756 300084
rect 130304 299062 130332 300084
rect 130292 299056 130344 299062
rect 130292 298998 130344 299004
rect 127716 297832 127768 297838
rect 127716 297774 127768 297780
rect 112260 297152 112312 297158
rect 112260 297094 112312 297100
rect 132880 297090 132908 300084
rect 133788 298784 133840 298790
rect 133788 298726 133840 298732
rect 133800 298042 133828 298726
rect 133788 298036 133840 298042
rect 133788 297978 133840 297984
rect 135456 297634 135484 300084
rect 138032 297906 138060 300084
rect 140608 298926 140636 300084
rect 140596 298920 140648 298926
rect 140596 298862 140648 298868
rect 138020 297900 138072 297906
rect 138020 297842 138072 297848
rect 135444 297628 135496 297634
rect 135444 297570 135496 297576
rect 143184 297566 143212 300084
rect 143448 298852 143500 298858
rect 143448 298794 143500 298800
rect 143460 297838 143488 298794
rect 145760 297945 145788 300084
rect 145746 297936 145802 297945
rect 145746 297871 145802 297880
rect 148336 297838 148364 300084
rect 143448 297832 143500 297838
rect 143448 297774 143500 297780
rect 148324 297832 148376 297838
rect 148324 297774 148376 297780
rect 143172 297560 143224 297566
rect 143172 297502 143224 297508
rect 150912 297498 150940 300084
rect 153212 300070 153502 300098
rect 150900 297492 150952 297498
rect 150900 297434 150952 297440
rect 132868 297084 132920 297090
rect 132868 297026 132920 297032
rect 111156 296540 111208 296546
rect 111156 296482 111208 296488
rect 153212 296478 153240 300070
rect 156064 298722 156092 300084
rect 156052 298716 156104 298722
rect 156052 298658 156104 298664
rect 158640 298042 158668 300084
rect 158628 298036 158680 298042
rect 158628 297978 158680 297984
rect 153200 296472 153252 296478
rect 153200 296414 153252 296420
rect 129740 296064 129792 296070
rect 129740 296006 129792 296012
rect 125600 295996 125652 296002
rect 125600 295938 125652 295944
rect 103520 289196 103572 289202
rect 103520 289138 103572 289144
rect 98000 279608 98052 279614
rect 98000 279550 98052 279556
rect 96620 275392 96672 275398
rect 96620 275334 96672 275340
rect 95884 33108 95936 33114
rect 95884 33050 95936 33056
rect 96632 16574 96660 275334
rect 98012 16574 98040 279550
rect 102140 278180 102192 278186
rect 102140 278122 102192 278128
rect 99380 272672 99432 272678
rect 99380 272614 99432 272620
rect 99392 16574 99420 272614
rect 100760 245064 100812 245070
rect 100760 245006 100812 245012
rect 93964 16546 94728 16574
rect 95252 16546 95832 16574
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 93872 6886 93992 6914
rect 93964 480 93992 6886
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94700 354 94728 16546
rect 95118 354 95230 480
rect 94700 326 95230 354
rect 95804 354 95832 16546
rect 97460 480 97488 16546
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 245006
rect 102152 6914 102180 278122
rect 102232 271244 102284 271250
rect 102232 271186 102284 271192
rect 102244 16574 102272 271186
rect 103532 16574 103560 289138
rect 114560 282260 114612 282266
rect 114560 282202 114612 282208
rect 107660 280900 107712 280906
rect 107660 280842 107712 280848
rect 106280 257508 106332 257514
rect 106280 257450 106332 257456
rect 104900 246628 104952 246634
rect 104900 246570 104952 246576
rect 104912 16574 104940 246570
rect 106292 16574 106320 257450
rect 107672 16574 107700 280842
rect 111800 276752 111852 276758
rect 111800 276694 111852 276700
rect 110420 269952 110472 269958
rect 110420 269894 110472 269900
rect 109040 245132 109092 245138
rect 109040 245074 109092 245080
rect 102244 16546 103376 16574
rect 103532 16546 104112 16574
rect 104912 16546 105768 16574
rect 106292 16546 106504 16574
rect 107672 16546 108160 16574
rect 102152 6886 102272 6914
rect 102244 480 102272 6886
rect 103348 480 103376 16546
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105740 480 105768 16546
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108132 480 108160 16546
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109052 354 109080 245074
rect 110432 6914 110460 269894
rect 110512 253360 110564 253366
rect 110512 253302 110564 253308
rect 110524 16574 110552 253302
rect 111812 16574 111840 276694
rect 113180 274100 113232 274106
rect 113180 274042 113232 274048
rect 113192 16574 113220 274042
rect 114572 16574 114600 282202
rect 115940 275460 115992 275466
rect 115940 275402 115992 275408
rect 115952 16574 115980 275402
rect 121460 265804 121512 265810
rect 121460 265746 121512 265752
rect 117320 257576 117372 257582
rect 117320 257518 117372 257524
rect 110524 16546 111656 16574
rect 111812 16546 112392 16574
rect 113192 16546 114048 16574
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 110432 6886 110552 6914
rect 110524 480 110552 6886
rect 111628 480 111656 16546
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114020 480 114048 16546
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 257518
rect 118700 256216 118752 256222
rect 118700 256158 118752 256164
rect 118712 3398 118740 256158
rect 118792 253428 118844 253434
rect 118792 253370 118844 253376
rect 118700 3392 118752 3398
rect 118700 3334 118752 3340
rect 118804 480 118832 253370
rect 120080 246696 120132 246702
rect 120080 246638 120132 246644
rect 120092 16574 120120 246638
rect 121472 16574 121500 265746
rect 124220 260432 124272 260438
rect 124220 260374 124272 260380
rect 122840 256284 122892 256290
rect 122840 256226 122892 256232
rect 122852 16574 122880 256226
rect 124232 16574 124260 260374
rect 120092 16546 120672 16574
rect 121472 16546 122328 16574
rect 122852 16546 123064 16574
rect 124232 16546 124720 16574
rect 119896 3392 119948 3398
rect 119896 3334 119948 3340
rect 119908 480 119936 3334
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 122300 480 122328 16546
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124692 480 124720 16546
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125612 354 125640 295938
rect 128360 291984 128412 291990
rect 128360 291926 128412 291932
rect 126980 280968 127032 280974
rect 126980 280910 127032 280916
rect 126992 480 127020 280910
rect 127072 275528 127124 275534
rect 127072 275470 127124 275476
rect 127084 16574 127112 275470
rect 128372 16574 128400 291926
rect 129752 16574 129780 296006
rect 135260 294704 135312 294710
rect 135260 294646 135312 294652
rect 132500 289264 132552 289270
rect 132500 289206 132552 289212
rect 131120 282328 131172 282334
rect 131120 282270 131172 282276
rect 131132 16574 131160 282270
rect 132512 16574 132540 289206
rect 133880 265872 133932 265878
rect 133880 265814 133932 265820
rect 127084 16546 128216 16574
rect 128372 16546 128952 16574
rect 129752 16546 130608 16574
rect 131132 16546 131344 16574
rect 132512 16546 133000 16574
rect 128188 480 128216 16546
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 16546
rect 130580 480 130608 16546
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 132972 480 133000 16546
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 133892 354 133920 265814
rect 135272 3806 135300 294646
rect 143540 290624 143592 290630
rect 143540 290566 143592 290572
rect 139400 287768 139452 287774
rect 139400 287710 139452 287716
rect 138020 283688 138072 283694
rect 138020 283630 138072 283636
rect 136640 276820 136692 276826
rect 136640 276762 136692 276768
rect 135352 250776 135404 250782
rect 135352 250718 135404 250724
rect 135260 3800 135312 3806
rect 135260 3742 135312 3748
rect 135364 3482 135392 250718
rect 136652 16574 136680 276762
rect 138032 16574 138060 283630
rect 139412 16574 139440 287710
rect 142160 263016 142212 263022
rect 142160 262958 142212 262964
rect 140780 247988 140832 247994
rect 140780 247930 140832 247936
rect 140792 16574 140820 247930
rect 136652 16546 137232 16574
rect 138032 16546 138888 16574
rect 139412 16546 139624 16574
rect 140792 16546 141280 16574
rect 136456 3800 136508 3806
rect 136456 3742 136508 3748
rect 135272 3454 135392 3482
rect 135272 480 135300 3454
rect 136468 480 136496 3742
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 16546
rect 138860 480 138888 16546
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 139596 354 139624 16546
rect 141252 480 141280 16546
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142172 354 142200 262958
rect 143552 480 143580 290566
rect 146300 286544 146352 286550
rect 146300 286486 146352 286492
rect 143632 268456 143684 268462
rect 143632 268398 143684 268404
rect 143644 16574 143672 268398
rect 144920 261656 144972 261662
rect 144920 261598 144972 261604
rect 144932 16574 144960 261598
rect 146312 16574 146340 286486
rect 150440 285184 150492 285190
rect 150440 285126 150492 285132
rect 147680 278248 147732 278254
rect 147680 278190 147732 278196
rect 147692 16574 147720 278190
rect 149060 264308 149112 264314
rect 149060 264250 149112 264256
rect 149072 16574 149100 264250
rect 150452 16574 150480 285126
rect 153200 283756 153252 283762
rect 153200 283698 153252 283704
rect 151820 270020 151872 270026
rect 151820 269962 151872 269968
rect 143644 16546 144776 16574
rect 144932 16546 145512 16574
rect 146312 16546 147168 16574
rect 147692 16546 147904 16574
rect 149072 16546 149560 16574
rect 150452 16546 150664 16574
rect 144748 480 144776 16546
rect 142406 354 142518 480
rect 142172 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 147140 480 147168 16546
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 149532 480 149560 16546
rect 150636 480 150664 16546
rect 151832 480 151860 269962
rect 151912 268524 151964 268530
rect 151912 268466 151964 268472
rect 151924 16574 151952 268466
rect 153212 16574 153240 283698
rect 157340 282396 157392 282402
rect 157340 282338 157392 282344
rect 154580 264376 154632 264382
rect 154580 264318 154632 264324
rect 154592 16574 154620 264318
rect 155960 252000 156012 252006
rect 155960 251942 156012 251948
rect 155972 16574 156000 251942
rect 157352 16574 157380 282338
rect 158720 261724 158772 261730
rect 158720 261666 158772 261672
rect 158732 16574 158760 261666
rect 151924 16546 153056 16574
rect 153212 16546 153792 16574
rect 154592 16546 155448 16574
rect 155972 16546 156184 16574
rect 157352 16546 157840 16574
rect 158732 16546 158944 16574
rect 153028 480 153056 16546
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 16546
rect 155420 480 155448 16546
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156156 354 156184 16546
rect 157812 480 157840 16546
rect 158916 480 158944 16546
rect 160112 11762 160140 300183
rect 161216 298654 161244 300084
rect 161204 298648 161256 298654
rect 161204 298590 161256 298596
rect 163792 298586 163820 300084
rect 163780 298580 163832 298586
rect 163780 298522 163832 298528
rect 161480 292052 161532 292058
rect 161480 291994 161532 292000
rect 160192 252068 160244 252074
rect 160192 252010 160244 252016
rect 160100 11756 160152 11762
rect 160100 11698 160152 11704
rect 160204 6914 160232 252010
rect 161492 16574 161520 291994
rect 162860 274168 162912 274174
rect 162860 274110 162912 274116
rect 162872 16574 162900 274110
rect 164252 16574 164280 300319
rect 166368 298110 166396 300084
rect 166356 298104 166408 298110
rect 166356 298046 166408 298052
rect 169864 298042 169892 306274
rect 170404 305856 170456 305862
rect 170404 305798 170456 305804
rect 170036 304632 170088 304638
rect 170036 304574 170088 304580
rect 169944 303476 169996 303482
rect 169944 303418 169996 303424
rect 169852 298036 169904 298042
rect 169852 297978 169904 297984
rect 169956 297770 169984 303418
rect 169944 297764 169996 297770
rect 169944 297706 169996 297712
rect 170048 297362 170076 304574
rect 170036 297356 170088 297362
rect 170036 297298 170088 297304
rect 168380 294772 168432 294778
rect 168380 294714 168432 294720
rect 165620 279676 165672 279682
rect 165620 279618 165672 279624
rect 165632 16574 165660 279618
rect 167000 271312 167052 271318
rect 167000 271254 167052 271260
rect 167012 16574 167040 271254
rect 161492 16546 162072 16574
rect 162872 16546 163728 16574
rect 164252 16546 164464 16574
rect 165632 16546 166120 16574
rect 167012 16546 167224 16574
rect 161296 11756 161348 11762
rect 161296 11698 161348 11704
rect 160112 6886 160232 6914
rect 160112 480 160140 6886
rect 161308 480 161336 11698
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 354 162072 16546
rect 163700 480 163728 16546
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164436 354 164464 16546
rect 166092 480 166120 16546
rect 167196 480 167224 16546
rect 168392 480 168420 294714
rect 169760 254924 169812 254930
rect 169760 254866 169812 254872
rect 168472 245200 168524 245206
rect 168472 245142 168524 245148
rect 168484 16574 168512 245142
rect 169772 16574 169800 254866
rect 168484 16546 169616 16574
rect 169772 16546 170352 16574
rect 169588 480 169616 16546
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170324 354 170352 16546
rect 170416 3534 170444 305798
rect 170494 303104 170550 303113
rect 170494 303039 170550 303048
rect 170508 3738 170536 303039
rect 170600 298110 170628 307090
rect 170588 298104 170640 298110
rect 170588 298046 170640 298052
rect 170496 3732 170548 3738
rect 170496 3674 170548 3680
rect 170404 3528 170456 3534
rect 170404 3470 170456 3476
rect 171152 3466 171180 345034
rect 171322 323232 171378 323241
rect 171322 323167 171378 323176
rect 171336 322998 171364 323167
rect 171324 322992 171376 322998
rect 171324 322934 171376 322940
rect 171506 320512 171562 320521
rect 171506 320447 171562 320456
rect 171520 320210 171548 320447
rect 171508 320204 171560 320210
rect 171508 320146 171560 320152
rect 171506 317792 171562 317801
rect 171506 317727 171562 317736
rect 171520 317490 171548 317727
rect 171508 317484 171560 317490
rect 171508 317426 171560 317432
rect 171416 307692 171468 307698
rect 171416 307634 171468 307640
rect 171428 306921 171456 307634
rect 171796 307630 171824 374410
rect 172334 369472 172390 369481
rect 172334 369407 172390 369416
rect 172348 368558 172376 369407
rect 172336 368552 172388 368558
rect 172336 368494 172388 368500
rect 172426 366752 172482 366761
rect 172426 366687 172482 366696
rect 172440 365770 172468 366687
rect 172428 365764 172480 365770
rect 172428 365706 172480 365712
rect 172334 364032 172390 364041
rect 172334 363967 172390 363976
rect 172348 362982 172376 363967
rect 172336 362976 172388 362982
rect 172336 362918 172388 362924
rect 171874 361312 171930 361321
rect 171874 361247 171930 361256
rect 171888 311302 171916 361247
rect 171966 355872 172022 355881
rect 171966 355807 172022 355816
rect 171876 311296 171928 311302
rect 171876 311238 171928 311244
rect 171980 310078 172008 355807
rect 172426 353152 172482 353161
rect 172426 353087 172482 353096
rect 172440 351966 172468 353087
rect 172428 351960 172480 351966
rect 172428 351902 172480 351908
rect 172426 347712 172482 347721
rect 172426 347647 172482 347656
rect 172440 346458 172468 347647
rect 172428 346452 172480 346458
rect 172428 346394 172480 346400
rect 172058 344992 172114 345001
rect 172058 344927 172114 344936
rect 172072 310865 172100 344927
rect 172150 342272 172206 342281
rect 172150 342207 172206 342216
rect 172058 310856 172114 310865
rect 172058 310791 172114 310800
rect 172164 310622 172192 342207
rect 172242 339552 172298 339561
rect 172242 339487 172298 339496
rect 172256 311234 172284 339487
rect 172426 336832 172482 336841
rect 172426 336767 172428 336776
rect 172480 336767 172482 336776
rect 172428 336738 172480 336744
rect 172426 334112 172482 334121
rect 172426 334047 172482 334056
rect 172440 334014 172468 334047
rect 172428 334008 172480 334014
rect 172428 333950 172480 333956
rect 172426 331392 172482 331401
rect 172426 331327 172482 331336
rect 172440 331294 172468 331327
rect 172428 331288 172480 331294
rect 172428 331230 172480 331236
rect 172334 328672 172390 328681
rect 172334 328607 172390 328616
rect 172348 311438 172376 328607
rect 172426 325952 172482 325961
rect 172426 325887 172482 325896
rect 172440 325718 172468 325887
rect 172428 325712 172480 325718
rect 172428 325654 172480 325660
rect 172426 315072 172482 315081
rect 172426 315007 172482 315016
rect 172440 314702 172468 315007
rect 172428 314696 172480 314702
rect 172428 314638 172480 314644
rect 172426 312352 172482 312361
rect 172426 312287 172482 312296
rect 172440 311914 172468 312287
rect 172428 311908 172480 311914
rect 172428 311850 172480 311856
rect 172336 311432 172388 311438
rect 172336 311374 172388 311380
rect 172244 311228 172296 311234
rect 172244 311170 172296 311176
rect 172152 310616 172204 310622
rect 172152 310558 172204 310564
rect 171968 310072 172020 310078
rect 171968 310014 172020 310020
rect 172242 309632 172298 309641
rect 172242 309567 172298 309576
rect 172256 309194 172284 309567
rect 172244 309188 172296 309194
rect 172244 309130 172296 309136
rect 171784 307624 171836 307630
rect 171784 307566 171836 307572
rect 173176 307018 173204 374818
rect 180064 374332 180116 374338
rect 180064 374274 180116 374280
rect 174544 373108 174596 373114
rect 174544 373050 174596 373056
rect 173256 373040 173308 373046
rect 173256 372982 173308 372988
rect 173268 308281 173296 372982
rect 173440 372972 173492 372978
rect 173440 372914 173492 372920
rect 173452 308961 173480 372914
rect 173438 308952 173494 308961
rect 173438 308887 173494 308896
rect 174556 308582 174584 373050
rect 174636 371680 174688 371686
rect 174636 371622 174688 371628
rect 174544 308576 174596 308582
rect 174544 308518 174596 308524
rect 174648 308378 174676 371622
rect 178684 345092 178736 345098
rect 178684 345034 178736 345040
rect 178696 311166 178724 345034
rect 178684 311160 178736 311166
rect 178684 311102 178736 311108
rect 174636 308372 174688 308378
rect 174636 308314 174688 308320
rect 173254 308272 173310 308281
rect 173254 308207 173310 308216
rect 180076 307494 180104 374274
rect 180064 307488 180116 307494
rect 180064 307430 180116 307436
rect 173164 307012 173216 307018
rect 173164 306954 173216 306960
rect 171414 306912 171470 306921
rect 171414 306847 171470 306856
rect 178040 305652 178092 305658
rect 178040 305594 178092 305600
rect 171692 305448 171744 305454
rect 171692 305390 171744 305396
rect 171704 297430 171732 305390
rect 172336 304972 172388 304978
rect 172336 304914 172388 304920
rect 171968 304564 172020 304570
rect 171968 304506 172020 304512
rect 171784 304360 171836 304366
rect 171784 304302 171836 304308
rect 171692 297424 171744 297430
rect 171692 297366 171744 297372
rect 171232 245268 171284 245274
rect 171232 245210 171284 245216
rect 171244 16574 171272 245210
rect 171244 16546 171732 16574
rect 171704 3482 171732 16546
rect 171796 3670 171824 304302
rect 171980 297566 172008 304506
rect 172244 304496 172296 304502
rect 172244 304438 172296 304444
rect 172256 297634 172284 304438
rect 172348 304201 172376 304914
rect 172334 304192 172390 304201
rect 172334 304127 172390 304136
rect 172428 302184 172480 302190
rect 172428 302126 172480 302132
rect 172440 301481 172468 302126
rect 172426 301472 172482 301481
rect 172426 301407 172482 301416
rect 172244 297628 172296 297634
rect 172244 297570 172296 297576
rect 171968 297560 172020 297566
rect 171968 297502 172020 297508
rect 176660 258868 176712 258874
rect 176660 258810 176712 258816
rect 173900 258732 173952 258738
rect 173900 258674 173952 258680
rect 172520 252136 172572 252142
rect 172520 252078 172572 252084
rect 172532 16574 172560 252078
rect 172532 16546 172744 16574
rect 171784 3664 171836 3670
rect 171784 3606 171836 3612
rect 171140 3460 171192 3466
rect 171704 3454 172008 3482
rect 171140 3402 171192 3408
rect 171980 480 172008 3454
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173912 354 173940 258674
rect 175280 246764 175332 246770
rect 175280 246706 175332 246712
rect 175292 16574 175320 246706
rect 175292 16546 175504 16574
rect 175476 480 175504 16546
rect 176672 11762 176700 258810
rect 176752 253564 176804 253570
rect 176752 253506 176804 253512
rect 176660 11756 176712 11762
rect 176660 11698 176712 11704
rect 176764 6914 176792 253506
rect 178052 16574 178080 305594
rect 189080 304292 189132 304298
rect 189080 304234 189132 304240
rect 184938 302968 184994 302977
rect 184938 302903 184994 302912
rect 182178 302832 182234 302841
rect 182178 302767 182234 302776
rect 181444 287904 181496 287910
rect 181444 287846 181496 287852
rect 180800 272740 180852 272746
rect 180800 272682 180852 272688
rect 180812 16574 180840 272682
rect 178052 16546 178632 16574
rect 180812 16546 181024 16574
rect 177856 11756 177908 11762
rect 177856 11698 177908 11704
rect 176672 6886 176792 6914
rect 176672 480 176700 6886
rect 177868 480 177896 11698
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 173134 -960 173246 326
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 180248 4140 180300 4146
rect 180248 4082 180300 4088
rect 180260 480 180288 4082
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 181456 4146 181484 287846
rect 181444 4140 181496 4146
rect 181444 4082 181496 4088
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 182192 354 182220 302767
rect 184952 11762 184980 302903
rect 187700 290692 187752 290698
rect 187700 290634 187752 290640
rect 185032 249416 185084 249422
rect 185032 249358 185084 249364
rect 184940 11756 184992 11762
rect 184940 11698 184992 11704
rect 185044 6914 185072 249358
rect 187712 16574 187740 290634
rect 188344 278316 188396 278322
rect 188344 278258 188396 278264
rect 187712 16546 188292 16574
rect 186136 11756 186188 11762
rect 186136 11698 186188 11704
rect 184952 6886 185072 6914
rect 183744 3664 183796 3670
rect 183744 3606 183796 3612
rect 183756 480 183784 3606
rect 184952 480 184980 6886
rect 186148 480 186176 11698
rect 187332 3528 187384 3534
rect 187332 3470 187384 3476
rect 188264 3482 188292 16546
rect 188356 3670 188384 278258
rect 189092 16574 189120 304234
rect 191840 265940 191892 265946
rect 191840 265882 191892 265888
rect 191852 16574 191880 265882
rect 192496 97986 192524 445878
rect 199384 444780 199436 444786
rect 199384 444722 199436 444728
rect 196716 443216 196768 443222
rect 196716 443158 196768 443164
rect 195980 305720 196032 305726
rect 195980 305662 196032 305668
rect 193220 301504 193272 301510
rect 193220 301446 193272 301452
rect 192484 97980 192536 97986
rect 192484 97922 192536 97928
rect 189092 16546 189304 16574
rect 191852 16546 192064 16574
rect 188344 3664 188396 3670
rect 188344 3606 188396 3612
rect 187344 480 187372 3470
rect 188264 3454 188568 3482
rect 188540 480 188568 3454
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189276 354 189304 16546
rect 190828 3460 190880 3466
rect 190828 3402 190880 3408
rect 190840 480 190868 3402
rect 192036 480 192064 16546
rect 193232 480 193260 301446
rect 193312 275596 193364 275602
rect 193312 275538 193364 275544
rect 193324 16574 193352 275538
rect 195992 16574 196020 305662
rect 196624 276888 196676 276894
rect 196624 276830 196676 276836
rect 193324 16546 194456 16574
rect 195992 16546 196572 16574
rect 194428 480 194456 16546
rect 195980 3800 196032 3806
rect 195980 3742 196032 3748
rect 195992 3534 196020 3742
rect 195980 3528 196032 3534
rect 195980 3470 196032 3476
rect 196544 3482 196572 16546
rect 196636 3806 196664 276830
rect 196728 202842 196756 443158
rect 198004 442128 198056 442134
rect 198004 442070 198056 442076
rect 197360 274236 197412 274242
rect 197360 274178 197412 274184
rect 196716 202836 196768 202842
rect 196716 202778 196768 202784
rect 197372 16574 197400 274178
rect 198016 150414 198044 442070
rect 198740 281036 198792 281042
rect 198740 280978 198792 280984
rect 198096 245336 198148 245342
rect 198096 245278 198148 245284
rect 198004 150408 198056 150414
rect 198004 150350 198056 150356
rect 197372 16546 197952 16574
rect 196624 3800 196676 3806
rect 196624 3742 196676 3748
rect 196544 3454 196848 3482
rect 195612 3052 195664 3058
rect 195612 2994 195664 3000
rect 195624 480 195652 2994
rect 196820 480 196848 3454
rect 197924 480 197952 16546
rect 198108 3058 198136 245278
rect 198096 3052 198148 3058
rect 198096 2994 198148 3000
rect 189694 354 189806 480
rect 189276 326 189806 354
rect 189694 -960 189806 326
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 280978
rect 199396 45558 199424 444722
rect 200764 442196 200816 442202
rect 200764 442138 200816 442144
rect 200120 307080 200172 307086
rect 200120 307022 200172 307028
rect 199384 45552 199436 45558
rect 199384 45494 199436 45500
rect 200132 16574 200160 307022
rect 200776 85542 200804 442138
rect 202880 293412 202932 293418
rect 202880 293354 202932 293360
rect 201500 272808 201552 272814
rect 201500 272750 201552 272756
rect 200764 85536 200816 85542
rect 200764 85478 200816 85484
rect 200132 16546 200344 16574
rect 200316 480 200344 16546
rect 201512 480 201540 272750
rect 201592 248056 201644 248062
rect 201592 247998 201644 248004
rect 201604 16574 201632 247998
rect 202892 16574 202920 293354
rect 203524 286612 203576 286618
rect 203524 286554 203576 286560
rect 201604 16546 202736 16574
rect 202892 16546 203472 16574
rect 202708 480 202736 16546
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203444 354 203472 16546
rect 203536 3466 203564 286554
rect 203628 189038 203656 445946
rect 205640 289332 205692 289338
rect 205640 289274 205692 289280
rect 203616 189032 203668 189038
rect 203616 188974 203668 188980
rect 205652 16574 205680 289274
rect 206296 137970 206324 446014
rect 217796 443698 217824 565082
rect 217888 478650 217916 700266
rect 217876 478644 217928 478650
rect 217876 478586 217928 478592
rect 217980 478582 218008 700334
rect 217968 478576 218020 478582
rect 217968 478518 218020 478524
rect 218072 464438 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 219348 700460 219400 700466
rect 219348 700402 219400 700408
rect 219070 512816 219126 512825
rect 219070 512751 219126 512760
rect 218978 508192 219034 508201
rect 218978 508127 219034 508136
rect 218886 488336 218942 488345
rect 218886 488271 218942 488280
rect 218900 465866 218928 488271
rect 218992 478310 219020 508127
rect 218980 478304 219032 478310
rect 218980 478246 219032 478252
rect 219084 475454 219112 512751
rect 219162 511048 219218 511057
rect 219162 510983 219218 510992
rect 219072 475448 219124 475454
rect 219072 475390 219124 475396
rect 219176 472802 219204 510983
rect 219254 509960 219310 509969
rect 219254 509895 219310 509904
rect 219164 472796 219216 472802
rect 219164 472738 219216 472744
rect 219268 468654 219296 509895
rect 219256 468648 219308 468654
rect 219256 468590 219308 468596
rect 218888 465860 218940 465866
rect 218888 465802 218940 465808
rect 218060 464432 218112 464438
rect 218060 464374 218112 464380
rect 219360 443766 219388 700402
rect 234632 565146 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 700466 267688 703520
rect 267648 700460 267700 700466
rect 267648 700402 267700 700408
rect 283852 700398 283880 703520
rect 283840 700392 283892 700398
rect 283840 700334 283892 700340
rect 300136 700330 300164 703520
rect 332520 700330 332548 703520
rect 348804 700398 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 348792 700392 348844 700398
rect 348792 700334 348844 700340
rect 358820 700392 358872 700398
rect 358820 700334 358872 700340
rect 300124 700324 300176 700330
rect 300124 700266 300176 700272
rect 332508 700324 332560 700330
rect 332508 700266 332560 700272
rect 357440 700324 357492 700330
rect 357440 700266 357492 700272
rect 234620 565140 234672 565146
rect 234620 565082 234672 565088
rect 269948 478644 270000 478650
rect 269948 478586 270000 478592
rect 268660 478508 268712 478514
rect 268660 478450 268712 478456
rect 256884 478236 256936 478242
rect 256884 478178 256936 478184
rect 238482 477320 238538 477329
rect 238482 477255 238538 477264
rect 238496 476814 238524 477255
rect 242806 477184 242862 477193
rect 242806 477119 242862 477128
rect 253754 477184 253810 477193
rect 253754 477119 253810 477128
rect 240046 476912 240102 476921
rect 240046 476847 240102 476856
rect 241426 476912 241482 476921
rect 241426 476847 241428 476856
rect 238484 476808 238536 476814
rect 237286 476776 237342 476785
rect 238484 476750 238536 476756
rect 237286 476711 237288 476720
rect 237340 476711 237342 476720
rect 239404 476740 239456 476746
rect 237288 476682 237340 476688
rect 239404 476682 239456 476688
rect 237194 476232 237250 476241
rect 237194 476167 237250 476176
rect 237208 454850 237236 476167
rect 239416 460358 239444 476682
rect 240060 476134 240088 476847
rect 241480 476847 241482 476856
rect 241428 476818 241480 476824
rect 242820 476678 242848 477119
rect 242808 476672 242860 476678
rect 242808 476614 242860 476620
rect 245566 476368 245622 476377
rect 245566 476303 245622 476312
rect 248234 476368 248290 476377
rect 248234 476303 248290 476312
rect 251086 476368 251142 476377
rect 251086 476303 251142 476312
rect 252374 476368 252430 476377
rect 252374 476303 252430 476312
rect 244186 476232 244242 476241
rect 244186 476167 244242 476176
rect 245474 476232 245530 476241
rect 245474 476167 245530 476176
rect 240048 476128 240100 476134
rect 240048 476070 240100 476076
rect 244200 463146 244228 476167
rect 244188 463140 244240 463146
rect 244188 463082 244240 463088
rect 239404 460352 239456 460358
rect 239404 460294 239456 460300
rect 237196 454844 237248 454850
rect 237196 454786 237248 454792
rect 245488 449682 245516 476167
rect 245580 449750 245608 476303
rect 246946 476232 247002 476241
rect 246946 476167 247002 476176
rect 246960 464506 246988 476167
rect 248248 468722 248276 476303
rect 248326 476232 248382 476241
rect 248326 476167 248382 476176
rect 249706 476232 249762 476241
rect 249706 476167 249762 476176
rect 250994 476232 251050 476241
rect 250994 476167 251050 476176
rect 248236 468716 248288 468722
rect 248236 468658 248288 468664
rect 246948 464500 247000 464506
rect 246948 464442 247000 464448
rect 248340 453626 248368 476167
rect 249720 463078 249748 476167
rect 249708 463072 249760 463078
rect 249708 463014 249760 463020
rect 251008 460426 251036 476167
rect 250996 460420 251048 460426
rect 250996 460362 251048 460368
rect 251100 457638 251128 476303
rect 252388 467362 252416 476303
rect 252466 476232 252522 476241
rect 252466 476167 252522 476176
rect 252376 467356 252428 467362
rect 252376 467298 252428 467304
rect 251088 457632 251140 457638
rect 251088 457574 251140 457580
rect 252284 456816 252336 456822
rect 252284 456758 252336 456764
rect 248328 453620 248380 453626
rect 248328 453562 248380 453568
rect 245568 449744 245620 449750
rect 245568 449686 245620 449692
rect 245476 449676 245528 449682
rect 245476 449618 245528 449624
rect 243726 445904 243782 445913
rect 235908 445868 235960 445874
rect 243726 445839 243782 445848
rect 235908 445810 235960 445816
rect 231124 444916 231176 444922
rect 231124 444858 231176 444864
rect 225604 444848 225656 444854
rect 225604 444790 225656 444796
rect 219348 443760 219400 443766
rect 219348 443702 219400 443708
rect 217784 443692 217836 443698
rect 217784 443634 217836 443640
rect 224224 443284 224276 443290
rect 224224 443226 224276 443232
rect 207664 440632 207716 440638
rect 207664 440574 207716 440580
rect 207020 304428 207072 304434
rect 207020 304370 207072 304376
rect 206284 137964 206336 137970
rect 206284 137906 206336 137912
rect 205652 16546 206232 16574
rect 203524 3460 203576 3466
rect 203524 3402 203576 3408
rect 205086 3360 205142 3369
rect 205086 3295 205142 3304
rect 205100 480 205128 3295
rect 206204 480 206232 16546
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 304370
rect 207676 71738 207704 440574
rect 224236 378826 224264 443226
rect 224224 378820 224276 378826
rect 224224 378762 224276 378768
rect 224224 351960 224276 351966
rect 224224 351902 224276 351908
rect 220084 346452 220136 346458
rect 220084 346394 220136 346400
rect 214838 308408 214894 308417
rect 214838 308343 214894 308352
rect 213644 305992 213696 305998
rect 213644 305934 213696 305940
rect 210976 305788 211028 305794
rect 210976 305730 211028 305736
rect 210792 301776 210844 301782
rect 210792 301718 210844 301724
rect 210608 300076 210660 300082
rect 210608 300018 210660 300024
rect 209780 296132 209832 296138
rect 209780 296074 209832 296080
rect 209688 295112 209740 295118
rect 209688 295054 209740 295060
rect 207664 71732 207716 71738
rect 207664 71674 207716 71680
rect 208584 4140 208636 4146
rect 208584 4082 208636 4088
rect 208596 480 208624 4082
rect 209700 3534 209728 295054
rect 209792 3670 209820 296074
rect 209872 250844 209924 250850
rect 209872 250786 209924 250792
rect 209780 3664 209832 3670
rect 209780 3606 209832 3612
rect 209688 3528 209740 3534
rect 209884 3482 209912 250786
rect 210620 189038 210648 300018
rect 210700 297424 210752 297430
rect 210700 297366 210752 297372
rect 210608 189032 210660 189038
rect 210608 188974 210660 188980
rect 210712 155446 210740 297366
rect 210700 155440 210752 155446
rect 210700 155382 210752 155388
rect 210804 155281 210832 301718
rect 210884 301572 210936 301578
rect 210884 301514 210936 301520
rect 210896 155514 210924 301514
rect 210988 155650 211016 305730
rect 212172 302932 212224 302938
rect 212172 302874 212224 302880
rect 211068 301844 211120 301850
rect 211068 301786 211120 301792
rect 210976 155644 211028 155650
rect 210976 155586 211028 155592
rect 210884 155508 210936 155514
rect 210884 155450 210936 155456
rect 210790 155272 210846 155281
rect 210790 155207 210846 155216
rect 211080 3738 211108 301786
rect 211712 301640 211764 301646
rect 211712 301582 211764 301588
rect 211160 283824 211212 283830
rect 211160 283766 211212 283772
rect 211172 16574 211200 283766
rect 211724 158778 211752 301582
rect 211986 300520 212042 300529
rect 211986 300455 212042 300464
rect 211804 271380 211856 271386
rect 211804 271322 211856 271328
rect 211712 158772 211764 158778
rect 211712 158714 211764 158720
rect 211172 16546 211752 16574
rect 211068 3732 211120 3738
rect 211068 3674 211120 3680
rect 210976 3664 211028 3670
rect 210976 3606 211028 3612
rect 209688 3470 209740 3476
rect 209792 3454 209912 3482
rect 209792 480 209820 3454
rect 210988 480 211016 3606
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 16546
rect 211816 4146 211844 271322
rect 211896 246832 211948 246838
rect 211896 246774 211948 246780
rect 211804 4140 211856 4146
rect 211804 4082 211856 4088
rect 211908 3602 211936 246774
rect 212000 158642 212028 300455
rect 212078 297392 212134 297401
rect 212078 297327 212134 297336
rect 211988 158636 212040 158642
rect 211988 158578 212040 158584
rect 212092 155854 212120 297327
rect 212184 159458 212212 302874
rect 212448 301980 212500 301986
rect 212448 301922 212500 301928
rect 212264 301912 212316 301918
rect 212264 301854 212316 301860
rect 212172 159452 212224 159458
rect 212172 159394 212224 159400
rect 212080 155848 212132 155854
rect 212080 155790 212132 155796
rect 212276 155310 212304 301854
rect 212356 297356 212408 297362
rect 212356 297298 212408 297304
rect 212264 155304 212316 155310
rect 212264 155246 212316 155252
rect 212368 4146 212396 297298
rect 212356 4140 212408 4146
rect 212356 4082 212408 4088
rect 212460 3602 212488 301922
rect 213460 297764 213512 297770
rect 213460 297706 213512 297712
rect 213366 297664 213422 297673
rect 213366 297599 213422 297608
rect 213184 297560 213236 297566
rect 213184 297502 213236 297508
rect 212540 261792 212592 261798
rect 212540 261734 212592 261740
rect 212552 16574 212580 261734
rect 213196 158710 213224 297502
rect 213276 294840 213328 294846
rect 213276 294782 213328 294788
rect 213184 158704 213236 158710
rect 213184 158646 213236 158652
rect 213288 155242 213316 294782
rect 213380 158506 213408 297599
rect 213368 158500 213420 158506
rect 213368 158442 213420 158448
rect 213472 155582 213500 297706
rect 213550 297528 213606 297537
rect 213550 297463 213606 297472
rect 213564 155786 213592 297463
rect 213656 159662 213684 305934
rect 214656 303612 214708 303618
rect 214656 303554 214708 303560
rect 214564 303136 214616 303142
rect 214564 303078 214616 303084
rect 214472 297696 214524 297702
rect 214472 297638 214524 297644
rect 213828 297628 213880 297634
rect 213828 297570 213880 297576
rect 213736 297492 213788 297498
rect 213736 297434 213788 297440
rect 213644 159656 213696 159662
rect 213644 159598 213696 159604
rect 213552 155780 213604 155786
rect 213552 155722 213604 155728
rect 213460 155576 213512 155582
rect 213460 155518 213512 155524
rect 213276 155236 213328 155242
rect 213276 155178 213328 155184
rect 212552 16546 213408 16574
rect 211896 3596 211948 3602
rect 211896 3538 211948 3544
rect 212448 3596 212500 3602
rect 212448 3538 212500 3544
rect 213380 480 213408 16546
rect 213748 4010 213776 297434
rect 213840 4078 213868 297570
rect 214380 294908 214432 294914
rect 214380 294850 214432 294856
rect 214392 195702 214420 294850
rect 214380 195696 214432 195702
rect 214380 195638 214432 195644
rect 214484 159594 214512 297638
rect 214472 159588 214524 159594
rect 214472 159530 214524 159536
rect 214576 158234 214604 303078
rect 214564 158228 214616 158234
rect 214564 158170 214616 158176
rect 214668 157865 214696 303554
rect 214748 303340 214800 303346
rect 214748 303282 214800 303288
rect 214760 157962 214788 303282
rect 214852 159390 214880 308343
rect 220096 307426 220124 346394
rect 220084 307420 220136 307426
rect 220084 307362 220136 307368
rect 224236 307290 224264 351902
rect 224224 307284 224276 307290
rect 224224 307226 224276 307232
rect 215208 306264 215260 306270
rect 215208 306206 215260 306212
rect 215024 303204 215076 303210
rect 215024 303146 215076 303152
rect 214932 295044 214984 295050
rect 214932 294986 214984 294992
rect 214840 159384 214892 159390
rect 214840 159326 214892 159332
rect 214748 157956 214800 157962
rect 214748 157898 214800 157904
rect 214654 157856 214710 157865
rect 214654 157791 214710 157800
rect 213828 4072 213880 4078
rect 213828 4014 213880 4020
rect 213736 4004 213788 4010
rect 213736 3946 213788 3952
rect 214944 3874 214972 294986
rect 214932 3868 214984 3874
rect 214932 3810 214984 3816
rect 214470 3496 214526 3505
rect 214470 3431 214526 3440
rect 214484 480 214512 3431
rect 215036 3398 215064 303146
rect 215116 302864 215168 302870
rect 215116 302806 215168 302812
rect 215024 3392 215076 3398
rect 215024 3334 215076 3340
rect 215128 3330 215156 302806
rect 215220 3369 215248 306206
rect 218980 306196 219032 306202
rect 218980 306138 219032 306144
rect 216404 306128 216456 306134
rect 216404 306070 216456 306076
rect 216312 306060 216364 306066
rect 216312 306002 216364 306008
rect 215944 303544 215996 303550
rect 215944 303486 215996 303492
rect 215852 302796 215904 302802
rect 215852 302738 215904 302744
rect 215760 294976 215812 294982
rect 215760 294918 215812 294924
rect 215772 193186 215800 294918
rect 215760 193180 215812 193186
rect 215760 193122 215812 193128
rect 215864 157826 215892 302738
rect 215956 158574 215984 303486
rect 216036 303272 216088 303278
rect 216036 303214 216088 303220
rect 215944 158568 215996 158574
rect 215944 158510 215996 158516
rect 216048 158370 216076 303214
rect 216220 302116 216272 302122
rect 216220 302058 216272 302064
rect 216128 302048 216180 302054
rect 216128 301990 216180 301996
rect 216036 158364 216088 158370
rect 216036 158306 216088 158312
rect 215852 157820 215904 157826
rect 215852 157762 215904 157768
rect 216140 155038 216168 301990
rect 216232 155718 216260 302058
rect 216324 158098 216352 306002
rect 216416 158302 216444 306070
rect 216588 305924 216640 305930
rect 216588 305866 216640 305872
rect 216496 302728 216548 302734
rect 216496 302670 216548 302676
rect 216404 158296 216456 158302
rect 216404 158238 216456 158244
rect 216312 158092 216364 158098
rect 216312 158034 216364 158040
rect 216220 155712 216272 155718
rect 216220 155654 216272 155660
rect 216128 155032 216180 155038
rect 216128 154974 216180 154980
rect 215666 3496 215722 3505
rect 215666 3431 215722 3440
rect 215206 3360 215262 3369
rect 215116 3324 215168 3330
rect 215206 3295 215262 3304
rect 215116 3266 215168 3272
rect 215680 480 215708 3431
rect 216508 3194 216536 302670
rect 216600 3466 216628 305866
rect 218888 305516 218940 305522
rect 218888 305458 218940 305464
rect 217968 303408 218020 303414
rect 217968 303350 218020 303356
rect 217784 299940 217836 299946
rect 217784 299882 217836 299888
rect 217692 287836 217744 287842
rect 217692 287778 217744 287784
rect 217324 267232 217376 267238
rect 217324 267174 217376 267180
rect 217140 256352 217192 256358
rect 217140 256294 217192 256300
rect 217152 192817 217180 256294
rect 217232 249348 217284 249354
rect 217232 249290 217284 249296
rect 217138 192808 217194 192817
rect 217138 192743 217194 192752
rect 216680 189032 216732 189038
rect 216680 188974 216732 188980
rect 216692 188193 216720 188974
rect 216678 188184 216734 188193
rect 216678 188119 216734 188128
rect 217244 168065 217272 249290
rect 217336 195945 217364 267174
rect 217600 258800 217652 258806
rect 217600 258742 217652 258748
rect 217416 254856 217468 254862
rect 217416 254798 217468 254804
rect 217322 195936 217378 195945
rect 217322 195871 217378 195880
rect 217324 195696 217376 195702
rect 217324 195638 217376 195644
rect 217230 168056 217286 168065
rect 217230 167991 217286 168000
rect 217336 3670 217364 195638
rect 217428 168337 217456 254798
rect 217508 243568 217560 243574
rect 217508 243510 217560 243516
rect 217414 168328 217470 168337
rect 217414 168263 217470 168272
rect 217520 155174 217548 243510
rect 217612 169969 217640 258742
rect 217704 196897 217732 287778
rect 217690 196888 217746 196897
rect 217690 196823 217746 196832
rect 217796 193769 217824 299882
rect 217876 297288 217928 297294
rect 217876 297230 217928 297236
rect 217782 193760 217838 193769
rect 217782 193695 217838 193704
rect 217598 169960 217654 169969
rect 217598 169895 217654 169904
rect 217888 159526 217916 297230
rect 217876 159520 217928 159526
rect 217876 159462 217928 159468
rect 217980 158166 218008 303350
rect 218428 301708 218480 301714
rect 218428 301650 218480 301656
rect 218440 191049 218468 301650
rect 218796 297220 218848 297226
rect 218796 297162 218848 297168
rect 218612 257644 218664 257650
rect 218612 257586 218664 257592
rect 218520 253496 218572 253502
rect 218520 253438 218572 253444
rect 218426 191040 218482 191049
rect 218426 190975 218482 190984
rect 218532 189961 218560 253438
rect 218624 193225 218652 257586
rect 218610 193216 218666 193225
rect 218610 193151 218666 193160
rect 218704 193180 218756 193186
rect 218704 193122 218756 193128
rect 218518 189952 218574 189961
rect 218518 189887 218574 189896
rect 217968 158160 218020 158166
rect 217968 158102 218020 158108
rect 217508 155168 217560 155174
rect 217508 155110 217560 155116
rect 218716 3806 218744 193122
rect 218808 155378 218836 297162
rect 218900 157894 218928 305458
rect 218992 158030 219020 306138
rect 219072 305584 219124 305590
rect 219072 305526 219124 305532
rect 219084 158438 219112 305526
rect 219164 303068 219216 303074
rect 219164 303010 219216 303016
rect 219072 158432 219124 158438
rect 219072 158374 219124 158380
rect 218980 158024 219032 158030
rect 218980 157966 219032 157972
rect 218888 157888 218940 157894
rect 218888 157830 218940 157836
rect 218796 155372 218848 155378
rect 218796 155314 218848 155320
rect 219176 155106 219204 303010
rect 219348 295180 219400 295186
rect 219348 295122 219400 295128
rect 219256 243636 219308 243642
rect 219256 243578 219308 243584
rect 219164 155100 219216 155106
rect 219164 155042 219216 155048
rect 219268 6914 219296 243578
rect 219176 6886 219296 6914
rect 218704 3800 218756 3806
rect 218704 3742 218756 3748
rect 217324 3664 217376 3670
rect 217324 3606 217376 3612
rect 219176 3534 219204 6886
rect 219360 3942 219388 295122
rect 225616 267714 225644 444790
rect 229744 443352 229796 443358
rect 229744 443294 229796 443300
rect 229756 377466 229784 443294
rect 231136 398818 231164 444858
rect 234618 444680 234674 444689
rect 234618 444615 234674 444624
rect 233976 443080 234028 443086
rect 232686 443048 232742 443057
rect 233976 443022 234028 443028
rect 232686 442983 232742 442992
rect 231216 442536 231268 442542
rect 231216 442478 231268 442484
rect 231228 411262 231256 442478
rect 232700 441524 232728 442983
rect 233332 441652 233384 441658
rect 233332 441594 233384 441600
rect 233344 441524 233372 441594
rect 233988 441524 234016 443022
rect 234632 441524 234660 444615
rect 235262 443320 235318 443329
rect 235262 443255 235318 443264
rect 235276 441524 235304 443255
rect 235920 441524 235948 445810
rect 237838 445768 237894 445777
rect 237838 445703 237894 445712
rect 236550 444408 236606 444417
rect 236550 444343 236606 444352
rect 236564 441524 236592 444343
rect 237196 441720 237248 441726
rect 237196 441662 237248 441668
rect 237208 441524 237236 441662
rect 237852 441524 237880 445703
rect 238574 444544 238630 444553
rect 238574 444479 238630 444488
rect 238588 441524 238616 444479
rect 239220 443896 239272 443902
rect 239220 443838 239272 443844
rect 239232 441524 239260 443838
rect 241152 443556 241204 443562
rect 241152 443498 241204 443504
rect 239862 443184 239918 443193
rect 239862 443119 239918 443128
rect 239876 441524 239904 443119
rect 241164 441524 241192 443498
rect 241796 441924 241848 441930
rect 241796 441866 241848 441872
rect 241808 441524 241836 441866
rect 242440 441788 242492 441794
rect 242440 441730 242492 441736
rect 242452 441524 242480 441730
rect 243082 441688 243138 441697
rect 243082 441623 243138 441632
rect 243096 441524 243124 441623
rect 243740 441524 243768 445839
rect 249708 444712 249760 444718
rect 249708 444654 249760 444660
rect 244464 444440 244516 444446
rect 244464 444382 244516 444388
rect 244476 441524 244504 444382
rect 245752 444168 245804 444174
rect 245752 444110 245804 444116
rect 245108 443488 245160 443494
rect 245108 443430 245160 443436
rect 245120 441524 245148 443430
rect 245764 441524 245792 444110
rect 246396 443624 246448 443630
rect 246396 443566 246448 443572
rect 246408 441524 246436 443566
rect 248328 443420 248380 443426
rect 248328 443362 248380 443368
rect 246948 443080 247000 443086
rect 246948 443022 247000 443028
rect 246960 442241 246988 443022
rect 246946 442232 247002 442241
rect 246946 442167 247002 442176
rect 247040 441992 247092 441998
rect 247040 441934 247092 441940
rect 247052 441524 247080 441934
rect 248340 441524 248368 443362
rect 248972 442060 249024 442066
rect 248972 442002 249024 442008
rect 248984 441524 249012 442002
rect 249720 441524 249748 444654
rect 250352 443148 250404 443154
rect 250352 443090 250404 443096
rect 250364 441524 250392 443090
rect 250996 443012 251048 443018
rect 250996 442954 251048 442960
rect 251008 441524 251036 442954
rect 252296 441524 252324 456758
rect 252480 447982 252508 476167
rect 253768 474230 253796 477119
rect 256606 477048 256662 477057
rect 256606 476983 256662 476992
rect 256620 476474 256648 476983
rect 256608 476468 256660 476474
rect 256608 476410 256660 476416
rect 253846 476232 253902 476241
rect 253846 476167 253902 476176
rect 255226 476232 255282 476241
rect 255226 476167 255282 476176
rect 256514 476232 256570 476241
rect 256514 476167 256570 476176
rect 253756 474224 253808 474230
rect 253756 474166 253808 474172
rect 252928 472728 252980 472734
rect 252928 472670 252980 472676
rect 252468 447976 252520 447982
rect 252468 447918 252520 447924
rect 252560 443964 252612 443970
rect 252560 443906 252612 443912
rect 252572 441182 252600 443906
rect 252940 441524 252968 472670
rect 253204 470620 253256 470626
rect 253204 470562 253256 470568
rect 253216 443358 253244 470562
rect 253860 470082 253888 476167
rect 254860 474088 254912 474094
rect 254860 474030 254912 474036
rect 253848 470076 253900 470082
rect 253848 470018 253900 470024
rect 254216 450628 254268 450634
rect 254216 450570 254268 450576
rect 253204 443352 253256 443358
rect 253204 443294 253256 443300
rect 253572 443352 253624 443358
rect 253572 443294 253624 443300
rect 253584 441524 253612 443294
rect 254228 441524 254256 450570
rect 254872 441524 254900 474030
rect 255240 470014 255268 476167
rect 255596 475380 255648 475386
rect 255596 475322 255648 475328
rect 255228 470008 255280 470014
rect 255228 469950 255280 469956
rect 255608 441524 255636 475322
rect 256528 457570 256556 476167
rect 256516 457564 256568 457570
rect 256516 457506 256568 457512
rect 256240 451988 256292 451994
rect 256240 451930 256292 451936
rect 256252 441524 256280 451930
rect 256896 441524 256924 478178
rect 259366 476776 259422 476785
rect 259366 476711 259422 476720
rect 257986 476232 258042 476241
rect 257986 476167 258042 476176
rect 259274 476232 259330 476241
rect 259274 476167 259330 476176
rect 258000 448050 258028 476167
rect 259288 472870 259316 476167
rect 259276 472864 259328 472870
rect 259276 472806 259328 472812
rect 258816 465792 258868 465798
rect 258816 465734 258868 465740
rect 258172 453348 258224 453354
rect 258172 453290 258224 453296
rect 257988 448044 258040 448050
rect 257988 447986 258040 447992
rect 257528 446412 257580 446418
rect 257528 446354 257580 446360
rect 257540 441524 257568 446354
rect 258184 441524 258212 453290
rect 258828 441524 258856 465734
rect 259380 458998 259408 476711
rect 266266 476640 266322 476649
rect 266266 476575 266322 476584
rect 266280 476542 266308 476575
rect 266268 476536 266320 476542
rect 262126 476504 262182 476513
rect 266268 476478 266320 476484
rect 262126 476439 262182 476448
rect 262140 476406 262168 476439
rect 262128 476400 262180 476406
rect 260654 476368 260710 476377
rect 262128 476342 262180 476348
rect 264794 476368 264850 476377
rect 260654 476303 260710 476312
rect 264794 476303 264850 476312
rect 267646 476368 267702 476377
rect 267646 476303 267702 476312
rect 259368 458992 259420 458998
rect 259368 458934 259420 458940
rect 260668 456142 260696 476303
rect 260746 476232 260802 476241
rect 260746 476167 260802 476176
rect 262034 476232 262090 476241
rect 262034 476167 262090 476176
rect 263506 476232 263562 476241
rect 263506 476167 263562 476176
rect 260656 456136 260708 456142
rect 260656 456078 260708 456084
rect 260104 454776 260156 454782
rect 260104 454718 260156 454724
rect 259460 446480 259512 446486
rect 259460 446422 259512 446428
rect 259472 441524 259500 446422
rect 260116 441524 260144 454718
rect 260760 450702 260788 476167
rect 261484 469940 261536 469946
rect 261484 469882 261536 469888
rect 260840 463004 260892 463010
rect 260840 462946 260892 462952
rect 260748 450696 260800 450702
rect 260748 450638 260800 450644
rect 260852 441524 260880 462946
rect 261496 441524 261524 469882
rect 262048 461786 262076 476167
rect 262772 467220 262824 467226
rect 262772 467162 262824 467168
rect 262036 461780 262088 461786
rect 262036 461722 262088 461728
rect 262128 456068 262180 456074
rect 262128 456010 262180 456016
rect 262140 441524 262168 456010
rect 262784 441524 262812 467162
rect 263520 449410 263548 476167
rect 264808 471442 264836 476303
rect 264886 476232 264942 476241
rect 264886 476167 264942 476176
rect 266174 476232 266230 476241
rect 266174 476167 266230 476176
rect 267554 476232 267610 476241
rect 267554 476167 267610 476176
rect 264796 471436 264848 471442
rect 264796 471378 264848 471384
rect 264704 468580 264756 468586
rect 264704 468522 264756 468528
rect 264060 458856 264112 458862
rect 264060 458798 264112 458804
rect 263508 449404 263560 449410
rect 263508 449346 263560 449352
rect 263416 446616 263468 446622
rect 263416 446558 263468 446564
rect 263428 441524 263456 446558
rect 264072 441524 264100 458798
rect 264716 441524 264744 468522
rect 264900 449546 264928 476167
rect 265992 460284 266044 460290
rect 265992 460226 266044 460232
rect 264888 449540 264940 449546
rect 264888 449482 264940 449488
rect 265348 446684 265400 446690
rect 265348 446626 265400 446632
rect 265360 441524 265388 446626
rect 266004 441524 266032 460226
rect 266188 449614 266216 476167
rect 266728 464364 266780 464370
rect 266728 464306 266780 464312
rect 266176 449608 266228 449614
rect 266176 449550 266228 449556
rect 266740 441524 266768 464306
rect 267568 449206 267596 476167
rect 267660 449478 267688 476303
rect 268016 461712 268068 461718
rect 268016 461654 268068 461660
rect 267648 449472 267700 449478
rect 267648 449414 267700 449420
rect 267556 449200 267608 449206
rect 267556 449142 267608 449148
rect 267372 446752 267424 446758
rect 267372 446694 267424 446700
rect 267384 441524 267412 446694
rect 268028 441524 268056 461654
rect 268568 443012 268620 443018
rect 268568 442954 268620 442960
rect 268580 442270 268608 442954
rect 268568 442264 268620 442270
rect 268568 442206 268620 442212
rect 268672 441524 268700 478450
rect 269304 478440 269356 478446
rect 269304 478382 269356 478388
rect 268934 476368 268990 476377
rect 268934 476303 268990 476312
rect 268948 466002 268976 476303
rect 269026 476232 269082 476241
rect 269026 476167 269082 476176
rect 268936 465996 268988 466002
rect 268936 465938 268988 465944
rect 269040 449342 269068 476167
rect 269028 449336 269080 449342
rect 269028 449278 269080 449284
rect 269028 443080 269080 443086
rect 269028 443022 269080 443028
rect 269040 442338 269068 443022
rect 269028 442332 269080 442338
rect 269028 442274 269080 442280
rect 269316 441524 269344 478382
rect 269960 441524 269988 478586
rect 271236 478576 271288 478582
rect 271236 478518 271288 478524
rect 270406 476232 270462 476241
rect 270406 476167 270462 476176
rect 270420 449274 270448 476167
rect 270408 449268 270460 449274
rect 270408 449210 270460 449216
rect 270592 443760 270644 443766
rect 270592 443702 270644 443708
rect 270604 441524 270632 443702
rect 271248 441524 271276 478518
rect 357452 478514 357480 700266
rect 358084 510672 358136 510678
rect 358084 510614 358136 510620
rect 357440 478508 357492 478514
rect 357440 478450 357492 478456
rect 308588 478372 308640 478378
rect 308588 478314 308640 478320
rect 282368 478168 282420 478174
rect 282368 478110 282420 478116
rect 271786 476640 271842 476649
rect 271786 476575 271788 476584
rect 271840 476575 271842 476584
rect 271788 476546 271840 476552
rect 274546 476504 274602 476513
rect 274546 476439 274602 476448
rect 274454 476368 274510 476377
rect 274454 476303 274510 476312
rect 271694 476232 271750 476241
rect 271694 476167 271750 476176
rect 273166 476232 273222 476241
rect 273166 476167 273222 476176
rect 274362 476232 274418 476241
rect 274362 476167 274418 476176
rect 271708 453490 271736 476167
rect 272616 456204 272668 456210
rect 272616 456146 272668 456152
rect 271696 453484 271748 453490
rect 271696 453426 271748 453432
rect 271972 443692 272024 443698
rect 271972 443634 272024 443640
rect 271984 441524 272012 443634
rect 272628 441524 272656 456146
rect 273180 452130 273208 476167
rect 273260 464432 273312 464438
rect 273260 464374 273312 464380
rect 273168 452124 273220 452130
rect 273168 452066 273220 452072
rect 273272 441524 273300 464374
rect 273904 453416 273956 453422
rect 273904 453358 273956 453364
rect 273916 441524 273944 453358
rect 274376 447914 274404 476167
rect 274468 464438 274496 476303
rect 274560 475522 274588 476439
rect 277306 476368 277362 476377
rect 277306 476303 277362 476312
rect 278594 476368 278650 476377
rect 278594 476303 278650 476312
rect 275926 476232 275982 476241
rect 275926 476167 275982 476176
rect 277214 476232 277270 476241
rect 277214 476167 277270 476176
rect 274548 475516 274600 475522
rect 274548 475458 274600 475464
rect 275940 472666 275968 476167
rect 275192 472660 275244 472666
rect 275192 472602 275244 472608
rect 275928 472660 275980 472666
rect 275928 472602 275980 472608
rect 274456 464432 274508 464438
rect 274456 464374 274508 464380
rect 274548 458924 274600 458930
rect 274548 458866 274600 458872
rect 274364 447908 274416 447914
rect 274364 447850 274416 447856
rect 274560 441524 274588 458866
rect 274732 443556 274784 443562
rect 274732 443498 274784 443504
rect 274640 443012 274692 443018
rect 274640 442954 274692 442960
rect 274652 442474 274680 442954
rect 274640 442468 274692 442474
rect 274640 442410 274692 442416
rect 274744 442338 274772 443498
rect 274732 442332 274784 442338
rect 274732 442274 274784 442280
rect 275204 441524 275232 472602
rect 277228 465934 277256 476167
rect 277216 465928 277268 465934
rect 277216 465870 277268 465876
rect 276480 461644 276532 461650
rect 276480 461586 276532 461592
rect 275836 451920 275888 451926
rect 275836 451862 275888 451868
rect 275848 441524 275876 451862
rect 276112 443420 276164 443426
rect 276112 443362 276164 443368
rect 252560 441176 252612 441182
rect 252560 441118 252612 441124
rect 276124 441046 276152 443362
rect 276492 441524 276520 461586
rect 277320 450566 277348 476303
rect 278608 460222 278636 476303
rect 278686 476232 278742 476241
rect 278686 476167 278742 476176
rect 280066 476232 280122 476241
rect 280066 476167 280122 476176
rect 281446 476232 281502 476241
rect 281446 476167 281502 476176
rect 278504 460216 278556 460222
rect 278504 460158 278556 460164
rect 278596 460216 278648 460222
rect 278596 460158 278648 460164
rect 277860 454708 277912 454714
rect 277860 454650 277912 454656
rect 277124 450560 277176 450566
rect 277124 450502 277176 450508
rect 277308 450560 277360 450566
rect 277308 450502 277360 450508
rect 277136 441524 277164 450502
rect 277400 443624 277452 443630
rect 277400 443566 277452 443572
rect 277412 441046 277440 443566
rect 277872 441524 277900 454650
rect 278516 441524 278544 460158
rect 278700 456210 278728 476167
rect 279792 465724 279844 465730
rect 279792 465666 279844 465672
rect 279148 456272 279200 456278
rect 279148 456214 279200 456220
rect 278688 456204 278740 456210
rect 278688 456146 278740 456152
rect 279160 441524 279188 456214
rect 279516 443420 279568 443426
rect 279516 443362 279568 443368
rect 279528 442406 279556 443362
rect 279516 442400 279568 442406
rect 279516 442342 279568 442348
rect 279804 441524 279832 465666
rect 280080 454714 280108 476167
rect 281080 459060 281132 459066
rect 281080 459002 281132 459008
rect 280436 457496 280488 457502
rect 280436 457438 280488 457444
rect 280068 454708 280120 454714
rect 280068 454650 280120 454656
rect 280448 441524 280476 457438
rect 281092 441524 281120 459002
rect 281460 458930 281488 476167
rect 281724 467152 281776 467158
rect 281724 467094 281776 467100
rect 281448 458924 281500 458930
rect 281448 458866 281500 458872
rect 281736 441524 281764 467094
rect 282380 441524 282408 478110
rect 284206 476232 284262 476241
rect 284206 476167 284262 476176
rect 286506 476232 286562 476241
rect 286506 476167 286562 476176
rect 288346 476232 288402 476241
rect 288346 476167 288402 476176
rect 291106 476232 291162 476241
rect 291106 476167 291162 476176
rect 293866 476232 293922 476241
rect 293866 476167 293922 476176
rect 296626 476232 296682 476241
rect 296626 476167 296682 476176
rect 299386 476232 299442 476241
rect 299386 476167 299442 476176
rect 302146 476232 302202 476241
rect 302146 476167 302202 476176
rect 303526 476232 303582 476241
rect 303526 476167 303582 476176
rect 306286 476232 306342 476241
rect 306286 476167 306342 476176
rect 283748 468512 283800 468518
rect 283748 468454 283800 468460
rect 283012 453552 283064 453558
rect 283012 453494 283064 453500
rect 282920 443896 282972 443902
rect 282920 443838 282972 443844
rect 282932 442406 282960 443838
rect 282920 442400 282972 442406
rect 282920 442342 282972 442348
rect 283024 441524 283052 453494
rect 283760 441524 283788 468454
rect 284220 451926 284248 476167
rect 284392 474020 284444 474026
rect 284392 473962 284444 473968
rect 284208 451920 284260 451926
rect 284208 451862 284260 451868
rect 284404 441524 284432 473962
rect 286520 471306 286548 476167
rect 287612 474768 287664 474774
rect 287612 474710 287664 474716
rect 286324 471300 286376 471306
rect 286324 471242 286376 471248
rect 286508 471300 286560 471306
rect 286508 471242 286560 471248
rect 285680 469872 285732 469878
rect 285680 469814 285732 469820
rect 285036 461848 285088 461854
rect 285036 461790 285088 461796
rect 285048 441524 285076 461790
rect 285692 441524 285720 469814
rect 286336 441524 286364 471242
rect 286968 452056 287020 452062
rect 286968 451998 287020 452004
rect 286980 441524 287008 451998
rect 287624 441524 287652 474710
rect 288360 469878 288388 476167
rect 288348 469872 288400 469878
rect 288348 469814 288400 469820
rect 288992 462392 289044 462398
rect 288992 462334 289044 462340
rect 288256 446548 288308 446554
rect 288256 446490 288308 446496
rect 288268 441524 288296 446490
rect 288348 443488 288400 443494
rect 288348 443430 288400 443436
rect 288360 442474 288388 443430
rect 288348 442468 288400 442474
rect 288348 442410 288400 442416
rect 289004 441524 289032 462334
rect 291120 461650 291148 476167
rect 291844 465996 291896 466002
rect 291844 465938 291896 465944
rect 291108 461644 291160 461650
rect 291108 461586 291160 461592
rect 290280 444916 290332 444922
rect 290280 444858 290332 444864
rect 289636 444508 289688 444514
rect 289636 444450 289688 444456
rect 289648 441524 289676 444450
rect 290292 441524 290320 444858
rect 291568 444644 291620 444650
rect 291568 444586 291620 444592
rect 290924 442536 290976 442542
rect 290924 442478 290976 442484
rect 290936 441524 290964 442478
rect 291580 441524 291608 444586
rect 291856 443766 291884 465938
rect 293880 463214 293908 476167
rect 294604 472864 294656 472870
rect 294604 472806 294656 472812
rect 293868 463208 293920 463214
rect 293868 463150 293920 463156
rect 293500 444576 293552 444582
rect 293500 444518 293552 444524
rect 291844 443760 291896 443766
rect 291844 443702 291896 443708
rect 292856 443284 292908 443290
rect 292856 443226 292908 443232
rect 292212 443080 292264 443086
rect 292212 443022 292264 443028
rect 292224 441524 292252 443022
rect 292868 441524 292896 443226
rect 293512 441524 293540 444518
rect 294616 443902 294644 472806
rect 295984 471436 296036 471442
rect 295984 471378 296036 471384
rect 295524 444848 295576 444854
rect 295524 444790 295576 444796
rect 294604 443896 294656 443902
rect 294604 443838 294656 443844
rect 294880 443828 294932 443834
rect 294880 443770 294932 443776
rect 294144 443012 294196 443018
rect 294144 442954 294196 442960
rect 294156 441524 294184 442954
rect 294892 441524 294920 443770
rect 295536 441524 295564 444790
rect 295996 443834 296024 471378
rect 296640 468518 296668 476167
rect 296628 468512 296680 468518
rect 296628 468454 296680 468460
rect 299400 465730 299428 476167
rect 299388 465724 299440 465730
rect 299388 465666 299440 465672
rect 302160 453422 302188 476167
rect 302148 453416 302200 453422
rect 302148 453358 302200 453364
rect 300124 446072 300176 446078
rect 300124 446014 300176 446020
rect 298100 446004 298152 446010
rect 298100 445946 298152 445952
rect 296812 445800 296864 445806
rect 296812 445742 296864 445748
rect 295984 443828 296036 443834
rect 295984 443770 296036 443776
rect 296168 443420 296220 443426
rect 296168 443362 296220 443368
rect 296180 441524 296208 443362
rect 296824 441524 296852 445742
rect 297454 444952 297510 444961
rect 297454 444887 297510 444896
rect 297468 441524 297496 444887
rect 298112 441524 298140 445946
rect 299386 444816 299442 444825
rect 299386 444751 299442 444760
rect 298744 443216 298796 443222
rect 298744 443158 298796 443164
rect 298756 441524 298784 443158
rect 299400 441524 299428 444751
rect 300136 441524 300164 446014
rect 302700 445936 302752 445942
rect 302700 445878 302752 445884
rect 301412 443964 301464 443970
rect 301412 443906 301464 443912
rect 300768 442128 300820 442134
rect 300768 442070 300820 442076
rect 300780 441524 300808 442070
rect 301424 441524 301452 443906
rect 302056 442196 302108 442202
rect 302056 442138 302108 442144
rect 302068 441524 302096 442138
rect 302712 441524 302740 445878
rect 303540 443698 303568 476167
rect 306300 467158 306328 476167
rect 306288 467152 306340 467158
rect 306288 467094 306340 467100
rect 307300 465860 307352 465866
rect 307300 465802 307352 465808
rect 303988 444780 304040 444786
rect 303988 444722 304040 444728
rect 303528 443692 303580 443698
rect 303528 443634 303580 443640
rect 304000 441524 304028 444722
rect 306656 441856 306708 441862
rect 306010 441824 306066 441833
rect 306656 441798 306708 441804
rect 306010 441759 306066 441768
rect 306024 441524 306052 441759
rect 306668 441524 306696 441798
rect 307312 441524 307340 465802
rect 307944 447840 307996 447846
rect 307944 447782 307996 447788
rect 307956 441524 307984 447782
rect 308600 441524 308628 478314
rect 314476 478304 314528 478310
rect 314476 478246 314528 478252
rect 309046 476776 309102 476785
rect 309046 476711 309102 476720
rect 311256 476740 311308 476746
rect 309060 476338 309088 476711
rect 311256 476682 311308 476688
rect 309048 476332 309100 476338
rect 309048 476274 309100 476280
rect 309876 463140 309928 463146
rect 309876 463082 309928 463088
rect 309232 460352 309284 460358
rect 309232 460294 309284 460300
rect 309244 441524 309272 460294
rect 309888 441524 309916 463082
rect 310520 453620 310572 453626
rect 310520 453562 310572 453568
rect 310532 441524 310560 453562
rect 311268 441524 311296 476682
rect 311806 476368 311862 476377
rect 311806 476303 311862 476312
rect 311820 476270 311848 476303
rect 311808 476264 311860 476270
rect 311808 476206 311860 476212
rect 313832 476128 313884 476134
rect 313832 476070 313884 476076
rect 313188 460420 313240 460426
rect 313188 460362 313240 460368
rect 311900 454844 311952 454850
rect 311900 454786 311952 454792
rect 311912 441524 311940 454786
rect 312544 449744 312596 449750
rect 312544 449686 312596 449692
rect 312556 441524 312584 449686
rect 313200 441524 313228 460362
rect 313844 441524 313872 476070
rect 314488 441524 314516 478246
rect 321466 477048 321522 477057
rect 321466 476983 321522 476992
rect 316408 476808 316460 476814
rect 314566 476776 314622 476785
rect 316408 476750 316460 476756
rect 314566 476711 314622 476720
rect 314580 476134 314608 476711
rect 315946 476232 316002 476241
rect 315946 476167 315948 476176
rect 316000 476167 316002 476176
rect 315948 476138 316000 476144
rect 314568 476128 314620 476134
rect 314568 476070 314620 476076
rect 315764 470076 315816 470082
rect 315764 470018 315816 470024
rect 315120 449676 315172 449682
rect 315120 449618 315172 449624
rect 315132 441524 315160 449618
rect 315776 441524 315804 470018
rect 316420 441524 316448 476750
rect 319076 476672 319128 476678
rect 319076 476614 319128 476620
rect 318706 476504 318762 476513
rect 318432 476468 318484 476474
rect 318706 476439 318708 476448
rect 318432 476410 318484 476416
rect 318760 476439 318762 476448
rect 318708 476410 318760 476416
rect 317144 468648 317196 468654
rect 317144 468590 317196 468596
rect 317156 441524 317184 468590
rect 317788 464500 317840 464506
rect 317788 464442 317840 464448
rect 317800 441524 317828 464442
rect 318444 441524 318472 476410
rect 319088 441524 319116 476614
rect 321480 474026 321508 476983
rect 330208 476604 330260 476610
rect 330208 476546 330260 476552
rect 326896 476536 326948 476542
rect 324226 476504 324282 476513
rect 326896 476478 326948 476484
rect 326986 476504 327042 476513
rect 324226 476439 324282 476448
rect 323032 476400 323084 476406
rect 323032 476342 323084 476348
rect 321652 475448 321704 475454
rect 321652 475390 321704 475396
rect 321468 474020 321520 474026
rect 321468 473962 321520 473968
rect 319720 472796 319772 472802
rect 319720 472738 319772 472744
rect 319732 441524 319760 472738
rect 320364 468716 320416 468722
rect 320364 468658 320416 468664
rect 320376 441524 320404 468658
rect 321008 443896 321060 443902
rect 321008 443838 321060 443844
rect 321020 441524 321048 443838
rect 321664 441524 321692 475390
rect 322296 463072 322348 463078
rect 322296 463014 322348 463020
rect 322308 441524 322336 463014
rect 323044 441524 323072 476342
rect 324240 475454 324268 476439
rect 324228 475448 324280 475454
rect 324228 475390 324280 475396
rect 323676 474156 323728 474162
rect 323676 474098 323728 474104
rect 323688 441524 323716 474098
rect 326252 467356 326304 467362
rect 326252 467298 326304 467304
rect 325608 467288 325660 467294
rect 325608 467230 325660 467236
rect 324320 457632 324372 457638
rect 324320 457574 324372 457580
rect 324332 441524 324360 457574
rect 324964 443828 325016 443834
rect 324964 443770 325016 443776
rect 324976 441524 325004 443770
rect 325620 441524 325648 467230
rect 326264 441524 326292 467298
rect 326908 441524 326936 476478
rect 326986 476439 327042 476448
rect 327000 476406 327028 476439
rect 326988 476400 327040 476406
rect 326988 476342 327040 476348
rect 329104 476332 329156 476338
rect 329104 476274 329156 476280
rect 327540 471368 327592 471374
rect 327540 471310 327592 471316
rect 327552 441524 327580 471310
rect 328276 447976 328328 447982
rect 328276 447918 328328 447924
rect 328288 441524 328316 447918
rect 329116 443766 329144 476274
rect 329564 474224 329616 474230
rect 329564 474166 329616 474172
rect 328920 443760 328972 443766
rect 328920 443702 328972 443708
rect 329104 443760 329156 443766
rect 329104 443702 329156 443708
rect 328932 441524 328960 443702
rect 329576 441524 329604 474166
rect 330220 441524 330248 476546
rect 336004 476468 336056 476474
rect 336004 476410 336056 476416
rect 331864 476264 331916 476270
rect 331864 476206 331916 476212
rect 331496 475516 331548 475522
rect 331496 475458 331548 475464
rect 330852 470008 330904 470014
rect 330852 469950 330904 469956
rect 330864 441524 330892 469950
rect 331508 441524 331536 475458
rect 331876 443970 331904 476206
rect 334624 476196 334676 476202
rect 334624 476138 334676 476144
rect 333244 476128 333296 476134
rect 333244 476070 333296 476076
rect 332140 457564 332192 457570
rect 332140 457506 332192 457512
rect 331864 443964 331916 443970
rect 331864 443906 331916 443912
rect 332152 441524 332180 457506
rect 332784 450560 332836 450566
rect 332784 450502 332836 450508
rect 332796 441524 332824 450502
rect 333256 443902 333284 476070
rect 334164 456204 334216 456210
rect 334164 456146 334216 456152
rect 333428 448044 333480 448050
rect 333428 447986 333480 447992
rect 333244 443896 333296 443902
rect 333244 443838 333296 443844
rect 333440 441524 333468 447986
rect 334176 441524 334204 456146
rect 334636 444038 334664 476138
rect 334808 458992 334860 458998
rect 334808 458934 334860 458940
rect 334624 444032 334676 444038
rect 334624 443974 334676 443980
rect 334820 441524 334848 458934
rect 335452 458924 335504 458930
rect 335452 458866 335504 458872
rect 335464 441524 335492 458866
rect 336016 444106 336044 476410
rect 338764 476400 338816 476406
rect 338764 476342 338816 476348
rect 338028 471300 338080 471306
rect 338028 471242 338080 471248
rect 336096 456136 336148 456142
rect 336096 456078 336148 456084
rect 336004 444100 336056 444106
rect 336004 444042 336056 444048
rect 336108 441524 336136 456078
rect 336740 451920 336792 451926
rect 336740 451862 336792 451868
rect 336752 441524 336780 451862
rect 337384 450696 337436 450702
rect 337384 450638 337436 450644
rect 337396 441524 337424 450638
rect 338040 441524 338068 471242
rect 338672 461780 338724 461786
rect 338672 461722 338724 461728
rect 338684 441524 338712 461722
rect 338776 443834 338804 476342
rect 352564 475448 352616 475454
rect 352564 475390 352616 475396
rect 339408 469872 339460 469878
rect 339408 469814 339460 469820
rect 338764 443828 338816 443834
rect 338764 443770 338816 443776
rect 339420 441524 339448 469814
rect 343272 468512 343324 468518
rect 343272 468454 343324 468460
rect 341984 463208 342036 463214
rect 341984 463150 342036 463156
rect 340696 461644 340748 461650
rect 340696 461586 340748 461592
rect 340052 449404 340104 449410
rect 340052 449346 340104 449352
rect 340064 441524 340092 449346
rect 340708 441524 340736 461586
rect 341340 449540 341392 449546
rect 341340 449482 341392 449488
rect 341352 441524 341380 449482
rect 341996 441524 342024 463150
rect 342628 449608 342680 449614
rect 342628 449550 342680 449556
rect 342640 441524 342668 449550
rect 343284 441524 343312 468454
rect 348516 467152 348568 467158
rect 348516 467094 348568 467100
rect 344560 465724 344612 465730
rect 344560 465666 344612 465672
rect 343916 449472 343968 449478
rect 343916 449414 343968 449420
rect 343928 441524 343956 449414
rect 344572 441524 344600 465666
rect 345940 453416 345992 453422
rect 345940 453358 345992 453364
rect 345296 449200 345348 449206
rect 345296 449142 345348 449148
rect 345308 441524 345336 449142
rect 345952 441524 345980 453358
rect 346584 449336 346636 449342
rect 346584 449278 346636 449284
rect 346596 441524 346624 449278
rect 347872 449268 347924 449274
rect 347872 449210 347924 449216
rect 347228 443692 347280 443698
rect 347228 443634 347280 443640
rect 347240 441524 347268 443634
rect 347884 441524 347912 449210
rect 348528 441524 348556 467094
rect 351828 464432 351880 464438
rect 351828 464374 351880 464380
rect 349160 453484 349212 453490
rect 349160 453426 349212 453432
rect 349172 441524 349200 453426
rect 350540 452124 350592 452130
rect 350540 452066 350592 452072
rect 349804 443760 349856 443766
rect 349804 443702 349856 443708
rect 349816 441524 349844 443702
rect 350552 441524 350580 452066
rect 351184 443964 351236 443970
rect 351184 443906 351236 443912
rect 351196 441524 351224 443906
rect 351840 441524 351868 464374
rect 352472 443896 352524 443902
rect 352472 443838 352524 443844
rect 352484 441524 352512 443838
rect 352576 443698 352604 475390
rect 356428 474020 356480 474026
rect 356428 473962 356480 473968
rect 354404 472660 354456 472666
rect 354404 472602 354456 472608
rect 353116 447908 353168 447914
rect 353116 447850 353168 447856
rect 352564 443692 352616 443698
rect 352564 443634 352616 443640
rect 353128 441524 353156 447850
rect 353760 444032 353812 444038
rect 353760 443974 353812 443980
rect 353772 441524 353800 443974
rect 354416 441524 354444 472602
rect 355692 465928 355744 465934
rect 355692 465870 355744 465876
rect 355048 444100 355100 444106
rect 355048 444042 355100 444048
rect 355060 441524 355088 444042
rect 355704 441524 355732 465870
rect 356440 441524 356468 473962
rect 357072 460216 357124 460222
rect 357072 460158 357124 460164
rect 357084 441524 357112 460158
rect 358096 450634 358124 510614
rect 358832 478446 358860 700334
rect 359464 700324 359516 700330
rect 359464 700266 359516 700272
rect 358820 478440 358872 478446
rect 358820 478382 358872 478388
rect 359476 460290 359504 700266
rect 363604 616888 363656 616894
rect 363604 616830 363656 616836
rect 360844 563100 360896 563106
rect 360844 563042 360896 563048
rect 359464 460284 359516 460290
rect 359464 460226 359516 460232
rect 358360 454708 358412 454714
rect 358360 454650 358412 454656
rect 358084 450628 358136 450634
rect 358084 450570 358136 450576
rect 357716 443692 357768 443698
rect 357716 443634 357768 443640
rect 357728 441524 357756 443634
rect 358372 441524 358400 454650
rect 360856 451994 360884 563042
rect 363616 453354 363644 616830
rect 364352 461718 364380 702406
rect 397472 699718 397500 703520
rect 396724 699712 396776 699718
rect 396724 699654 396776 699660
rect 397460 699712 397512 699718
rect 397460 699654 397512 699660
rect 391204 696992 391256 696998
rect 391204 696934 391256 696940
rect 378784 683188 378836 683194
rect 378784 683130 378836 683136
rect 377404 670744 377456 670750
rect 377404 670686 377456 670692
rect 373264 643136 373316 643142
rect 373264 643078 373316 643084
rect 369124 536852 369176 536858
rect 369124 536794 369176 536800
rect 367744 484424 367796 484430
rect 367744 484366 367796 484372
rect 367756 472734 367784 484366
rect 369136 474094 369164 536794
rect 371884 524476 371936 524482
rect 371884 524418 371936 524424
rect 371896 475386 371924 524418
rect 371884 475380 371936 475386
rect 371884 475322 371936 475328
rect 369124 474088 369176 474094
rect 369124 474030 369176 474036
rect 367744 472728 367796 472734
rect 367744 472670 367796 472676
rect 373276 465798 373304 643078
rect 374644 590708 374696 590714
rect 374644 590650 374696 590656
rect 374656 478242 374684 590650
rect 374644 478236 374696 478242
rect 374644 478178 374696 478184
rect 373264 465792 373316 465798
rect 373264 465734 373316 465740
rect 364340 461712 364392 461718
rect 364340 461654 364392 461660
rect 377416 454782 377444 670686
rect 378796 469946 378824 683130
rect 378784 469940 378836 469946
rect 378784 469882 378836 469888
rect 391216 463010 391244 696934
rect 396736 464370 396764 699654
rect 396724 464364 396776 464370
rect 396724 464306 396776 464312
rect 391204 463004 391256 463010
rect 391204 462946 391256 462952
rect 377404 454776 377456 454782
rect 377404 454718 377456 454724
rect 363604 453348 363656 453354
rect 363604 453290 363656 453296
rect 360844 451988 360896 451994
rect 360844 451930 360896 451936
rect 412652 446758 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 429856 700330 429884 703520
rect 429844 700324 429896 700330
rect 429844 700266 429896 700272
rect 442264 700324 442316 700330
rect 442264 700266 442316 700272
rect 442276 456074 442304 700266
rect 462332 468586 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 462320 468580 462372 468586
rect 462320 468522 462372 468528
rect 442264 456068 442316 456074
rect 442264 456010 442316 456016
rect 412640 446752 412692 446758
rect 412640 446694 412692 446700
rect 477512 446690 477540 702406
rect 494072 458862 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 527192 467226 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 527180 467220 527232 467226
rect 527180 467162 527232 467168
rect 494060 458856 494112 458862
rect 494060 458798 494112 458804
rect 477500 446684 477552 446690
rect 477500 446626 477552 446632
rect 542372 446622 542400 702406
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580262 630864 580318 630873
rect 580262 630799 580318 630808
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580184 590714 580212 590951
rect 580172 590708 580224 590714
rect 580172 590650 580224 590656
rect 579894 564360 579950 564369
rect 579894 564295 579950 564304
rect 579908 563106 579936 564295
rect 579896 563100 579948 563106
rect 579896 563042 579948 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 580184 470626 580212 471407
rect 580172 470620 580224 470626
rect 580172 470562 580224 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 542360 446616 542412 446622
rect 542360 446558 542412 446564
rect 580276 446486 580304 630799
rect 580354 577688 580410 577697
rect 580354 577623 580410 577632
rect 580264 446480 580316 446486
rect 580264 446422 580316 446428
rect 580368 446418 580396 577623
rect 580356 446412 580408 446418
rect 580356 446354 580408 446360
rect 373264 445868 373316 445874
rect 373264 445810 373316 445816
rect 362224 444168 362276 444174
rect 362224 444110 362276 444116
rect 359004 443828 359056 443834
rect 359004 443770 359056 443776
rect 359016 441524 359044 443770
rect 359648 443216 359700 443222
rect 359648 443158 359700 443164
rect 359660 441524 359688 443158
rect 360292 443080 360344 443086
rect 360292 443022 360344 443028
rect 360304 441524 360332 443022
rect 360936 443012 360988 443018
rect 360936 442954 360988 442960
rect 360948 441524 360976 442954
rect 290004 441448 290056 441454
rect 290004 441390 290056 441396
rect 294604 441448 294656 441454
rect 294604 441390 294656 441396
rect 289818 441280 289874 441289
rect 289818 441215 289874 441224
rect 289832 441046 289860 441215
rect 290016 441046 290044 441390
rect 293592 441312 293644 441318
rect 293592 441254 293644 441260
rect 293774 441280 293830 441289
rect 293408 441244 293460 441250
rect 293408 441186 293460 441192
rect 290740 441176 290792 441182
rect 290738 441144 290740 441153
rect 290792 441144 290794 441153
rect 290738 441079 290794 441088
rect 293420 441046 293448 441186
rect 293604 441046 293632 441254
rect 294616 441250 294644 441390
rect 293774 441215 293830 441224
rect 294604 441244 294656 441250
rect 293682 441144 293738 441153
rect 293682 441079 293738 441088
rect 293696 441046 293724 441079
rect 293788 441046 293816 441215
rect 294604 441186 294656 441192
rect 240784 441040 240836 441046
rect 240534 440988 240784 440994
rect 247960 441040 248012 441046
rect 240534 440982 240836 440988
rect 247710 440988 247960 440994
rect 252008 441040 252060 441046
rect 247710 440982 248012 440988
rect 251666 440988 252008 440994
rect 251666 440982 252060 440988
rect 276112 441040 276164 441046
rect 276112 440982 276164 440988
rect 277400 441040 277452 441046
rect 277400 440982 277452 440988
rect 289820 441040 289872 441046
rect 289820 440982 289872 440988
rect 290004 441040 290056 441046
rect 290004 440982 290056 440988
rect 293408 441040 293460 441046
rect 293408 440982 293460 440988
rect 293592 441040 293644 441046
rect 293592 440982 293644 440988
rect 293684 441040 293736 441046
rect 293684 440982 293736 440988
rect 293776 441040 293828 441046
rect 293776 440982 293828 440988
rect 303068 441040 303120 441046
rect 304356 441040 304408 441046
rect 303120 440988 303370 440994
rect 303068 440982 303370 440988
rect 304998 441008 305054 441017
rect 304408 440988 304658 440994
rect 304356 440982 304658 440988
rect 240534 440966 240824 440982
rect 247710 440966 248000 440982
rect 251666 440966 252048 440982
rect 303080 440966 303370 440982
rect 304368 440966 304658 440982
rect 305054 440966 305302 440994
rect 304998 440943 305054 440952
rect 231216 411256 231268 411262
rect 231216 411198 231268 411204
rect 231124 398812 231176 398818
rect 231124 398754 231176 398760
rect 229744 377460 229796 377466
rect 229744 377402 229796 377408
rect 228364 374808 228416 374814
rect 228364 374750 228416 374756
rect 227076 374536 227128 374542
rect 227076 374478 227128 374484
rect 226984 372904 227036 372910
rect 226984 372846 227036 372852
rect 225696 336796 225748 336802
rect 225696 336738 225748 336744
rect 225708 310010 225736 336738
rect 225788 334008 225840 334014
rect 225788 333950 225840 333956
rect 225800 310593 225828 333950
rect 225786 310584 225842 310593
rect 225786 310519 225842 310528
rect 225696 310004 225748 310010
rect 225696 309946 225748 309952
rect 226996 308854 227024 372846
rect 227088 310554 227116 374478
rect 227076 310548 227128 310554
rect 227076 310490 227128 310496
rect 226984 308848 227036 308854
rect 226984 308790 227036 308796
rect 228376 307766 228404 374750
rect 229836 374740 229888 374746
rect 229836 374682 229888 374688
rect 228548 374400 228600 374406
rect 228548 374342 228600 374348
rect 228456 372768 228508 372774
rect 228456 372710 228508 372716
rect 228468 308786 228496 372710
rect 228560 309641 228588 374342
rect 229744 374196 229796 374202
rect 229744 374138 229796 374144
rect 228640 371612 228692 371618
rect 228640 371554 228692 371560
rect 228546 309632 228602 309641
rect 228546 309567 228602 309576
rect 228456 308780 228508 308786
rect 228456 308722 228508 308728
rect 228652 308689 228680 371554
rect 228732 357468 228784 357474
rect 228732 357410 228784 357416
rect 228744 309602 228772 357410
rect 228732 309596 228784 309602
rect 228732 309538 228784 309544
rect 228638 308680 228694 308689
rect 228638 308615 228694 308624
rect 228364 307760 228416 307766
rect 228364 307702 228416 307708
rect 229756 307562 229784 374138
rect 229744 307556 229796 307562
rect 229744 307498 229796 307504
rect 229848 307358 229876 374682
rect 231216 374264 231268 374270
rect 231216 374206 231268 374212
rect 231124 372836 231176 372842
rect 231124 372778 231176 372784
rect 229928 372700 229980 372706
rect 229928 372642 229980 372648
rect 229940 309058 229968 372642
rect 230020 371544 230072 371550
rect 230020 371486 230072 371492
rect 230032 309126 230060 371486
rect 230112 362976 230164 362982
rect 230112 362918 230164 362924
rect 230124 310350 230152 362918
rect 230204 331288 230256 331294
rect 230204 331230 230256 331236
rect 230112 310344 230164 310350
rect 230112 310286 230164 310292
rect 230216 309806 230244 331230
rect 231032 320204 231084 320210
rect 231032 320146 231084 320152
rect 230388 314696 230440 314702
rect 230388 314638 230440 314644
rect 230400 310758 230428 314638
rect 230848 311432 230900 311438
rect 230848 311374 230900 311380
rect 230388 310752 230440 310758
rect 230388 310694 230440 310700
rect 230756 310616 230808 310622
rect 230756 310558 230808 310564
rect 230204 309800 230256 309806
rect 230204 309742 230256 309748
rect 230020 309120 230072 309126
rect 230020 309062 230072 309068
rect 229928 309052 229980 309058
rect 229928 308994 229980 309000
rect 230768 308922 230796 310558
rect 230860 310146 230888 311374
rect 230940 311228 230992 311234
rect 230940 311170 230992 311176
rect 230952 310282 230980 311170
rect 230940 310276 230992 310282
rect 230940 310218 230992 310224
rect 230848 310140 230900 310146
rect 230848 310082 230900 310088
rect 231044 309330 231072 320146
rect 231032 309324 231084 309330
rect 231032 309266 231084 309272
rect 230756 308916 230808 308922
rect 230756 308858 230808 308864
rect 231136 308718 231164 372778
rect 231228 309913 231256 374206
rect 231308 371476 231360 371482
rect 231308 371418 231360 371424
rect 231214 309904 231270 309913
rect 231214 309839 231270 309848
rect 231320 309097 231348 371418
rect 231492 371408 231544 371414
rect 231492 371350 231544 371356
rect 231400 371340 231452 371346
rect 231400 371282 231452 371288
rect 231306 309088 231362 309097
rect 231306 309023 231362 309032
rect 231412 308990 231440 371282
rect 231400 308984 231452 308990
rect 231400 308926 231452 308932
rect 231504 308825 231532 371350
rect 231584 371272 231636 371278
rect 231584 371214 231636 371220
rect 231490 308816 231546 308825
rect 231490 308751 231546 308760
rect 231124 308712 231176 308718
rect 231124 308654 231176 308660
rect 231596 308242 231624 371214
rect 232228 368552 232280 368558
rect 232228 368494 232280 368500
rect 231676 365764 231728 365770
rect 231676 365706 231728 365712
rect 231688 309466 231716 365706
rect 232240 364334 232268 368494
rect 232240 364306 232360 364334
rect 232228 325712 232280 325718
rect 232228 325654 232280 325660
rect 231768 322992 231820 322998
rect 231768 322934 231820 322940
rect 231780 309942 231808 322934
rect 232240 321554 232268 325654
rect 231964 321526 232268 321554
rect 231860 317484 231912 317490
rect 231860 317426 231912 317432
rect 231872 310214 231900 317426
rect 231964 310418 231992 321526
rect 232044 311908 232096 311914
rect 232332 311894 232360 364306
rect 232044 311850 232096 311856
rect 232148 311866 232360 311894
rect 231952 310412 232004 310418
rect 231952 310354 232004 310360
rect 232056 310282 232084 311850
rect 231952 310276 232004 310282
rect 231952 310218 232004 310224
rect 232044 310276 232096 310282
rect 232044 310218 232096 310224
rect 231860 310208 231912 310214
rect 231860 310150 231912 310156
rect 231768 309936 231820 309942
rect 231768 309878 231820 309884
rect 231676 309460 231728 309466
rect 231676 309402 231728 309408
rect 231584 308236 231636 308242
rect 231584 308178 231636 308184
rect 231964 308038 231992 310218
rect 232044 310140 232096 310146
rect 232044 310082 232096 310088
rect 232056 308106 232084 310082
rect 232148 309534 232176 311866
rect 232228 311296 232280 311302
rect 232226 311264 232228 311273
rect 232280 311264 232282 311273
rect 232226 311199 232282 311208
rect 232228 311160 232280 311166
rect 232228 311102 232280 311108
rect 232240 310570 232268 311102
rect 233698 310584 233754 310593
rect 232240 310542 232530 310570
rect 233698 310519 233754 310528
rect 234066 310584 234122 310593
rect 255608 310554 255806 310570
rect 273732 310554 273930 310570
rect 234066 310519 234122 310528
rect 235448 310548 235500 310554
rect 232596 310480 232648 310486
rect 232410 310448 232466 310457
rect 232596 310422 232648 310428
rect 232410 310383 232466 310392
rect 232136 309528 232188 309534
rect 232136 309470 232188 309476
rect 232424 308514 232452 310383
rect 232608 310298 232636 310422
rect 232700 310298 232728 310420
rect 232884 310321 232912 310420
rect 233252 310350 233280 310420
rect 233240 310344 233292 310350
rect 232608 310270 232728 310298
rect 232870 310312 232926 310321
rect 233240 310286 233292 310292
rect 232870 310247 232926 310256
rect 233620 309126 233648 310420
rect 233712 310298 233740 310519
rect 233804 310298 233832 310420
rect 233712 310270 233832 310298
rect 233608 309120 233660 309126
rect 233608 309062 233660 309068
rect 232412 308508 232464 308514
rect 232412 308450 232464 308456
rect 232044 308100 232096 308106
rect 232044 308042 232096 308048
rect 231952 308032 232004 308038
rect 231952 307974 232004 307980
rect 229836 307352 229888 307358
rect 229836 307294 229888 307300
rect 233988 302234 234016 310420
rect 234080 309126 234108 310519
rect 235448 310490 235500 310496
rect 255412 310548 255464 310554
rect 255412 310490 255464 310496
rect 255596 310548 255806 310554
rect 255648 310542 255806 310548
rect 273536 310548 273588 310554
rect 255596 310490 255648 310496
rect 273536 310490 273588 310496
rect 273720 310548 273930 310554
rect 273772 310542 273930 310548
rect 314870 310554 315068 310570
rect 314870 310548 315080 310554
rect 314870 310542 315028 310548
rect 273720 310490 273772 310496
rect 315028 310490 315080 310496
rect 315396 310548 315448 310554
rect 315396 310490 315448 310496
rect 234172 309262 234200 310420
rect 234160 309256 234212 309262
rect 234160 309198 234212 309204
rect 234068 309120 234120 309126
rect 234068 309062 234120 309068
rect 233344 302206 234016 302234
rect 233344 300014 233372 302206
rect 233332 300008 233384 300014
rect 233332 299950 233384 299956
rect 234356 299305 234384 310420
rect 234540 308961 234568 310420
rect 234526 308952 234582 308961
rect 234526 308887 234582 308896
rect 234342 299296 234398 299305
rect 234342 299231 234398 299240
rect 234724 298586 234752 310420
rect 234908 308394 234936 310420
rect 234816 308366 234936 308394
rect 235000 310406 235198 310434
rect 234712 298580 234764 298586
rect 234712 298522 234764 298528
rect 234816 296614 234844 308366
rect 235000 305454 235028 310406
rect 235368 309058 235396 310420
rect 235460 310298 235488 310490
rect 235552 310298 235580 310420
rect 235460 310270 235580 310298
rect 235736 309097 235764 310420
rect 235920 309194 235948 310420
rect 235908 309188 235960 309194
rect 235908 309130 235960 309136
rect 235722 309088 235778 309097
rect 235356 309052 235408 309058
rect 235722 309023 235778 309032
rect 235356 308994 235408 309000
rect 236104 308310 236132 310420
rect 236288 310282 236316 310420
rect 236276 310276 236328 310282
rect 236276 310218 236328 310224
rect 236184 308440 236236 308446
rect 236472 308394 236500 310420
rect 236184 308382 236236 308388
rect 236092 308304 236144 308310
rect 236092 308246 236144 308252
rect 236092 308168 236144 308174
rect 236092 308110 236144 308116
rect 236104 306374 236132 308110
rect 235920 306346 236132 306374
rect 234988 305448 235040 305454
rect 234988 305390 235040 305396
rect 235920 297158 235948 306346
rect 236196 300150 236224 308382
rect 236288 308366 236500 308394
rect 236288 301617 236316 308366
rect 236368 308304 236420 308310
rect 236368 308246 236420 308252
rect 236274 301608 236330 301617
rect 236274 301543 236330 301552
rect 236184 300144 236236 300150
rect 236184 300086 236236 300092
rect 236380 297838 236408 308246
rect 236656 308174 236684 310420
rect 236840 308446 236868 310420
rect 237024 308990 237052 310420
rect 237012 308984 237064 308990
rect 237012 308926 237064 308932
rect 237104 308984 237156 308990
rect 237104 308926 237156 308932
rect 237116 308718 237144 308926
rect 237104 308712 237156 308718
rect 237104 308654 237156 308660
rect 236828 308440 236880 308446
rect 236828 308382 236880 308388
rect 236644 308168 236696 308174
rect 236644 308110 236696 308116
rect 236368 297832 236420 297838
rect 236368 297774 236420 297780
rect 235908 297152 235960 297158
rect 235908 297094 235960 297100
rect 237208 296714 237236 310420
rect 237288 308712 237340 308718
rect 237288 308654 237340 308660
rect 237300 308514 237328 308654
rect 237288 308508 237340 308514
rect 237288 308450 237340 308456
rect 237392 308394 237420 310420
rect 237590 310406 237788 310434
rect 237472 310072 237524 310078
rect 237472 310014 237524 310020
rect 237484 309194 237512 310014
rect 237472 309188 237524 309194
rect 237472 309130 237524 309136
rect 237392 308366 237696 308394
rect 237564 308304 237616 308310
rect 237564 308246 237616 308252
rect 237576 299441 237604 308246
rect 237562 299432 237618 299441
rect 237562 299367 237618 299376
rect 237668 297974 237696 308366
rect 237760 300218 237788 310406
rect 237852 308310 237880 310420
rect 237932 308508 237984 308514
rect 237932 308450 237984 308456
rect 237840 308304 237892 308310
rect 237840 308246 237892 308252
rect 237944 308106 237972 308450
rect 237932 308100 237984 308106
rect 237932 308042 237984 308048
rect 237748 300212 237800 300218
rect 237748 300154 237800 300160
rect 238036 299266 238064 310420
rect 238220 308378 238248 310420
rect 238208 308372 238260 308378
rect 238208 308314 238260 308320
rect 238404 307154 238432 310420
rect 238588 309126 238616 310420
rect 238772 309126 238800 310420
rect 238956 310010 238984 310420
rect 238944 310004 238996 310010
rect 238944 309946 238996 309952
rect 238576 309120 238628 309126
rect 238576 309062 238628 309068
rect 238760 309120 238812 309126
rect 238760 309062 238812 309068
rect 238852 308440 238904 308446
rect 239140 308394 239168 310420
rect 239324 308446 239352 310420
rect 239508 309942 239536 310420
rect 239496 309936 239548 309942
rect 239496 309878 239548 309884
rect 238852 308382 238904 308388
rect 238392 307148 238444 307154
rect 238392 307090 238444 307096
rect 238024 299260 238076 299266
rect 238024 299202 238076 299208
rect 238864 298994 238892 308382
rect 238944 308372 238996 308378
rect 238944 308314 238996 308320
rect 239048 308366 239168 308394
rect 239312 308440 239364 308446
rect 239312 308382 239364 308388
rect 238956 300286 238984 308314
rect 238944 300280 238996 300286
rect 238944 300222 238996 300228
rect 238852 298988 238904 298994
rect 238852 298930 238904 298936
rect 237656 297968 237708 297974
rect 237656 297910 237708 297916
rect 239048 297906 239076 308366
rect 239692 307018 239720 310420
rect 239772 309052 239824 309058
rect 239772 308994 239824 309000
rect 239784 308650 239812 308994
rect 239772 308644 239824 308650
rect 239772 308586 239824 308592
rect 239876 308378 239904 310420
rect 239864 308372 239916 308378
rect 239864 308314 239916 308320
rect 239680 307012 239732 307018
rect 239680 306954 239732 306960
rect 240060 304638 240088 310420
rect 240336 309913 240364 310420
rect 240322 309904 240378 309913
rect 240322 309839 240378 309848
rect 240140 308508 240192 308514
rect 240140 308450 240192 308456
rect 240048 304632 240100 304638
rect 240048 304574 240100 304580
rect 240152 300354 240180 308450
rect 240232 308440 240284 308446
rect 240520 308394 240548 310420
rect 240704 308446 240732 310420
rect 240232 308382 240284 308388
rect 240140 300348 240192 300354
rect 240140 300290 240192 300296
rect 240244 299334 240272 308382
rect 240324 308372 240376 308378
rect 240324 308314 240376 308320
rect 240428 308366 240548 308394
rect 240692 308440 240744 308446
rect 240692 308382 240744 308388
rect 240888 308378 240916 310420
rect 241072 308514 241100 310420
rect 241256 310049 241284 310420
rect 241242 310040 241298 310049
rect 241242 309975 241298 309984
rect 241060 308508 241112 308514
rect 241060 308450 241112 308456
rect 240876 308372 240928 308378
rect 240336 300422 240364 308314
rect 240428 302190 240456 308366
rect 240876 308314 240928 308320
rect 241440 306374 241468 310420
rect 241624 308718 241652 310420
rect 241808 310298 241836 310420
rect 241716 310270 241836 310298
rect 241716 309806 241744 310270
rect 241796 310208 241848 310214
rect 241796 310150 241848 310156
rect 241704 309800 241756 309806
rect 241704 309742 241756 309748
rect 241808 309398 241836 310150
rect 241796 309392 241848 309398
rect 241796 309334 241848 309340
rect 241612 308712 241664 308718
rect 241612 308654 241664 308660
rect 241992 308582 242020 310420
rect 242176 308786 242204 310420
rect 242164 308780 242216 308786
rect 242164 308722 242216 308728
rect 242360 308650 242388 310420
rect 242348 308644 242400 308650
rect 242348 308586 242400 308592
rect 241980 308576 242032 308582
rect 241980 308518 242032 308524
rect 242544 307426 242572 310420
rect 242532 307420 242584 307426
rect 242532 307362 242584 307368
rect 240520 306346 241468 306374
rect 240416 302184 240468 302190
rect 240416 302126 240468 302132
rect 240324 300416 240376 300422
rect 240324 300358 240376 300364
rect 240232 299328 240284 299334
rect 240232 299270 240284 299276
rect 239036 297900 239088 297906
rect 239036 297842 239088 297848
rect 236472 296686 237236 296714
rect 234804 296608 234856 296614
rect 234804 296550 234856 296556
rect 236472 296546 236500 296686
rect 240520 296682 240548 306346
rect 242728 300490 242756 310420
rect 243004 309602 243032 310420
rect 242992 309596 243044 309602
rect 242992 309538 243044 309544
rect 242808 308576 242860 308582
rect 242808 308518 242860 308524
rect 242820 300626 242848 308518
rect 242992 308440 243044 308446
rect 242992 308382 243044 308388
rect 243188 308394 243216 310420
rect 243372 308854 243400 310420
rect 243360 308848 243412 308854
rect 243360 308790 243412 308796
rect 243556 308446 243584 310420
rect 243544 308440 243596 308446
rect 242808 300620 242860 300626
rect 242808 300562 242860 300568
rect 242716 300484 242768 300490
rect 242716 300426 242768 300432
rect 243004 299402 243032 308382
rect 243188 308366 243308 308394
rect 243544 308382 243596 308388
rect 243176 308304 243228 308310
rect 243176 308246 243228 308252
rect 243084 307148 243136 307154
rect 243084 307090 243136 307096
rect 243096 300558 243124 307090
rect 243084 300552 243136 300558
rect 243084 300494 243136 300500
rect 242992 299396 243044 299402
rect 242992 299338 243044 299344
rect 243188 298790 243216 308246
rect 243280 306338 243308 308366
rect 243740 307290 243768 310420
rect 243728 307284 243780 307290
rect 243728 307226 243780 307232
rect 243924 307154 243952 310420
rect 244108 308310 244136 310420
rect 244096 308304 244148 308310
rect 244096 308246 244148 308252
rect 244292 307630 244320 310420
rect 244476 310350 244504 310420
rect 244464 310344 244516 310350
rect 244464 310286 244516 310292
rect 244660 309369 244688 310420
rect 244646 309360 244702 309369
rect 244646 309295 244702 309304
rect 244280 307624 244332 307630
rect 244280 307566 244332 307572
rect 244844 307494 244872 310420
rect 244832 307488 244884 307494
rect 244832 307430 244884 307436
rect 243912 307148 243964 307154
rect 243912 307090 243964 307096
rect 243268 306332 243320 306338
rect 243268 306274 243320 306280
rect 245028 302234 245056 310420
rect 245212 304978 245240 310420
rect 245200 304972 245252 304978
rect 245200 304914 245252 304920
rect 245488 304570 245516 310420
rect 245476 304564 245528 304570
rect 245476 304506 245528 304512
rect 244476 302206 245056 302234
rect 244476 299198 244504 302206
rect 245672 300801 245700 310420
rect 245856 308038 245884 310420
rect 245844 308032 245896 308038
rect 245844 307974 245896 307980
rect 246040 303482 246068 310420
rect 246028 303476 246080 303482
rect 246028 303418 246080 303424
rect 245658 300792 245714 300801
rect 245658 300727 245714 300736
rect 246224 300694 246252 310420
rect 246304 308712 246356 308718
rect 246304 308654 246356 308660
rect 246212 300688 246264 300694
rect 246212 300630 246264 300636
rect 244464 299192 244516 299198
rect 244464 299134 244516 299140
rect 243176 298784 243228 298790
rect 243176 298726 243228 298732
rect 240508 296676 240560 296682
rect 240508 296618 240560 296624
rect 236460 296540 236512 296546
rect 236460 296482 236512 296488
rect 225604 267708 225656 267714
rect 225604 267650 225656 267656
rect 246316 260166 246344 308654
rect 246408 308378 246436 310420
rect 246396 308372 246448 308378
rect 246396 308314 246448 308320
rect 246592 307766 246620 310420
rect 246776 309058 246804 310420
rect 246764 309052 246816 309058
rect 246764 308994 246816 309000
rect 246580 307760 246632 307766
rect 246580 307702 246632 307708
rect 246960 307698 246988 310420
rect 247144 308990 247172 310420
rect 247328 309777 247356 310420
rect 247314 309768 247370 309777
rect 247314 309703 247370 309712
rect 247512 309466 247540 310420
rect 247500 309460 247552 309466
rect 247500 309402 247552 309408
rect 247132 308984 247184 308990
rect 247132 308926 247184 308932
rect 246948 307692 247000 307698
rect 246948 307634 247000 307640
rect 247696 306354 247724 310420
rect 247776 307828 247828 307834
rect 247776 307770 247828 307776
rect 247132 306332 247184 306338
rect 247132 306274 247184 306280
rect 247328 306326 247724 306354
rect 247144 299130 247172 306274
rect 247328 299470 247356 306326
rect 247684 302660 247736 302666
rect 247684 302602 247736 302608
rect 247316 299464 247368 299470
rect 247316 299406 247368 299412
rect 247132 299124 247184 299130
rect 247132 299066 247184 299072
rect 247696 265674 247724 302602
rect 247788 298654 247816 307770
rect 247880 306338 247908 310420
rect 248156 309641 248184 310420
rect 248142 309632 248198 309641
rect 248142 309567 248198 309576
rect 248340 308825 248368 310420
rect 248326 308816 248382 308825
rect 247960 308780 248012 308786
rect 248326 308751 248382 308760
rect 247960 308722 248012 308728
rect 247868 306332 247920 306338
rect 247868 306274 247920 306280
rect 247972 302666 248000 308722
rect 248524 307834 248552 310420
rect 248512 307828 248564 307834
rect 248512 307770 248564 307776
rect 248512 306400 248564 306406
rect 248512 306342 248564 306348
rect 247960 302660 248012 302666
rect 247960 302602 248012 302608
rect 248524 298858 248552 306342
rect 248604 306332 248656 306338
rect 248604 306274 248656 306280
rect 248616 301209 248644 306274
rect 248602 301200 248658 301209
rect 248602 301135 248658 301144
rect 248512 298852 248564 298858
rect 248512 298794 248564 298800
rect 247776 298648 247828 298654
rect 247776 298590 247828 298596
rect 248708 296478 248736 310420
rect 248892 304502 248920 310420
rect 249076 309534 249104 310420
rect 249064 309528 249116 309534
rect 249064 309470 249116 309476
rect 249260 306406 249288 310420
rect 249248 306400 249300 306406
rect 249248 306342 249300 306348
rect 249444 306338 249472 310420
rect 249628 309398 249656 310420
rect 249616 309392 249668 309398
rect 249616 309334 249668 309340
rect 249812 309330 249840 310420
rect 249800 309324 249852 309330
rect 249800 309266 249852 309272
rect 249996 307222 250024 310420
rect 249984 307216 250036 307222
rect 249984 307158 250036 307164
rect 250180 306354 250208 310420
rect 250364 308281 250392 310420
rect 250456 310406 250654 310434
rect 250350 308272 250406 308281
rect 250350 308207 250406 308216
rect 250456 308122 250484 310406
rect 250272 308094 250484 308122
rect 250272 307562 250300 308094
rect 250824 307986 250852 310420
rect 250904 308644 250956 308650
rect 250904 308586 250956 308592
rect 250364 307958 250852 307986
rect 250260 307556 250312 307562
rect 250260 307498 250312 307504
rect 249432 306332 249484 306338
rect 249432 306274 249484 306280
rect 249904 306326 250208 306354
rect 248880 304496 248932 304502
rect 248880 304438 248932 304444
rect 249904 300830 249932 306326
rect 250364 302234 250392 307958
rect 250916 307902 250944 308586
rect 251008 308553 251036 310420
rect 251088 308848 251140 308854
rect 251088 308790 251140 308796
rect 250994 308544 251050 308553
rect 250994 308479 251050 308488
rect 251100 307970 251128 308790
rect 251088 307964 251140 307970
rect 251088 307906 251140 307912
rect 250444 307896 250496 307902
rect 250444 307838 250496 307844
rect 250536 307896 250588 307902
rect 250536 307838 250588 307844
rect 250904 307896 250956 307902
rect 250904 307838 250956 307844
rect 249996 302206 250392 302234
rect 249892 300824 249944 300830
rect 249892 300766 249944 300772
rect 249996 299062 250024 302206
rect 249984 299056 250036 299062
rect 249984 298998 250036 299004
rect 248696 296472 248748 296478
rect 248696 296414 248748 296420
rect 247684 265668 247736 265674
rect 247684 265610 247736 265616
rect 246304 260160 246356 260166
rect 246304 260102 246356 260108
rect 250456 244934 250484 307838
rect 250548 275330 250576 307838
rect 250628 307828 250680 307834
rect 250628 307770 250680 307776
rect 250640 298926 250668 307770
rect 251192 306354 251220 310420
rect 251376 307834 251404 310420
rect 251364 307828 251416 307834
rect 251364 307770 251416 307776
rect 251192 306326 251496 306354
rect 251364 305448 251416 305454
rect 251364 305390 251416 305396
rect 251376 300762 251404 305390
rect 251364 300756 251416 300762
rect 251364 300698 251416 300704
rect 250628 298920 250680 298926
rect 250628 298862 250680 298868
rect 251468 297090 251496 306326
rect 251560 303006 251588 310420
rect 251744 309233 251772 310420
rect 251730 309224 251786 309233
rect 251730 309159 251786 309168
rect 251928 306490 251956 310420
rect 252008 307896 252060 307902
rect 252008 307838 252060 307844
rect 251652 306462 251956 306490
rect 251652 305454 251680 306462
rect 251732 306332 251784 306338
rect 251732 306274 251784 306280
rect 251640 305448 251692 305454
rect 251640 305390 251692 305396
rect 251548 303000 251600 303006
rect 251548 302942 251600 302948
rect 251744 298722 251772 306274
rect 252020 304994 252048 307838
rect 252112 306338 252140 310420
rect 252192 307964 252244 307970
rect 252192 307906 252244 307912
rect 252100 306332 252152 306338
rect 252100 306274 252152 306280
rect 251836 304966 252048 304994
rect 251732 298716 251784 298722
rect 251732 298658 251784 298664
rect 251456 297084 251508 297090
rect 251456 297026 251508 297032
rect 250536 275324 250588 275330
rect 250536 275266 250588 275272
rect 251836 257582 251864 304966
rect 252204 302234 252232 307906
rect 252296 307358 252324 310420
rect 252480 308582 252508 310420
rect 252664 308689 252692 310420
rect 252848 308922 252876 310420
rect 252836 308916 252888 308922
rect 252836 308858 252888 308864
rect 252650 308680 252706 308689
rect 252650 308615 252706 308624
rect 252468 308576 252520 308582
rect 252468 308518 252520 308524
rect 252284 307352 252336 307358
rect 252284 307294 252336 307300
rect 253032 307018 253060 310420
rect 253124 310406 253322 310434
rect 253020 307012 253072 307018
rect 253020 306954 253072 306960
rect 252836 306808 252888 306814
rect 252836 306750 252888 306756
rect 252744 306536 252796 306542
rect 252744 306478 252796 306484
rect 252652 306468 252704 306474
rect 252652 306410 252704 306416
rect 251928 302206 252232 302234
rect 251928 260438 251956 302206
rect 251916 260432 251968 260438
rect 251916 260374 251968 260380
rect 251824 257576 251876 257582
rect 251824 257518 251876 257524
rect 252664 247722 252692 306410
rect 252756 262886 252784 306478
rect 252848 284986 252876 306750
rect 253124 306542 253152 310406
rect 253204 308576 253256 308582
rect 253204 308518 253256 308524
rect 253112 306536 253164 306542
rect 253112 306478 253164 306484
rect 253112 306332 253164 306338
rect 253112 306274 253164 306280
rect 253124 306218 253152 306274
rect 252940 306190 253152 306218
rect 252940 286346 252968 306190
rect 253020 305448 253072 305454
rect 253020 305390 253072 305396
rect 252928 286340 252980 286346
rect 252928 286282 252980 286288
rect 252836 284980 252888 284986
rect 252836 284922 252888 284928
rect 252744 262880 252796 262886
rect 252744 262822 252796 262828
rect 252652 247716 252704 247722
rect 252652 247658 252704 247664
rect 253032 246362 253060 305390
rect 253216 247926 253244 308518
rect 253492 306474 253520 310420
rect 253480 306468 253532 306474
rect 253480 306410 253532 306416
rect 253676 306338 253704 310420
rect 253664 306332 253716 306338
rect 253664 306274 253716 306280
rect 253860 305454 253888 310420
rect 253940 306332 253992 306338
rect 253940 306274 253992 306280
rect 253952 305862 253980 306274
rect 254044 305862 254072 310420
rect 254228 306320 254256 310420
rect 254412 308786 254440 310420
rect 254400 308780 254452 308786
rect 254400 308722 254452 308728
rect 254596 306354 254624 310420
rect 254136 306292 254256 306320
rect 254320 306326 254624 306354
rect 253940 305856 253992 305862
rect 253940 305798 253992 305804
rect 254032 305856 254084 305862
rect 254032 305798 254084 305804
rect 253848 305448 253900 305454
rect 253848 305390 253900 305396
rect 254032 305448 254084 305454
rect 254032 305390 254084 305396
rect 254044 273970 254072 305390
rect 254136 289134 254164 306292
rect 254216 305856 254268 305862
rect 254216 305798 254268 305804
rect 254228 290494 254256 305798
rect 254320 293282 254348 306326
rect 254780 305454 254808 310420
rect 254768 305448 254820 305454
rect 254768 305390 254820 305396
rect 254964 302234 254992 310420
rect 255148 306338 255176 310420
rect 255332 306338 255360 310420
rect 255136 306332 255188 306338
rect 255136 306274 255188 306280
rect 255320 306332 255372 306338
rect 255320 306274 255372 306280
rect 254412 302206 254992 302234
rect 254308 293276 254360 293282
rect 254308 293218 254360 293224
rect 254216 290488 254268 290494
rect 254216 290430 254268 290436
rect 254124 289128 254176 289134
rect 254124 289070 254176 289076
rect 254032 273964 254084 273970
rect 254032 273906 254084 273912
rect 254412 261526 254440 302206
rect 254400 261520 254452 261526
rect 254400 261462 254452 261468
rect 255424 257446 255452 310490
rect 255530 310406 255728 310434
rect 255596 306332 255648 306338
rect 255596 306274 255648 306280
rect 255504 305380 255556 305386
rect 255504 305322 255556 305328
rect 255412 257440 255464 257446
rect 255412 257382 255464 257388
rect 255516 257378 255544 305322
rect 255608 283626 255636 306274
rect 255700 305862 255728 310406
rect 255976 308718 256004 310420
rect 255964 308712 256016 308718
rect 255964 308654 256016 308660
rect 256160 306354 256188 310420
rect 256240 307964 256292 307970
rect 256240 307906 256292 307912
rect 255792 306326 256188 306354
rect 255688 305856 255740 305862
rect 255688 305798 255740 305804
rect 255688 305448 255740 305454
rect 255688 305390 255740 305396
rect 255700 287706 255728 305390
rect 255792 300121 255820 306326
rect 255872 305856 255924 305862
rect 255872 305798 255924 305804
rect 255778 300112 255834 300121
rect 255778 300047 255834 300056
rect 255688 287700 255740 287706
rect 255688 287642 255740 287648
rect 255596 283620 255648 283626
rect 255596 283562 255648 283568
rect 255504 257372 255556 257378
rect 255504 257314 255556 257320
rect 255884 256018 255912 305798
rect 256252 296714 256280 307906
rect 256344 305454 256372 310420
rect 256332 305448 256384 305454
rect 256332 305390 256384 305396
rect 256528 305386 256556 310420
rect 256608 306536 256660 306542
rect 256608 306478 256660 306484
rect 256516 305380 256568 305386
rect 256516 305322 256568 305328
rect 256620 304230 256648 306478
rect 256712 304366 256740 310420
rect 256792 306468 256844 306474
rect 256792 306410 256844 306416
rect 256700 304360 256752 304366
rect 256700 304302 256752 304308
rect 256608 304224 256660 304230
rect 256608 304166 256660 304172
rect 256804 302234 256832 306410
rect 256896 304366 256924 310420
rect 257080 306898 257108 310420
rect 256988 306870 257108 306898
rect 256988 306626 257016 306870
rect 256988 306598 257200 306626
rect 257172 305862 257200 306598
rect 257264 306542 257292 310420
rect 257252 306536 257304 306542
rect 257252 306478 257304 306484
rect 257448 306474 257476 310420
rect 257436 306468 257488 306474
rect 257436 306410 257488 306416
rect 257632 306354 257660 310420
rect 257816 308854 257844 310420
rect 257804 308848 257856 308854
rect 257804 308790 257856 308796
rect 257712 307828 257764 307834
rect 257712 307770 257764 307776
rect 257264 306326 257660 306354
rect 257160 305856 257212 305862
rect 257160 305798 257212 305804
rect 257160 305448 257212 305454
rect 257160 305390 257212 305396
rect 256884 304360 256936 304366
rect 256884 304302 256936 304308
rect 257068 304360 257120 304366
rect 257068 304302 257120 304308
rect 256976 304224 257028 304230
rect 256976 304166 257028 304172
rect 256804 302206 256924 302234
rect 255976 296686 256280 296714
rect 255872 256012 255924 256018
rect 255872 255954 255924 255960
rect 255976 250714 256004 296686
rect 256896 260302 256924 302206
rect 256988 276690 257016 304166
rect 257080 285054 257108 304302
rect 257068 285048 257120 285054
rect 257068 284990 257120 284996
rect 256976 276684 257028 276690
rect 256976 276626 257028 276632
rect 256884 260296 256936 260302
rect 256884 260238 256936 260244
rect 255964 250708 256016 250714
rect 255964 250650 256016 250656
rect 253204 247920 253256 247926
rect 253204 247862 253256 247868
rect 257172 247790 257200 305390
rect 257264 260234 257292 306326
rect 257724 306218 257752 307770
rect 257356 306190 257752 306218
rect 257356 279478 257384 306190
rect 257436 305856 257488 305862
rect 257436 305798 257488 305804
rect 257448 291854 257476 305798
rect 258000 305454 258028 310420
rect 258184 308938 258212 310420
rect 258092 308910 258212 308938
rect 258276 310406 258474 310434
rect 258092 305862 258120 308910
rect 258172 308780 258224 308786
rect 258172 308722 258224 308728
rect 258080 305856 258132 305862
rect 258080 305798 258132 305804
rect 257988 305448 258040 305454
rect 257988 305390 258040 305396
rect 257436 291848 257488 291854
rect 257436 291790 257488 291796
rect 257344 279472 257396 279478
rect 257344 279414 257396 279420
rect 258184 265742 258212 308722
rect 258276 278050 258304 310406
rect 258540 306332 258592 306338
rect 258540 306274 258592 306280
rect 258356 305856 258408 305862
rect 258356 305798 258408 305804
rect 258448 305856 258500 305862
rect 258448 305798 258500 305804
rect 258368 280838 258396 305798
rect 258460 286414 258488 305798
rect 258448 286408 258500 286414
rect 258448 286350 258500 286356
rect 258356 280832 258408 280838
rect 258356 280774 258408 280780
rect 258264 278044 258316 278050
rect 258264 277986 258316 277992
rect 258172 265736 258224 265742
rect 258172 265678 258224 265684
rect 257252 260228 257304 260234
rect 257252 260170 257304 260176
rect 258552 247858 258580 306274
rect 258644 294642 258672 310420
rect 258828 308786 258856 310420
rect 258816 308780 258868 308786
rect 258816 308722 258868 308728
rect 258816 308576 258868 308582
rect 258816 308518 258868 308524
rect 258828 307902 258856 308518
rect 258816 307896 258868 307902
rect 258816 307838 258868 307844
rect 259012 307834 259040 310420
rect 259000 307828 259052 307834
rect 259000 307770 259052 307776
rect 259196 305862 259224 310420
rect 259380 306338 259408 310420
rect 259564 308854 259592 310420
rect 259552 308848 259604 308854
rect 259552 308790 259604 308796
rect 259748 306456 259776 310420
rect 259564 306428 259776 306456
rect 259368 306332 259420 306338
rect 259368 306274 259420 306280
rect 259184 305856 259236 305862
rect 259184 305798 259236 305804
rect 258632 294636 258684 294642
rect 258632 294578 258684 294584
rect 259564 251870 259592 306428
rect 259644 306332 259696 306338
rect 259932 306320 259960 310420
rect 259644 306274 259696 306280
rect 259748 306292 259960 306320
rect 259656 251938 259684 306274
rect 259748 282198 259776 306292
rect 260116 303113 260144 310420
rect 260102 303104 260158 303113
rect 260102 303039 260158 303048
rect 260300 302954 260328 310420
rect 259840 302926 260328 302954
rect 259840 286482 259868 302926
rect 260484 302234 260512 310420
rect 260564 308644 260616 308650
rect 260564 308586 260616 308592
rect 260024 302206 260512 302234
rect 259828 286476 259880 286482
rect 259828 286418 259880 286424
rect 259736 282192 259788 282198
rect 259736 282134 259788 282140
rect 259644 251932 259696 251938
rect 259644 251874 259696 251880
rect 259552 251864 259604 251870
rect 259552 251806 259604 251812
rect 258540 247852 258592 247858
rect 258540 247794 258592 247800
rect 257160 247784 257212 247790
rect 257160 247726 257212 247732
rect 260024 246430 260052 302206
rect 260576 296714 260604 308586
rect 260668 306338 260696 310420
rect 260852 310406 260958 310434
rect 260656 306332 260708 306338
rect 260656 306274 260708 306280
rect 260852 305454 260880 310406
rect 261128 306762 261156 310420
rect 260944 306734 261156 306762
rect 260840 305448 260892 305454
rect 260840 305390 260892 305396
rect 260840 305312 260892 305318
rect 260840 305254 260892 305260
rect 260116 296686 260604 296714
rect 260116 272678 260144 296686
rect 260852 293350 260880 305254
rect 260840 293344 260892 293350
rect 260840 293286 260892 293292
rect 260104 272672 260156 272678
rect 260104 272614 260156 272620
rect 260944 250510 260972 306734
rect 261312 306626 261340 310420
rect 261036 306598 261340 306626
rect 261036 262954 261064 306598
rect 261496 306490 261524 310420
rect 261220 306462 261524 306490
rect 261116 305380 261168 305386
rect 261116 305322 261168 305328
rect 261128 271182 261156 305322
rect 261220 272542 261248 306462
rect 261680 306354 261708 310420
rect 261760 307896 261812 307902
rect 261760 307838 261812 307844
rect 261404 306326 261708 306354
rect 261300 305448 261352 305454
rect 261300 305390 261352 305396
rect 261312 290562 261340 305390
rect 261300 290556 261352 290562
rect 261300 290498 261352 290504
rect 261208 272536 261260 272542
rect 261208 272478 261260 272484
rect 261116 271176 261168 271182
rect 261116 271118 261168 271124
rect 261024 262948 261076 262954
rect 261024 262890 261076 262896
rect 260932 250504 260984 250510
rect 260932 250446 260984 250452
rect 261404 249082 261432 306326
rect 261772 302234 261800 307838
rect 261864 305318 261892 310420
rect 262048 305386 262076 310420
rect 262036 305380 262088 305386
rect 262036 305322 262088 305328
rect 261852 305312 261904 305318
rect 261852 305254 261904 305260
rect 261496 302206 261800 302234
rect 262232 302234 262260 310420
rect 262416 307970 262444 310420
rect 262404 307964 262456 307970
rect 262404 307906 262456 307912
rect 262600 306898 262628 310420
rect 262324 306870 262628 306898
rect 262324 302326 262352 306870
rect 262404 306332 262456 306338
rect 262784 306320 262812 310420
rect 262404 306274 262456 306280
rect 262508 306292 262812 306320
rect 262312 302320 262364 302326
rect 262312 302262 262364 302268
rect 262232 302206 262352 302234
rect 261496 257514 261524 302206
rect 261484 257508 261536 257514
rect 261484 257450 261536 257456
rect 261392 249076 261444 249082
rect 261392 249018 261444 249024
rect 262324 246838 262352 302206
rect 262312 246832 262364 246838
rect 262312 246774 262364 246780
rect 262416 246498 262444 306274
rect 262508 249150 262536 306292
rect 262968 306218 262996 310420
rect 263152 306338 263180 310420
rect 263140 306332 263192 306338
rect 263140 306274 263192 306280
rect 262692 306190 262996 306218
rect 262588 305856 262640 305862
rect 262588 305798 262640 305804
rect 262600 250578 262628 305798
rect 262692 260370 262720 306190
rect 263336 305862 263364 310420
rect 263612 309134 263640 310420
rect 263520 309106 263640 309134
rect 263324 305856 263376 305862
rect 263324 305798 263376 305804
rect 263520 304366 263548 309106
rect 263796 305862 263824 310420
rect 263980 306354 264008 310420
rect 264164 306490 264192 310420
rect 263888 306326 264008 306354
rect 264072 306462 264192 306490
rect 263600 305856 263652 305862
rect 263600 305798 263652 305804
rect 263784 305856 263836 305862
rect 263784 305798 263836 305804
rect 263508 304360 263560 304366
rect 263508 304302 263560 304308
rect 262772 302252 262824 302258
rect 262772 302194 262824 302200
rect 262680 260364 262732 260370
rect 262680 260306 262732 260312
rect 262588 250572 262640 250578
rect 262588 250514 262640 250520
rect 262496 249144 262548 249150
rect 262496 249086 262548 249092
rect 262404 246492 262456 246498
rect 262404 246434 262456 246440
rect 260012 246424 260064 246430
rect 260012 246366 260064 246372
rect 253020 246356 253072 246362
rect 253020 246298 253072 246304
rect 262784 245002 262812 302194
rect 263612 291922 263640 305798
rect 263784 305448 263836 305454
rect 263784 305390 263836 305396
rect 263692 304360 263744 304366
rect 263692 304302 263744 304308
rect 263600 291916 263652 291922
rect 263600 291858 263652 291864
rect 263704 250646 263732 304302
rect 263796 261594 263824 305390
rect 263888 264246 263916 306326
rect 264072 306218 264100 306462
rect 264348 306354 264376 310420
rect 264428 307828 264480 307834
rect 264428 307770 264480 307776
rect 263980 306190 264100 306218
rect 264164 306326 264376 306354
rect 263980 267034 264008 306190
rect 264060 305856 264112 305862
rect 264060 305798 264112 305804
rect 264072 269822 264100 305798
rect 264164 279546 264192 306326
rect 264440 302234 264468 307770
rect 264532 305454 264560 310420
rect 264520 305448 264572 305454
rect 264520 305390 264572 305396
rect 264256 302206 264468 302234
rect 264152 279540 264204 279546
rect 264152 279482 264204 279488
rect 264060 269816 264112 269822
rect 264060 269758 264112 269764
rect 263968 267028 264020 267034
rect 263968 266970 264020 266976
rect 263876 264240 263928 264246
rect 263876 264182 263928 264188
rect 263784 261588 263836 261594
rect 263784 261530 263836 261536
rect 264256 254658 264284 302206
rect 264716 296714 264744 310420
rect 264900 305862 264928 310420
rect 264980 306400 265032 306406
rect 264980 306342 265032 306348
rect 264888 305856 264940 305862
rect 264888 305798 264940 305804
rect 264348 296686 264744 296714
rect 264244 254652 264296 254658
rect 264244 254594 264296 254600
rect 263692 250640 263744 250646
rect 263692 250582 263744 250588
rect 264348 249218 264376 296686
rect 264992 249286 265020 306342
rect 265084 305862 265112 310420
rect 265268 306354 265296 310420
rect 265176 306326 265296 306354
rect 265348 306332 265400 306338
rect 265072 305856 265124 305862
rect 265072 305798 265124 305804
rect 265072 305448 265124 305454
rect 265072 305390 265124 305396
rect 265084 253230 265112 305390
rect 265176 256086 265204 306326
rect 265348 306274 265400 306280
rect 265256 305856 265308 305862
rect 265256 305798 265308 305804
rect 265268 268394 265296 305798
rect 265360 272610 265388 306274
rect 265452 278118 265480 310420
rect 265636 305454 265664 310420
rect 265624 305448 265676 305454
rect 265624 305390 265676 305396
rect 265820 296714 265848 310420
rect 265912 310406 266110 310434
rect 265912 306406 265940 310406
rect 265900 306400 265952 306406
rect 265900 306342 265952 306348
rect 266280 306338 266308 310420
rect 266268 306332 266320 306338
rect 266268 306274 266320 306280
rect 265544 296686 265848 296714
rect 265544 285122 265572 296686
rect 265532 285116 265584 285122
rect 265532 285058 265584 285064
rect 265440 278112 265492 278118
rect 265440 278054 265492 278060
rect 265348 272604 265400 272610
rect 265348 272546 265400 272552
rect 265256 268388 265308 268394
rect 265256 268330 265308 268336
rect 265164 256080 265216 256086
rect 265164 256022 265216 256028
rect 266464 253298 266492 310420
rect 266648 306406 266676 310420
rect 266832 309134 266860 310420
rect 266740 309106 266860 309134
rect 266636 306400 266688 306406
rect 266636 306342 266688 306348
rect 266544 306332 266596 306338
rect 266544 306274 266596 306280
rect 266556 254726 266584 306274
rect 266740 305946 266768 309106
rect 267016 307834 267044 310420
rect 267096 308780 267148 308786
rect 267096 308722 267148 308728
rect 267004 307828 267056 307834
rect 267004 307770 267056 307776
rect 267004 306400 267056 306406
rect 267004 306342 267056 306348
rect 266648 305918 266768 305946
rect 266544 254720 266596 254726
rect 266544 254662 266596 254668
rect 266648 254590 266676 305918
rect 266728 305856 266780 305862
rect 267016 305844 267044 306342
rect 266728 305798 266780 305804
rect 266832 305816 267044 305844
rect 266740 256154 266768 305798
rect 266728 256148 266780 256154
rect 266728 256090 266780 256096
rect 266636 254584 266688 254590
rect 266636 254526 266688 254532
rect 266452 253292 266504 253298
rect 266452 253234 266504 253240
rect 265072 253224 265124 253230
rect 265072 253166 265124 253172
rect 264980 249280 265032 249286
rect 264980 249222 265032 249228
rect 264336 249212 264388 249218
rect 264336 249154 264388 249160
rect 266832 246566 266860 305816
rect 267108 302234 267136 308722
rect 267200 308718 267228 310420
rect 267188 308712 267240 308718
rect 267188 308654 267240 308660
rect 267384 306338 267412 310420
rect 267372 306332 267424 306338
rect 267372 306274 267424 306280
rect 267568 305862 267596 310420
rect 267752 306338 267780 310420
rect 267936 306746 267964 310420
rect 267924 306740 267976 306746
rect 267924 306682 267976 306688
rect 268120 306626 268148 310420
rect 267844 306598 268148 306626
rect 267740 306332 267792 306338
rect 267740 306274 267792 306280
rect 267556 305856 267608 305862
rect 267556 305798 267608 305804
rect 267016 302206 267136 302234
rect 267016 258874 267044 302206
rect 267004 258868 267056 258874
rect 267004 258810 267056 258816
rect 267844 254794 267872 306598
rect 267924 306468 267976 306474
rect 267924 306410 267976 306416
rect 267936 269890 267964 306410
rect 268304 306354 268332 310420
rect 268016 306332 268068 306338
rect 268016 306274 268068 306280
rect 268120 306326 268332 306354
rect 268028 274038 268056 306274
rect 268120 275398 268148 306326
rect 268488 302234 268516 310420
rect 268764 308650 268792 310420
rect 268752 308644 268804 308650
rect 268752 308586 268804 308592
rect 268212 302206 268516 302234
rect 268212 279614 268240 302206
rect 268948 296714 268976 310420
rect 269132 305862 269160 310420
rect 269212 306468 269264 306474
rect 269212 306410 269264 306416
rect 269120 305856 269172 305862
rect 269120 305798 269172 305804
rect 268304 296686 268976 296714
rect 268200 279608 268252 279614
rect 268200 279550 268252 279556
rect 268108 275392 268160 275398
rect 268108 275334 268160 275340
rect 268016 274032 268068 274038
rect 268016 273974 268068 273980
rect 267924 269884 267976 269890
rect 267924 269826 267976 269832
rect 267832 254788 267884 254794
rect 267832 254730 267884 254736
rect 266820 246560 266872 246566
rect 266820 246502 266872 246508
rect 268304 245070 268332 296686
rect 269224 246634 269252 306410
rect 269316 306354 269344 310420
rect 269500 306354 269528 310420
rect 269684 306474 269712 310420
rect 269868 307902 269896 310420
rect 269856 307896 269908 307902
rect 269856 307838 269908 307844
rect 269672 306468 269724 306474
rect 269672 306410 269724 306416
rect 269316 306326 269436 306354
rect 269500 306326 269804 306354
rect 269304 305380 269356 305386
rect 269304 305322 269356 305328
rect 269316 269958 269344 305322
rect 269408 271250 269436 306326
rect 269488 305856 269540 305862
rect 269488 305798 269540 305804
rect 269580 305856 269632 305862
rect 269580 305798 269632 305804
rect 269500 278186 269528 305798
rect 269592 280906 269620 305798
rect 269672 305448 269724 305454
rect 269672 305390 269724 305396
rect 269580 280900 269632 280906
rect 269580 280842 269632 280848
rect 269488 278180 269540 278186
rect 269488 278122 269540 278128
rect 269396 271244 269448 271250
rect 269396 271186 269448 271192
rect 269304 269952 269356 269958
rect 269304 269894 269356 269900
rect 269212 246628 269264 246634
rect 269212 246570 269264 246576
rect 269684 245138 269712 305390
rect 269776 289202 269804 306326
rect 270052 305862 270080 310420
rect 270040 305856 270092 305862
rect 270040 305798 270092 305804
rect 270236 305454 270264 310420
rect 270224 305448 270276 305454
rect 270224 305390 270276 305396
rect 270420 305386 270448 310420
rect 270604 305862 270632 310420
rect 270684 306468 270736 306474
rect 270684 306410 270736 306416
rect 270592 305856 270644 305862
rect 270592 305798 270644 305804
rect 270408 305380 270460 305386
rect 270408 305322 270460 305328
rect 270592 305380 270644 305386
rect 270592 305322 270644 305328
rect 269764 289196 269816 289202
rect 269764 289138 269816 289144
rect 270604 253434 270632 305322
rect 270696 274106 270724 306410
rect 270788 306354 270816 310420
rect 270972 306474 271000 310420
rect 271064 310406 271262 310434
rect 270960 306468 271012 306474
rect 270960 306410 271012 306416
rect 271064 306354 271092 310406
rect 271144 308508 271196 308514
rect 271144 308450 271196 308456
rect 270788 306326 270908 306354
rect 270776 305448 270828 305454
rect 270776 305390 270828 305396
rect 270788 275466 270816 305390
rect 270880 276758 270908 306326
rect 270972 306326 271092 306354
rect 270972 282266 271000 306326
rect 271052 305856 271104 305862
rect 271052 305798 271104 305804
rect 270960 282260 271012 282266
rect 270960 282202 271012 282208
rect 270868 276752 270920 276758
rect 270868 276694 270920 276700
rect 270776 275460 270828 275466
rect 270776 275402 270828 275408
rect 270684 274100 270736 274106
rect 270684 274042 270736 274048
rect 270592 253428 270644 253434
rect 270592 253370 270644 253376
rect 271064 253366 271092 305798
rect 271156 291990 271184 308450
rect 271432 305454 271460 310420
rect 271616 308582 271644 310420
rect 271604 308576 271656 308582
rect 271604 308518 271656 308524
rect 271420 305448 271472 305454
rect 271420 305390 271472 305396
rect 271800 305386 271828 310420
rect 271788 305380 271840 305386
rect 271788 305322 271840 305328
rect 271144 291984 271196 291990
rect 271144 291926 271196 291932
rect 271984 256222 272012 310420
rect 272168 306490 272196 310420
rect 272168 306462 272288 306490
rect 272156 306400 272208 306406
rect 272156 306342 272208 306348
rect 272064 306332 272116 306338
rect 272064 306274 272116 306280
rect 272076 256290 272104 306274
rect 272168 265810 272196 306342
rect 272260 306218 272288 306462
rect 272352 306406 272380 310420
rect 272340 306400 272392 306406
rect 272340 306342 272392 306348
rect 272536 306338 272564 310420
rect 272720 308446 272748 310420
rect 272708 308440 272760 308446
rect 272708 308382 272760 308388
rect 272524 306332 272576 306338
rect 272524 306274 272576 306280
rect 272260 306190 272380 306218
rect 272248 305856 272300 305862
rect 272248 305798 272300 305804
rect 272260 280974 272288 305798
rect 272248 280968 272300 280974
rect 272248 280910 272300 280916
rect 272156 265804 272208 265810
rect 272156 265746 272208 265752
rect 272064 256284 272116 256290
rect 272064 256226 272116 256232
rect 271972 256216 272024 256222
rect 271972 256158 272024 256164
rect 271052 253360 271104 253366
rect 271052 253302 271104 253308
rect 272352 246702 272380 306190
rect 272904 296714 272932 310420
rect 273088 305862 273116 310420
rect 273272 306354 273300 310420
rect 273456 308514 273484 310420
rect 273444 308508 273496 308514
rect 273444 308450 273496 308456
rect 273272 306326 273484 306354
rect 273076 305856 273128 305862
rect 273076 305798 273128 305804
rect 273352 305856 273404 305862
rect 273352 305798 273404 305804
rect 272444 296686 272932 296714
rect 272444 296002 272472 296686
rect 272432 295996 272484 296002
rect 272432 295938 272484 295944
rect 273364 265878 273392 305798
rect 273456 275534 273484 306326
rect 273548 282334 273576 310490
rect 273654 310406 273852 310434
rect 273720 306400 273772 306406
rect 273720 306342 273772 306348
rect 273628 306332 273680 306338
rect 273628 306274 273680 306280
rect 273640 289270 273668 306274
rect 273628 289264 273680 289270
rect 273628 289206 273680 289212
rect 273536 282328 273588 282334
rect 273536 282270 273588 282276
rect 273444 275528 273496 275534
rect 273444 275470 273496 275476
rect 273352 265872 273404 265878
rect 273352 265814 273404 265820
rect 273732 250782 273760 306342
rect 273824 296070 273852 310406
rect 274100 306338 274128 310420
rect 274088 306332 274140 306338
rect 274088 306274 274140 306280
rect 274284 305862 274312 310420
rect 274468 306406 274496 310420
rect 274456 306400 274508 306406
rect 274456 306342 274508 306348
rect 274652 306354 274680 310420
rect 274836 306354 274864 310420
rect 274652 306326 274772 306354
rect 274836 306326 274956 306354
rect 274272 305856 274324 305862
rect 274272 305798 274324 305804
rect 274640 305856 274692 305862
rect 274640 305798 274692 305804
rect 273812 296064 273864 296070
rect 273812 296006 273864 296012
rect 274652 290630 274680 305798
rect 274744 294710 274772 306326
rect 274824 304020 274876 304026
rect 274824 303962 274876 303968
rect 274732 294704 274784 294710
rect 274732 294646 274784 294652
rect 274640 290624 274692 290630
rect 274640 290566 274692 290572
rect 274836 268462 274864 303962
rect 274928 276826 274956 306326
rect 275020 283694 275048 310420
rect 275204 306354 275232 310420
rect 275112 306326 275232 306354
rect 275112 287774 275140 306326
rect 275388 302234 275416 310420
rect 275204 302206 275416 302234
rect 275100 287768 275152 287774
rect 275100 287710 275152 287716
rect 275008 283688 275060 283694
rect 275008 283630 275060 283636
rect 274916 276820 274968 276826
rect 274916 276762 274968 276768
rect 274824 268456 274876 268462
rect 274824 268398 274876 268404
rect 273720 250776 273772 250782
rect 273720 250718 273772 250724
rect 275204 247994 275232 302206
rect 275572 296714 275600 310420
rect 275756 305862 275784 310420
rect 275744 305856 275796 305862
rect 275744 305798 275796 305804
rect 275836 305652 275888 305658
rect 275836 305594 275888 305600
rect 275848 305386 275876 305594
rect 275836 305380 275888 305386
rect 275836 305322 275888 305328
rect 275940 304026 275968 310420
rect 276124 306354 276152 310420
rect 276032 306326 276152 306354
rect 276308 310406 276414 310434
rect 276204 306332 276256 306338
rect 275928 304020 275980 304026
rect 275928 303962 275980 303968
rect 275296 296686 275600 296714
rect 275296 263022 275324 296686
rect 275284 263016 275336 263022
rect 275284 262958 275336 262964
rect 276032 261662 276060 306326
rect 276204 306274 276256 306280
rect 276216 306218 276244 306274
rect 276124 306190 276244 306218
rect 276124 264314 276152 306190
rect 276308 305862 276336 310406
rect 276584 306354 276612 310420
rect 276400 306326 276612 306354
rect 276768 306338 276796 310420
rect 276756 306332 276808 306338
rect 276296 305856 276348 305862
rect 276296 305798 276348 305804
rect 276296 305652 276348 305658
rect 276296 305594 276348 305600
rect 276204 305448 276256 305454
rect 276204 305390 276256 305396
rect 276216 268530 276244 305390
rect 276308 270026 276336 305594
rect 276400 278254 276428 306326
rect 276756 306274 276808 306280
rect 276952 306082 276980 310420
rect 276492 306054 276980 306082
rect 276492 285190 276520 306054
rect 276848 305856 276900 305862
rect 276848 305798 276900 305804
rect 276860 296714 276888 305798
rect 277136 305658 277164 310420
rect 277124 305652 277176 305658
rect 277124 305594 277176 305600
rect 277320 305454 277348 310420
rect 277400 306468 277452 306474
rect 277400 306410 277452 306416
rect 277308 305448 277360 305454
rect 277308 305390 277360 305396
rect 276584 296686 276888 296714
rect 276584 286550 276612 296686
rect 276572 286544 276624 286550
rect 276572 286486 276624 286492
rect 276480 285184 276532 285190
rect 276480 285126 276532 285132
rect 276388 278248 276440 278254
rect 276388 278190 276440 278196
rect 276296 270020 276348 270026
rect 276296 269962 276348 269968
rect 276204 268524 276256 268530
rect 276204 268466 276256 268472
rect 276112 264308 276164 264314
rect 276112 264250 276164 264256
rect 276020 261656 276072 261662
rect 276020 261598 276072 261604
rect 277412 252006 277440 306410
rect 277504 305862 277532 310420
rect 277584 306332 277636 306338
rect 277584 306274 277636 306280
rect 277492 305856 277544 305862
rect 277492 305798 277544 305804
rect 277492 305652 277544 305658
rect 277492 305594 277544 305600
rect 277504 252074 277532 305594
rect 277596 261730 277624 306274
rect 277688 264382 277716 310420
rect 277872 306474 277900 310420
rect 277860 306468 277912 306474
rect 277860 306410 277912 306416
rect 278056 306354 278084 310420
rect 277780 306326 278084 306354
rect 278240 306338 278268 310420
rect 278228 306332 278280 306338
rect 277780 282402 277808 306326
rect 278228 306274 278280 306280
rect 277860 305856 277912 305862
rect 277860 305798 277912 305804
rect 277872 283762 277900 305798
rect 278424 305658 278452 310420
rect 278412 305652 278464 305658
rect 278412 305594 278464 305600
rect 278608 300257 278636 310420
rect 278806 310406 278912 310434
rect 278780 306468 278832 306474
rect 278780 306410 278832 306416
rect 278594 300248 278650 300257
rect 278594 300183 278650 300192
rect 278792 294778 278820 306410
rect 278884 306338 278912 310406
rect 278976 310406 279082 310434
rect 278872 306332 278924 306338
rect 278872 306274 278924 306280
rect 278872 305652 278924 305658
rect 278872 305594 278924 305600
rect 278780 294772 278832 294778
rect 278780 294714 278832 294720
rect 277860 283756 277912 283762
rect 277860 283698 277912 283704
rect 277768 282396 277820 282402
rect 277768 282338 277820 282344
rect 278884 271318 278912 305594
rect 278976 274174 279004 310406
rect 279056 306400 279108 306406
rect 279056 306342 279108 306348
rect 279252 306354 279280 310420
rect 279436 306406 279464 310420
rect 279424 306400 279476 306406
rect 279068 279682 279096 306342
rect 279148 306332 279200 306338
rect 279252 306326 279372 306354
rect 279424 306342 279476 306348
rect 279148 306274 279200 306280
rect 279160 292058 279188 306274
rect 279240 305856 279292 305862
rect 279240 305798 279292 305804
rect 279148 292052 279200 292058
rect 279148 291994 279200 292000
rect 279056 279676 279108 279682
rect 279056 279618 279108 279624
rect 278964 274168 279016 274174
rect 278964 274110 279016 274116
rect 278872 271312 278924 271318
rect 278872 271254 278924 271260
rect 277676 264376 277728 264382
rect 277676 264318 277728 264324
rect 277584 261724 277636 261730
rect 277584 261666 277636 261672
rect 277492 252068 277544 252074
rect 277492 252010 277544 252016
rect 277400 252000 277452 252006
rect 277400 251942 277452 251948
rect 275192 247988 275244 247994
rect 275192 247930 275244 247936
rect 272340 246696 272392 246702
rect 272340 246638 272392 246644
rect 279252 245206 279280 305798
rect 279344 300393 279372 306326
rect 279620 305658 279648 310420
rect 279804 306474 279832 310420
rect 279792 306468 279844 306474
rect 279792 306410 279844 306416
rect 279988 305862 280016 310420
rect 279976 305856 280028 305862
rect 279976 305798 280028 305804
rect 279608 305652 279660 305658
rect 279608 305594 279660 305600
rect 280172 305454 280200 310420
rect 280356 306474 280384 310420
rect 280344 306468 280396 306474
rect 280344 306410 280396 306416
rect 280540 306218 280568 310420
rect 280448 306190 280568 306218
rect 280448 305946 280476 306190
rect 280356 305918 280476 305946
rect 280252 305652 280304 305658
rect 280252 305594 280304 305600
rect 280160 305448 280212 305454
rect 280160 305390 280212 305396
rect 279330 300384 279386 300393
rect 279330 300319 279386 300328
rect 280264 246770 280292 305594
rect 280356 252142 280384 305918
rect 280436 305856 280488 305862
rect 280436 305798 280488 305804
rect 280448 253570 280476 305798
rect 280528 305448 280580 305454
rect 280528 305390 280580 305396
rect 280540 254930 280568 305390
rect 280724 302234 280752 310420
rect 280804 306468 280856 306474
rect 280804 306410 280856 306416
rect 280632 302206 280752 302234
rect 280632 258738 280660 302206
rect 280816 296714 280844 306410
rect 280908 305658 280936 310420
rect 281092 305862 281120 310420
rect 281276 308786 281304 310420
rect 281264 308780 281316 308786
rect 281264 308722 281316 308728
rect 281080 305856 281132 305862
rect 281080 305798 281132 305804
rect 280896 305652 280948 305658
rect 280896 305594 280948 305600
rect 281552 305386 281580 310420
rect 281736 307018 281764 310420
rect 281724 307012 281776 307018
rect 281724 306954 281776 306960
rect 281920 305946 281948 310420
rect 282000 307012 282052 307018
rect 282000 306954 282052 306960
rect 281644 305918 281948 305946
rect 281540 305380 281592 305386
rect 281540 305322 281592 305328
rect 280724 296686 280844 296714
rect 280620 258732 280672 258738
rect 280620 258674 280672 258680
rect 280528 254924 280580 254930
rect 280528 254866 280580 254872
rect 280436 253564 280488 253570
rect 280436 253506 280488 253512
rect 280344 252136 280396 252142
rect 280344 252078 280396 252084
rect 280252 246764 280304 246770
rect 280252 246706 280304 246712
rect 280724 245274 280752 296686
rect 281644 272746 281672 305918
rect 281816 305856 281868 305862
rect 281816 305798 281868 305804
rect 281724 305652 281776 305658
rect 281724 305594 281776 305600
rect 281736 276894 281764 305594
rect 281828 278322 281856 305798
rect 282012 299474 282040 306954
rect 282104 302841 282132 310420
rect 282288 305862 282316 310420
rect 282276 305856 282328 305862
rect 282276 305798 282328 305804
rect 282090 302832 282146 302841
rect 282090 302767 282146 302776
rect 281920 299446 282040 299474
rect 281920 287910 281948 299446
rect 282472 296714 282500 310420
rect 282656 302977 282684 310420
rect 282840 305658 282868 310420
rect 283024 308224 283052 310420
rect 282932 308196 283052 308224
rect 282932 307902 282960 308196
rect 283208 308156 283236 310420
rect 283024 308128 283236 308156
rect 282920 307896 282972 307902
rect 282920 307838 282972 307844
rect 282920 307760 282972 307766
rect 282920 307702 282972 307708
rect 282828 305652 282880 305658
rect 282828 305594 282880 305600
rect 282642 302968 282698 302977
rect 282642 302903 282698 302912
rect 282932 301510 282960 307702
rect 283024 304298 283052 308128
rect 283392 307986 283420 310420
rect 283208 307958 283420 307986
rect 283104 307080 283156 307086
rect 283104 307022 283156 307028
rect 283012 304292 283064 304298
rect 283012 304234 283064 304240
rect 282920 301504 282972 301510
rect 282920 301446 282972 301452
rect 282196 296686 282500 296714
rect 281908 287904 281960 287910
rect 281908 287846 281960 287852
rect 281816 278316 281868 278322
rect 281816 278258 281868 278264
rect 281724 276888 281776 276894
rect 281724 276830 281776 276836
rect 281632 272740 281684 272746
rect 281632 272682 281684 272688
rect 282196 249422 282224 296686
rect 283116 275602 283144 307022
rect 283208 286618 283236 307958
rect 283288 307896 283340 307902
rect 283288 307838 283340 307844
rect 283380 307896 283432 307902
rect 283380 307838 283432 307844
rect 283300 290698 283328 307838
rect 283288 290692 283340 290698
rect 283288 290634 283340 290640
rect 283196 286612 283248 286618
rect 283196 286554 283248 286560
rect 283104 275596 283156 275602
rect 283104 275538 283156 275544
rect 282184 249416 282236 249422
rect 282184 249358 282236 249364
rect 283392 245342 283420 307838
rect 283576 296714 283604 310420
rect 283760 307766 283788 310420
rect 283748 307760 283800 307766
rect 283748 307702 283800 307708
rect 283944 307086 283972 310420
rect 284036 310406 284234 310434
rect 284036 307902 284064 310406
rect 284300 308440 284352 308446
rect 284300 308382 284352 308388
rect 284024 307896 284076 307902
rect 284024 307838 284076 307844
rect 283932 307080 283984 307086
rect 283932 307022 283984 307028
rect 284312 306374 284340 308382
rect 284404 307834 284432 310420
rect 284588 308394 284616 310420
rect 284496 308366 284616 308394
rect 284392 307828 284444 307834
rect 284392 307770 284444 307776
rect 284312 306346 284432 306374
rect 283484 296686 283604 296714
rect 283484 265946 283512 296686
rect 284404 272814 284432 306346
rect 284496 274242 284524 308366
rect 284772 308292 284800 310420
rect 284588 308264 284800 308292
rect 284588 281042 284616 308264
rect 284668 308168 284720 308174
rect 284668 308110 284720 308116
rect 284680 293418 284708 308110
rect 284760 308100 284812 308106
rect 284760 308042 284812 308048
rect 284668 293412 284720 293418
rect 284668 293354 284720 293360
rect 284576 281036 284628 281042
rect 284576 280978 284628 280984
rect 284484 274236 284536 274242
rect 284484 274178 284536 274184
rect 284392 272808 284444 272814
rect 284392 272750 284444 272756
rect 283472 265940 283524 265946
rect 283472 265882 283524 265888
rect 284772 248062 284800 308042
rect 284852 307828 284904 307834
rect 284852 307770 284904 307776
rect 284864 305726 284892 307770
rect 284956 307154 284984 310420
rect 285140 308446 285168 310420
rect 285128 308440 285180 308446
rect 285128 308382 285180 308388
rect 285324 308106 285352 310420
rect 285508 308174 285536 310420
rect 285496 308168 285548 308174
rect 285496 308110 285548 308116
rect 285312 308100 285364 308106
rect 285312 308042 285364 308048
rect 285692 307902 285720 310420
rect 285876 308174 285904 310420
rect 286060 308292 286088 310420
rect 286140 308440 286192 308446
rect 286140 308382 286192 308388
rect 285968 308264 286088 308292
rect 285864 308168 285916 308174
rect 285864 308110 285916 308116
rect 285968 307986 285996 308264
rect 286048 308168 286100 308174
rect 286048 308110 286100 308116
rect 285784 307958 285996 307986
rect 285680 307896 285732 307902
rect 285680 307838 285732 307844
rect 285680 307760 285732 307766
rect 285680 307702 285732 307708
rect 284944 307148 284996 307154
rect 284944 307090 284996 307096
rect 284852 305720 284904 305726
rect 284852 305662 284904 305668
rect 285692 296138 285720 307702
rect 285784 304434 285812 307958
rect 285956 307896 286008 307902
rect 285956 307838 286008 307844
rect 285864 307828 285916 307834
rect 285864 307770 285916 307776
rect 285772 304428 285824 304434
rect 285772 304370 285824 304376
rect 285680 296132 285732 296138
rect 285680 296074 285732 296080
rect 285876 283830 285904 307770
rect 285968 284889 285996 307838
rect 286060 289338 286088 308110
rect 286048 289332 286100 289338
rect 286048 289274 286100 289280
rect 285954 284880 286010 284889
rect 285954 284815 286010 284824
rect 285864 283824 285916 283830
rect 285864 283766 285916 283772
rect 286152 250850 286180 308382
rect 286244 271386 286272 310420
rect 286428 308446 286456 310420
rect 286520 310406 286718 310434
rect 286416 308440 286468 308446
rect 286416 308382 286468 308388
rect 286520 307766 286548 310406
rect 286888 307834 286916 310420
rect 286968 310004 287020 310010
rect 286968 309946 287020 309952
rect 286980 309482 287008 309946
rect 287072 309618 287100 310420
rect 287072 309590 287192 309618
rect 286980 309454 287100 309482
rect 286876 307828 286928 307834
rect 286876 307770 286928 307776
rect 286508 307760 286560 307766
rect 286508 307702 286560 307708
rect 286232 271380 286284 271386
rect 286232 271322 286284 271328
rect 286140 250844 286192 250850
rect 286140 250786 286192 250792
rect 287072 250481 287100 309454
rect 287164 308650 287192 309590
rect 287256 308718 287284 310420
rect 287244 308712 287296 308718
rect 287244 308654 287296 308660
rect 287152 308644 287204 308650
rect 287152 308586 287204 308592
rect 287440 308530 287468 310420
rect 287624 310010 287652 310420
rect 287612 310004 287664 310010
rect 287612 309946 287664 309952
rect 287520 308712 287572 308718
rect 287520 308654 287572 308660
rect 287164 308502 287468 308530
rect 287164 255921 287192 308502
rect 287336 308304 287388 308310
rect 287336 308246 287388 308252
rect 287428 308304 287480 308310
rect 287428 308246 287480 308252
rect 287244 308236 287296 308242
rect 287244 308178 287296 308184
rect 287256 257650 287284 308178
rect 287348 261798 287376 308246
rect 287440 295118 287468 308246
rect 287532 303249 287560 308654
rect 287808 308514 287836 310420
rect 287992 308514 288020 310420
rect 287796 308508 287848 308514
rect 287796 308450 287848 308456
rect 287980 308508 288032 308514
rect 287980 308450 288032 308456
rect 288176 308394 288204 310420
rect 287624 308366 288204 308394
rect 287624 303385 287652 308366
rect 288360 306241 288388 310420
rect 288544 308650 288572 310420
rect 288532 308644 288584 308650
rect 288532 308586 288584 308592
rect 288728 308530 288756 310420
rect 288452 308502 288756 308530
rect 288346 306232 288402 306241
rect 288346 306167 288402 306176
rect 288452 303618 288480 308502
rect 288808 308440 288860 308446
rect 288808 308382 288860 308388
rect 288532 308372 288584 308378
rect 288532 308314 288584 308320
rect 288544 306270 288572 308314
rect 288624 308304 288676 308310
rect 288624 308246 288676 308252
rect 288532 306264 288584 306270
rect 288532 306206 288584 306212
rect 288440 303612 288492 303618
rect 288440 303554 288492 303560
rect 287610 303376 287666 303385
rect 287610 303311 287666 303320
rect 287518 303240 287574 303249
rect 287518 303175 287574 303184
rect 288636 302870 288664 308246
rect 288716 308236 288768 308242
rect 288716 308178 288768 308184
rect 288728 305969 288756 308178
rect 288714 305960 288770 305969
rect 288714 305895 288770 305904
rect 288624 302864 288676 302870
rect 288624 302806 288676 302812
rect 288820 302802 288848 308382
rect 288912 306105 288940 310420
rect 289096 308310 289124 310420
rect 289188 310406 289386 310434
rect 289084 308304 289136 308310
rect 289084 308246 289136 308252
rect 288898 306096 288954 306105
rect 288898 306031 288954 306040
rect 288808 302796 288860 302802
rect 288808 302738 288860 302744
rect 289188 302734 289216 310406
rect 289556 308242 289584 310420
rect 289740 308446 289768 310420
rect 289820 308508 289872 308514
rect 289820 308450 289872 308456
rect 289728 308440 289780 308446
rect 289728 308382 289780 308388
rect 289544 308236 289596 308242
rect 289544 308178 289596 308184
rect 289832 307986 289860 308450
rect 289924 308122 289952 310420
rect 289924 308094 290044 308122
rect 289832 307958 289952 307986
rect 289820 307896 289872 307902
rect 289820 307838 289872 307844
rect 289832 305522 289860 307838
rect 289820 305516 289872 305522
rect 289820 305458 289872 305464
rect 289924 303346 289952 307958
rect 289912 303340 289964 303346
rect 289912 303282 289964 303288
rect 289176 302728 289228 302734
rect 289176 302670 289228 302676
rect 290016 300529 290044 308094
rect 290108 305833 290136 310420
rect 290292 308514 290320 310420
rect 290280 308508 290332 308514
rect 290280 308450 290332 308456
rect 290476 308394 290504 310420
rect 290200 308366 290504 308394
rect 290094 305824 290150 305833
rect 290094 305759 290150 305768
rect 290002 300520 290058 300529
rect 290002 300455 290058 300464
rect 290200 297673 290228 308366
rect 290280 308304 290332 308310
rect 290280 308246 290332 308252
rect 290186 297664 290242 297673
rect 290186 297599 290242 297608
rect 290292 297401 290320 308246
rect 290660 307902 290688 310420
rect 290648 307896 290700 307902
rect 290648 307838 290700 307844
rect 290844 303550 290872 310420
rect 291028 308310 291056 310420
rect 291212 308310 291240 310420
rect 291292 308508 291344 308514
rect 291292 308450 291344 308456
rect 291016 308304 291068 308310
rect 291016 308246 291068 308252
rect 291200 308304 291252 308310
rect 291200 308246 291252 308252
rect 291200 308168 291252 308174
rect 291200 308110 291252 308116
rect 290832 303544 290884 303550
rect 290832 303486 290884 303492
rect 291212 303278 291240 308110
rect 291304 305590 291332 308450
rect 291292 305584 291344 305590
rect 291292 305526 291344 305532
rect 291200 303272 291252 303278
rect 291200 303214 291252 303220
rect 291396 303210 291424 310420
rect 291476 308440 291528 308446
rect 291476 308382 291528 308388
rect 291488 306134 291516 308382
rect 291476 306128 291528 306134
rect 291476 306070 291528 306076
rect 291384 303204 291436 303210
rect 291384 303146 291436 303152
rect 291580 297537 291608 310420
rect 291672 310406 291870 310434
rect 291672 308514 291700 310406
rect 291660 308508 291712 308514
rect 291660 308450 291712 308456
rect 291660 308372 291712 308378
rect 291660 308314 291712 308320
rect 291566 297528 291622 297537
rect 291566 297463 291622 297472
rect 290278 297392 290334 297401
rect 291672 297362 291700 308314
rect 291752 308304 291804 308310
rect 291752 308246 291804 308252
rect 291764 305697 291792 308246
rect 292040 308174 292068 310420
rect 292224 308378 292252 310420
rect 292408 308446 292436 310420
rect 292396 308440 292448 308446
rect 292396 308382 292448 308388
rect 292212 308372 292264 308378
rect 292212 308314 292264 308320
rect 292028 308168 292080 308174
rect 292028 308110 292080 308116
rect 291750 305688 291806 305697
rect 291750 305623 291806 305632
rect 292592 303142 292620 310420
rect 292776 305946 292804 310420
rect 292960 306066 292988 310420
rect 293144 306082 293172 310420
rect 292948 306060 293000 306066
rect 293144 306054 293264 306082
rect 292948 306002 293000 306008
rect 292776 305918 293172 305946
rect 293040 305856 293092 305862
rect 293040 305798 293092 305804
rect 292948 305788 293000 305794
rect 292948 305730 293000 305736
rect 292580 303136 292632 303142
rect 292580 303078 292632 303084
rect 292960 297430 292988 305730
rect 293052 297770 293080 305798
rect 293144 302122 293172 305918
rect 293236 303414 293264 306054
rect 293224 303408 293276 303414
rect 293224 303350 293276 303356
rect 293132 302116 293184 302122
rect 293132 302058 293184 302064
rect 293328 297809 293356 310420
rect 293512 306202 293540 310420
rect 293500 306196 293552 306202
rect 293500 306138 293552 306144
rect 293696 305862 293724 310420
rect 293684 305856 293736 305862
rect 293684 305798 293736 305804
rect 293880 305794 293908 310420
rect 294064 305998 294092 310420
rect 294262 310406 294460 310434
rect 294144 306400 294196 306406
rect 294144 306342 294196 306348
rect 294052 305992 294104 305998
rect 294052 305934 294104 305940
rect 293868 305788 293920 305794
rect 293868 305730 293920 305736
rect 293314 297800 293370 297809
rect 293040 297764 293092 297770
rect 293314 297735 293370 297744
rect 293040 297706 293092 297712
rect 294156 297702 294184 306342
rect 294328 306332 294380 306338
rect 294328 306274 294380 306280
rect 294236 306264 294288 306270
rect 294236 306206 294288 306212
rect 294144 297696 294196 297702
rect 294144 297638 294196 297644
rect 292948 297424 293000 297430
rect 292948 297366 293000 297372
rect 290278 297327 290334 297336
rect 291660 297356 291712 297362
rect 291660 297298 291712 297304
rect 294248 297226 294276 306206
rect 294236 297220 294288 297226
rect 294236 297162 294288 297168
rect 287428 295112 287480 295118
rect 287428 295054 287480 295060
rect 294340 295050 294368 306274
rect 294432 297634 294460 310406
rect 294524 302938 294552 310420
rect 294512 302932 294564 302938
rect 294512 302874 294564 302880
rect 294420 297628 294472 297634
rect 294420 297570 294472 297576
rect 294708 297498 294736 310420
rect 294892 306406 294920 310420
rect 294880 306400 294932 306406
rect 294880 306342 294932 306348
rect 295076 306338 295104 310420
rect 295064 306332 295116 306338
rect 295064 306274 295116 306280
rect 295260 306270 295288 310420
rect 295444 306626 295472 310420
rect 295628 306746 295656 310420
rect 295616 306740 295668 306746
rect 295616 306682 295668 306688
rect 295812 306626 295840 310420
rect 295444 306598 295748 306626
rect 295812 306598 295932 306626
rect 295720 306490 295748 306598
rect 295616 306468 295668 306474
rect 295720 306462 295840 306490
rect 295616 306410 295668 306416
rect 295432 306400 295484 306406
rect 295432 306342 295484 306348
rect 295248 306264 295300 306270
rect 295248 306206 295300 306212
rect 295444 301782 295472 306342
rect 295524 306332 295576 306338
rect 295628 306320 295656 306410
rect 295628 306292 295748 306320
rect 295524 306274 295576 306280
rect 295536 301850 295564 306274
rect 295616 306196 295668 306202
rect 295616 306138 295668 306144
rect 295524 301844 295576 301850
rect 295524 301786 295576 301792
rect 295432 301776 295484 301782
rect 295432 301718 295484 301724
rect 295628 301578 295656 306138
rect 295616 301572 295668 301578
rect 295616 301514 295668 301520
rect 294696 297492 294748 297498
rect 294696 297434 294748 297440
rect 295720 295186 295748 306292
rect 295812 297294 295840 306462
rect 295904 305726 295932 306598
rect 295996 306338 296024 310420
rect 296180 306406 296208 310420
rect 296168 306400 296220 306406
rect 296168 306342 296220 306348
rect 295984 306332 296036 306338
rect 295984 306274 296036 306280
rect 296364 306202 296392 310420
rect 296352 306196 296404 306202
rect 296352 306138 296404 306144
rect 295892 305720 295944 305726
rect 295892 305662 295944 305668
rect 296548 301986 296576 310420
rect 296536 301980 296588 301986
rect 296536 301922 296588 301928
rect 296732 301918 296760 310420
rect 296916 310406 297022 310434
rect 296812 306332 296864 306338
rect 296812 306274 296864 306280
rect 296824 302054 296852 306274
rect 296812 302048 296864 302054
rect 296812 301990 296864 301996
rect 296720 301912 296772 301918
rect 296720 301854 296772 301860
rect 295800 297288 295852 297294
rect 295800 297230 295852 297236
rect 295708 295180 295760 295186
rect 295708 295122 295760 295128
rect 294328 295044 294380 295050
rect 294328 294986 294380 294992
rect 296916 294846 296944 310406
rect 297192 307018 297220 310420
rect 297180 307012 297232 307018
rect 297180 306954 297232 306960
rect 297088 306808 297140 306814
rect 297088 306750 297140 306756
rect 296996 300620 297048 300626
rect 296996 300562 297048 300568
rect 297008 294982 297036 300562
rect 296996 294976 297048 294982
rect 296996 294918 297048 294924
rect 297100 294914 297128 306750
rect 297180 302524 297232 302530
rect 297180 302466 297232 302472
rect 297088 294908 297140 294914
rect 297088 294850 297140 294856
rect 296904 294840 296956 294846
rect 296904 294782 296956 294788
rect 287336 261792 287388 261798
rect 287336 261734 287388 261740
rect 287244 257644 287296 257650
rect 287244 257586 287296 257592
rect 287150 255912 287206 255921
rect 287150 255847 287206 255856
rect 287058 250472 287114 250481
rect 287058 250407 287114 250416
rect 284760 248056 284812 248062
rect 284760 247998 284812 248004
rect 283380 245336 283432 245342
rect 283380 245278 283432 245284
rect 280712 245268 280764 245274
rect 280712 245210 280764 245216
rect 279240 245200 279292 245206
rect 279240 245142 279292 245148
rect 269672 245132 269724 245138
rect 269672 245074 269724 245080
rect 268292 245064 268344 245070
rect 268292 245006 268344 245012
rect 262772 244996 262824 245002
rect 262772 244938 262824 244944
rect 250444 244928 250496 244934
rect 250444 244870 250496 244876
rect 297192 243642 297220 302466
rect 297376 300626 297404 310420
rect 297560 306338 297588 310420
rect 297548 306332 297600 306338
rect 297548 306274 297600 306280
rect 297364 300620 297416 300626
rect 297364 300562 297416 300568
rect 297744 296714 297772 310420
rect 297928 302530 297956 310420
rect 298112 305969 298140 310420
rect 298296 308417 298324 310420
rect 298282 308408 298338 308417
rect 298282 308343 298338 308352
rect 298098 305960 298154 305969
rect 298480 305930 298508 310420
rect 298560 306332 298612 306338
rect 298560 306274 298612 306280
rect 298098 305895 298154 305904
rect 298468 305924 298520 305930
rect 298468 305866 298520 305872
rect 297916 302524 297968 302530
rect 297916 302466 297968 302472
rect 297284 296686 297772 296714
rect 297180 243636 297232 243642
rect 297180 243578 297232 243584
rect 297284 243574 297312 296686
rect 298572 243778 298600 306274
rect 298560 243772 298612 243778
rect 298560 243714 298612 243720
rect 297272 243568 297324 243574
rect 298664 243545 298692 310420
rect 298848 303385 298876 310420
rect 298834 303376 298890 303385
rect 298834 303311 298890 303320
rect 299032 303074 299060 310420
rect 299216 306338 299244 310420
rect 299204 306332 299256 306338
rect 299204 306274 299256 306280
rect 299020 303068 299072 303074
rect 299020 303010 299072 303016
rect 299400 302938 299428 310420
rect 299676 308446 299704 310420
rect 299664 308440 299716 308446
rect 299664 308382 299716 308388
rect 299572 306400 299624 306406
rect 299572 306342 299624 306348
rect 299480 306332 299532 306338
rect 299480 306274 299532 306280
rect 299388 302932 299440 302938
rect 299388 302874 299440 302880
rect 299492 243846 299520 306274
rect 299480 243840 299532 243846
rect 299480 243782 299532 243788
rect 299584 243574 299612 306342
rect 299860 306320 299888 310420
rect 299676 306292 299888 306320
rect 299676 243914 299704 306292
rect 300044 302234 300072 310420
rect 299768 302206 300072 302234
rect 299768 300121 299796 302206
rect 300228 300490 300256 310420
rect 300412 306338 300440 310420
rect 300596 306406 300624 310420
rect 300780 308514 300808 310420
rect 300768 308508 300820 308514
rect 300768 308450 300820 308456
rect 300860 306740 300912 306746
rect 300860 306682 300912 306688
rect 300584 306400 300636 306406
rect 300584 306342 300636 306348
rect 300400 306332 300452 306338
rect 300400 306274 300452 306280
rect 300216 300484 300268 300490
rect 300216 300426 300268 300432
rect 299754 300112 299810 300121
rect 299754 300047 299810 300056
rect 299664 243908 299716 243914
rect 299664 243850 299716 243856
rect 300872 243710 300900 306682
rect 300964 306626 300992 310420
rect 301148 306746 301176 310420
rect 301136 306740 301188 306746
rect 301136 306682 301188 306688
rect 300964 306598 301268 306626
rect 301044 306400 301096 306406
rect 301044 306342 301096 306348
rect 300952 303748 301004 303754
rect 300952 303690 301004 303696
rect 300860 243704 300912 243710
rect 300860 243646 300912 243652
rect 300964 243642 300992 303690
rect 301056 253638 301084 306342
rect 301136 306332 301188 306338
rect 301136 306274 301188 306280
rect 301148 253706 301176 306274
rect 301240 303006 301268 306598
rect 301228 303000 301280 303006
rect 301228 302942 301280 302948
rect 301332 302234 301360 310420
rect 301516 306338 301544 310420
rect 301700 308582 301728 310420
rect 301688 308576 301740 308582
rect 301688 308518 301740 308524
rect 301504 306332 301556 306338
rect 301504 306274 301556 306280
rect 301884 303754 301912 310420
rect 302068 306406 302096 310420
rect 302344 308650 302372 310420
rect 302332 308644 302384 308650
rect 302332 308586 302384 308592
rect 302056 306400 302108 306406
rect 302528 306354 302556 310420
rect 302712 308718 302740 310420
rect 302700 308712 302752 308718
rect 302700 308654 302752 308660
rect 302056 306342 302108 306348
rect 302240 306332 302292 306338
rect 302240 306274 302292 306280
rect 302344 306326 302556 306354
rect 301872 303748 301924 303754
rect 301872 303690 301924 303696
rect 301240 302206 301360 302234
rect 301240 300354 301268 302206
rect 301228 300348 301280 300354
rect 301228 300290 301280 300296
rect 301136 253700 301188 253706
rect 301136 253642 301188 253648
rect 301044 253632 301096 253638
rect 301044 253574 301096 253580
rect 302252 245274 302280 306274
rect 302344 247994 302372 306326
rect 302896 306218 302924 310420
rect 302436 306190 302924 306218
rect 302436 248334 302464 306190
rect 302516 304020 302568 304026
rect 302516 303962 302568 303968
rect 302424 248328 302476 248334
rect 302424 248270 302476 248276
rect 302528 248062 302556 303962
rect 303080 296714 303108 310420
rect 303264 306338 303292 310420
rect 303252 306332 303304 306338
rect 303252 306274 303304 306280
rect 303448 304026 303476 310420
rect 303436 304020 303488 304026
rect 303436 303962 303488 303968
rect 302620 296686 303108 296714
rect 302620 253842 302648 296686
rect 302608 253836 302660 253842
rect 302608 253778 302660 253784
rect 302516 248056 302568 248062
rect 302516 247998 302568 248004
rect 302332 247988 302384 247994
rect 302332 247930 302384 247936
rect 302240 245268 302292 245274
rect 302240 245210 302292 245216
rect 303632 243681 303660 310420
rect 303816 308786 303844 310420
rect 303804 308780 303856 308786
rect 303804 308722 303856 308728
rect 304000 306354 304028 310420
rect 303804 306332 303856 306338
rect 303804 306274 303856 306280
rect 303908 306326 304028 306354
rect 303712 302864 303764 302870
rect 303712 302806 303764 302812
rect 303724 247586 303752 302806
rect 303816 250481 303844 306274
rect 303908 250782 303936 306326
rect 303988 306264 304040 306270
rect 303988 306206 304040 306212
rect 304000 250889 304028 306206
rect 304184 296714 304212 310420
rect 304368 306338 304396 310420
rect 304356 306332 304408 306338
rect 304356 306274 304408 306280
rect 304552 302870 304580 310420
rect 304644 310406 304842 310434
rect 304644 306270 304672 310406
rect 304632 306264 304684 306270
rect 304632 306206 304684 306212
rect 305012 306134 305040 310420
rect 305092 306468 305144 306474
rect 305092 306410 305144 306416
rect 305000 306128 305052 306134
rect 305000 306070 305052 306076
rect 305000 305992 305052 305998
rect 305000 305934 305052 305940
rect 304540 302864 304592 302870
rect 304540 302806 304592 302812
rect 304092 296686 304212 296714
rect 304092 253774 304120 296686
rect 304080 253768 304132 253774
rect 304080 253710 304132 253716
rect 303986 250880 304042 250889
rect 303986 250815 304042 250824
rect 303896 250776 303948 250782
rect 303896 250718 303948 250724
rect 303802 250472 303858 250481
rect 303802 250407 303858 250416
rect 303712 247580 303764 247586
rect 303712 247522 303764 247528
rect 305012 244905 305040 305934
rect 305104 248198 305132 306410
rect 305196 306354 305224 310420
rect 305196 306326 305316 306354
rect 305184 306264 305236 306270
rect 305184 306206 305236 306212
rect 305092 248192 305144 248198
rect 305092 248134 305144 248140
rect 305196 245041 305224 306206
rect 305288 248169 305316 306326
rect 305380 306218 305408 310420
rect 305564 306490 305592 310420
rect 305472 306462 305592 306490
rect 305748 306474 305776 310420
rect 305736 306468 305788 306474
rect 305472 306338 305500 306462
rect 305736 306410 305788 306416
rect 305460 306332 305512 306338
rect 305460 306274 305512 306280
rect 305380 306190 305684 306218
rect 305368 306128 305420 306134
rect 305368 306070 305420 306076
rect 305460 306128 305512 306134
rect 305460 306070 305512 306076
rect 305274 248160 305330 248169
rect 305274 248095 305330 248104
rect 305380 245177 305408 306070
rect 305472 248130 305500 306070
rect 305552 299736 305604 299742
rect 305552 299678 305604 299684
rect 305564 250918 305592 299678
rect 305552 250912 305604 250918
rect 305552 250854 305604 250860
rect 305656 250374 305684 306190
rect 305932 299742 305960 310420
rect 306116 305998 306144 310420
rect 306300 306134 306328 310420
rect 306484 306490 306512 310420
rect 306392 306462 306512 306490
rect 306288 306128 306340 306134
rect 306288 306070 306340 306076
rect 306104 305992 306156 305998
rect 306104 305934 306156 305940
rect 306392 305862 306420 306462
rect 306668 306354 306696 310420
rect 306484 306326 306696 306354
rect 306380 305856 306432 305862
rect 306380 305798 306432 305804
rect 306380 305720 306432 305726
rect 306380 305662 306432 305668
rect 305920 299736 305972 299742
rect 305920 299678 305972 299684
rect 305644 250368 305696 250374
rect 305644 250310 305696 250316
rect 305460 248124 305512 248130
rect 305460 248066 305512 248072
rect 306392 245342 306420 305662
rect 306380 245336 306432 245342
rect 306484 245313 306512 306326
rect 306564 306264 306616 306270
rect 306852 306218 306880 310420
rect 306564 306206 306616 306212
rect 306576 248266 306604 306206
rect 306668 306190 306880 306218
rect 306668 248402 306696 306190
rect 307036 306082 307064 310420
rect 306760 306054 307064 306082
rect 306760 251122 306788 306054
rect 306840 305992 306892 305998
rect 306840 305934 306892 305940
rect 306748 251116 306800 251122
rect 306748 251058 306800 251064
rect 306852 251054 306880 305934
rect 306932 305856 306984 305862
rect 306932 305798 306984 305804
rect 306840 251048 306892 251054
rect 306840 250990 306892 250996
rect 306944 250986 306972 305798
rect 307220 305726 307248 310420
rect 307312 310406 307510 310434
rect 307312 306474 307340 310406
rect 307300 306468 307352 306474
rect 307300 306410 307352 306416
rect 307680 305998 307708 310420
rect 307864 306354 307892 310420
rect 307944 306468 307996 306474
rect 307944 306410 307996 306416
rect 307772 306326 307892 306354
rect 307668 305992 307720 305998
rect 307668 305934 307720 305940
rect 307208 305720 307260 305726
rect 307208 305662 307260 305668
rect 306932 250980 306984 250986
rect 306932 250922 306984 250928
rect 306656 248396 306708 248402
rect 306656 248338 306708 248344
rect 306564 248260 306616 248266
rect 306564 248202 306616 248208
rect 307772 245478 307800 306326
rect 307956 306218 307984 306410
rect 307864 306190 307984 306218
rect 307760 245472 307812 245478
rect 307760 245414 307812 245420
rect 307864 245410 307892 306190
rect 307944 306128 307996 306134
rect 307944 306070 307996 306076
rect 307956 245546 307984 306070
rect 308048 247654 308076 310420
rect 308232 306354 308260 310420
rect 308416 306474 308444 310420
rect 308404 306468 308456 306474
rect 308404 306410 308456 306416
rect 308128 306332 308180 306338
rect 308232 306326 308444 306354
rect 308600 306338 308628 310420
rect 308128 306274 308180 306280
rect 308140 247761 308168 306274
rect 308220 306264 308272 306270
rect 308220 306206 308272 306212
rect 308232 250617 308260 306206
rect 308416 250753 308444 306326
rect 308588 306332 308640 306338
rect 308588 306274 308640 306280
rect 308784 306270 308812 310420
rect 308772 306264 308824 306270
rect 308772 306206 308824 306212
rect 308968 306134 308996 310420
rect 309152 306354 309180 310420
rect 309336 306610 309364 310420
rect 309324 306604 309376 306610
rect 309324 306546 309376 306552
rect 309520 306490 309548 310420
rect 309336 306462 309548 306490
rect 309152 306326 309272 306354
rect 309140 306196 309192 306202
rect 309140 306138 309192 306144
rect 308956 306128 309008 306134
rect 308956 306070 309008 306076
rect 308402 250744 308458 250753
rect 308402 250679 308458 250688
rect 308218 250608 308274 250617
rect 308218 250543 308274 250552
rect 308126 247752 308182 247761
rect 308126 247687 308182 247696
rect 308036 247648 308088 247654
rect 308036 247590 308088 247596
rect 309152 245585 309180 306138
rect 309244 248033 309272 306326
rect 309230 248024 309286 248033
rect 309230 247959 309286 247968
rect 309138 245576 309194 245585
rect 307944 245540 307996 245546
rect 309138 245511 309194 245520
rect 307944 245482 307996 245488
rect 309336 245449 309364 306462
rect 309704 306354 309732 310420
rect 309428 306326 309732 306354
rect 309796 310406 309994 310434
rect 309428 247897 309456 306326
rect 309508 306264 309560 306270
rect 309508 306206 309560 306212
rect 309520 251190 309548 306206
rect 309796 296714 309824 310406
rect 310164 306202 310192 310420
rect 310348 308990 310376 310420
rect 310336 308984 310388 308990
rect 310336 308926 310388 308932
rect 310152 306196 310204 306202
rect 310152 306138 310204 306144
rect 309612 296686 309824 296714
rect 309508 251184 309560 251190
rect 309508 251126 309560 251132
rect 309612 250442 309640 296686
rect 309600 250436 309652 250442
rect 309600 250378 309652 250384
rect 309414 247888 309470 247897
rect 309414 247823 309470 247832
rect 309322 245440 309378 245449
rect 307852 245404 307904 245410
rect 309322 245375 309378 245384
rect 307852 245346 307904 245352
rect 306380 245278 306432 245284
rect 306470 245304 306526 245313
rect 306470 245239 306526 245248
rect 305366 245168 305422 245177
rect 305366 245103 305422 245112
rect 305182 245032 305238 245041
rect 305182 244967 305238 244976
rect 304998 244896 305054 244905
rect 304998 244831 305054 244840
rect 310532 244769 310560 310420
rect 310612 306468 310664 306474
rect 310612 306410 310664 306416
rect 310624 248305 310652 306410
rect 310716 306354 310744 310420
rect 310900 306474 310928 310420
rect 311084 308553 311112 310420
rect 311070 308544 311126 308553
rect 311070 308479 311126 308488
rect 310888 306468 310940 306474
rect 310888 306410 310940 306416
rect 310716 306326 310928 306354
rect 310704 306264 310756 306270
rect 310704 306206 310756 306212
rect 310716 251841 310744 306206
rect 310796 306196 310848 306202
rect 310796 306138 310848 306144
rect 310808 253201 310836 306138
rect 310794 253192 310850 253201
rect 310794 253127 310850 253136
rect 310900 251977 310928 306326
rect 310980 306332 311032 306338
rect 310980 306274 311032 306280
rect 310992 254697 311020 306274
rect 311268 306270 311296 310420
rect 311256 306264 311308 306270
rect 311256 306206 311308 306212
rect 311452 296714 311480 310420
rect 311636 306338 311664 310420
rect 311624 306332 311676 306338
rect 311624 306274 311676 306280
rect 311820 306202 311848 310420
rect 311900 306468 311952 306474
rect 311900 306410 311952 306416
rect 311808 306196 311860 306202
rect 311808 306138 311860 306144
rect 311084 296686 311480 296714
rect 311084 258777 311112 296686
rect 311070 258768 311126 258777
rect 311070 258703 311126 258712
rect 310978 254688 311034 254697
rect 310978 254623 311034 254632
rect 310886 251968 310942 251977
rect 310886 251903 310942 251912
rect 310702 251832 310758 251841
rect 310702 251767 310758 251776
rect 311912 250850 311940 306410
rect 312004 306320 312032 310420
rect 312188 308922 312216 310420
rect 312176 308916 312228 308922
rect 312176 308858 312228 308864
rect 312004 306292 312124 306320
rect 311992 306196 312044 306202
rect 311992 306138 312044 306144
rect 312004 285122 312032 306138
rect 312096 286385 312124 306292
rect 312372 303521 312400 310420
rect 312464 310406 312662 310434
rect 312464 306474 312492 310406
rect 312452 306468 312504 306474
rect 312452 306410 312504 306416
rect 312358 303512 312414 303521
rect 312358 303447 312414 303456
rect 312832 303362 312860 310420
rect 312188 303334 312860 303362
rect 312188 296274 312216 303334
rect 313016 302234 313044 310420
rect 313200 306202 313228 310420
rect 313280 306400 313332 306406
rect 313280 306342 313332 306348
rect 313188 306196 313240 306202
rect 313188 306138 313240 306144
rect 312280 302206 313044 302234
rect 312280 301782 312308 302206
rect 312268 301776 312320 301782
rect 312268 301718 312320 301724
rect 312176 296268 312228 296274
rect 312176 296210 312228 296216
rect 312082 286376 312138 286385
rect 312082 286311 312138 286320
rect 311992 285116 312044 285122
rect 311992 285058 312044 285064
rect 313292 254561 313320 306342
rect 313384 306320 313412 310420
rect 313568 306338 313596 310420
rect 313556 306332 313608 306338
rect 313384 306292 313504 306320
rect 313372 306128 313424 306134
rect 313372 306070 313424 306076
rect 313384 265878 313412 306070
rect 313476 282402 313504 306292
rect 313556 306274 313608 306280
rect 313556 306196 313608 306202
rect 313556 306138 313608 306144
rect 313568 287978 313596 306138
rect 313752 302234 313780 310420
rect 313936 306406 313964 310420
rect 314120 307222 314148 310420
rect 314108 307216 314160 307222
rect 314108 307158 314160 307164
rect 313924 306400 313976 306406
rect 313924 306342 313976 306348
rect 313832 306332 313884 306338
rect 313832 306274 313884 306280
rect 313660 302206 313780 302234
rect 313660 299062 313688 302206
rect 313844 300422 313872 306274
rect 314304 306202 314332 310420
rect 314292 306196 314344 306202
rect 314292 306138 314344 306144
rect 314488 306134 314516 310420
rect 314672 306134 314700 310420
rect 314948 310406 315146 310434
rect 314752 306332 314804 306338
rect 314948 306320 314976 310406
rect 315316 306320 315344 310420
rect 314752 306274 314804 306280
rect 314856 306292 314976 306320
rect 315040 306292 315344 306320
rect 314476 306128 314528 306134
rect 314476 306070 314528 306076
rect 314660 306128 314712 306134
rect 314660 306070 314712 306076
rect 314660 304700 314712 304706
rect 314660 304642 314712 304648
rect 313832 300416 313884 300422
rect 313832 300358 313884 300364
rect 313648 299056 313700 299062
rect 313648 298998 313700 299004
rect 313556 287972 313608 287978
rect 313556 287914 313608 287920
rect 313464 282396 313516 282402
rect 313464 282338 313516 282344
rect 313372 265872 313424 265878
rect 313372 265814 313424 265820
rect 314672 261866 314700 304642
rect 314764 264450 314792 306274
rect 314856 271250 314884 306292
rect 314936 306196 314988 306202
rect 314936 306138 314988 306144
rect 314948 283830 314976 306138
rect 315040 294778 315068 306292
rect 315120 306128 315172 306134
rect 315120 306070 315172 306076
rect 315132 298994 315160 306070
rect 315408 305833 315436 310490
rect 315500 306338 315528 310420
rect 315488 306332 315540 306338
rect 315488 306274 315540 306280
rect 315394 305824 315450 305833
rect 315394 305759 315450 305768
rect 315684 304706 315712 310420
rect 315868 306202 315896 310420
rect 316052 306406 316080 310420
rect 316236 306610 316264 310420
rect 316224 306604 316276 306610
rect 316224 306546 316276 306552
rect 316420 306490 316448 310420
rect 316144 306462 316448 306490
rect 316040 306400 316092 306406
rect 316040 306342 316092 306348
rect 316144 306252 316172 306462
rect 316224 306400 316276 306406
rect 316224 306342 316276 306348
rect 316052 306224 316172 306252
rect 315856 306196 315908 306202
rect 315856 306138 315908 306144
rect 315672 304700 315724 304706
rect 315672 304642 315724 304648
rect 315120 298988 315172 298994
rect 315120 298930 315172 298936
rect 315028 294772 315080 294778
rect 315028 294714 315080 294720
rect 314936 283824 314988 283830
rect 314936 283766 314988 283772
rect 314844 271244 314896 271250
rect 314844 271186 314896 271192
rect 314752 264444 314804 264450
rect 314752 264386 314804 264392
rect 314660 261860 314712 261866
rect 314660 261802 314712 261808
rect 313278 254552 313334 254561
rect 313278 254487 313334 254496
rect 316052 253570 316080 306224
rect 316132 303544 316184 303550
rect 316132 303486 316184 303492
rect 316144 254794 316172 303486
rect 316236 260370 316264 306342
rect 316604 306320 316632 310420
rect 316328 306292 316632 306320
rect 316224 260364 316276 260370
rect 316224 260306 316276 260312
rect 316328 260302 316356 306292
rect 316408 306196 316460 306202
rect 316408 306138 316460 306144
rect 316420 261798 316448 306138
rect 316788 302234 316816 310420
rect 316868 306604 316920 306610
rect 316868 306546 316920 306552
rect 316512 302206 316816 302234
rect 316512 263090 316540 302206
rect 316880 296714 316908 306546
rect 316972 303550 317000 310420
rect 317156 306202 317184 310420
rect 317340 307834 317368 310420
rect 317538 310406 317736 310434
rect 317328 307828 317380 307834
rect 317328 307770 317380 307776
rect 317708 306610 317736 310406
rect 317800 307154 317828 310420
rect 317788 307148 317840 307154
rect 317788 307090 317840 307096
rect 317696 306604 317748 306610
rect 317696 306546 317748 306552
rect 317984 306490 318012 310420
rect 318064 307828 318116 307834
rect 318064 307770 318116 307776
rect 317524 306462 318012 306490
rect 317420 306264 317472 306270
rect 317420 306206 317472 306212
rect 317144 306196 317196 306202
rect 317144 306138 317196 306144
rect 316960 303544 317012 303550
rect 316960 303486 317012 303492
rect 316604 296686 316908 296714
rect 316604 263158 316632 296686
rect 317432 267306 317460 306206
rect 317524 275534 317552 306462
rect 317696 306400 317748 306406
rect 317696 306342 317748 306348
rect 317604 306332 317656 306338
rect 317604 306274 317656 306280
rect 317616 279614 317644 306274
rect 317708 290698 317736 306342
rect 317788 306196 317840 306202
rect 317788 306138 317840 306144
rect 317800 291922 317828 306138
rect 317788 291916 317840 291922
rect 317788 291858 317840 291864
rect 317696 290692 317748 290698
rect 317696 290634 317748 290640
rect 317604 279608 317656 279614
rect 317604 279550 317656 279556
rect 317512 275528 317564 275534
rect 317512 275470 317564 275476
rect 318076 270026 318104 307770
rect 318168 306202 318196 310420
rect 318248 306604 318300 306610
rect 318248 306546 318300 306552
rect 318156 306196 318208 306202
rect 318156 306138 318208 306144
rect 318260 303249 318288 306546
rect 318352 306338 318380 310420
rect 318340 306332 318392 306338
rect 318340 306274 318392 306280
rect 318536 306270 318564 310420
rect 318720 306406 318748 310420
rect 318708 306400 318760 306406
rect 318708 306342 318760 306348
rect 318800 306400 318852 306406
rect 318800 306342 318852 306348
rect 318524 306264 318576 306270
rect 318524 306206 318576 306212
rect 318246 303240 318302 303249
rect 318246 303175 318302 303184
rect 318064 270020 318116 270026
rect 318064 269962 318116 269968
rect 317420 267300 317472 267306
rect 317420 267242 317472 267248
rect 316592 263152 316644 263158
rect 316592 263094 316644 263100
rect 316500 263084 316552 263090
rect 316500 263026 316552 263032
rect 316408 261792 316460 261798
rect 316408 261734 316460 261740
rect 316316 260296 316368 260302
rect 316316 260238 316368 260244
rect 316132 254788 316184 254794
rect 316132 254730 316184 254736
rect 316040 253564 316092 253570
rect 316040 253506 316092 253512
rect 311900 250844 311952 250850
rect 311900 250786 311952 250792
rect 318812 249490 318840 306342
rect 318904 306320 318932 310420
rect 319088 306474 319116 310420
rect 319076 306468 319128 306474
rect 319076 306410 319128 306416
rect 319168 306332 319220 306338
rect 318904 306292 319116 306320
rect 318984 306196 319036 306202
rect 318984 306138 319036 306144
rect 318892 306128 318944 306134
rect 318892 306070 318944 306076
rect 318904 250714 318932 306070
rect 318996 256426 319024 306138
rect 319088 278186 319116 306292
rect 319168 306274 319220 306280
rect 319180 282334 319208 306274
rect 319272 297634 319300 310420
rect 319352 306468 319404 306474
rect 319352 306410 319404 306416
rect 319364 306105 319392 306410
rect 319456 306406 319484 310420
rect 319444 306400 319496 306406
rect 319444 306342 319496 306348
rect 319640 306202 319668 310420
rect 319824 306338 319852 310420
rect 319812 306332 319864 306338
rect 319812 306274 319864 306280
rect 319628 306196 319680 306202
rect 319628 306138 319680 306144
rect 320008 306134 320036 310420
rect 320180 306332 320232 306338
rect 320180 306274 320232 306280
rect 319996 306128 320048 306134
rect 319350 306096 319406 306105
rect 319996 306070 320048 306076
rect 319350 306031 319406 306040
rect 319260 297628 319312 297634
rect 319260 297570 319312 297576
rect 319168 282328 319220 282334
rect 319168 282270 319220 282276
rect 319076 278180 319128 278186
rect 319076 278122 319128 278128
rect 318984 256420 319036 256426
rect 318984 256362 319036 256368
rect 318892 250708 318944 250714
rect 318892 250650 318944 250656
rect 318800 249484 318852 249490
rect 318800 249426 318852 249432
rect 310610 248296 310666 248305
rect 310610 248231 310666 248240
rect 320192 247926 320220 306274
rect 320284 306134 320312 310420
rect 320364 306400 320416 306406
rect 320364 306342 320416 306348
rect 320272 306128 320324 306134
rect 320272 306070 320324 306076
rect 320272 305992 320324 305998
rect 320272 305934 320324 305940
rect 320284 256290 320312 305934
rect 320376 269958 320404 306342
rect 320468 306184 320496 310420
rect 320652 306406 320680 310420
rect 320640 306400 320692 306406
rect 320640 306342 320692 306348
rect 320468 306156 320588 306184
rect 320456 306060 320508 306066
rect 320456 306002 320508 306008
rect 320468 279546 320496 306002
rect 320560 280906 320588 306156
rect 320640 306128 320692 306134
rect 320640 306070 320692 306076
rect 320652 290630 320680 306070
rect 320836 296714 320864 310420
rect 321020 306066 321048 310420
rect 321204 306338 321232 310420
rect 321192 306332 321244 306338
rect 321192 306274 321244 306280
rect 321008 306060 321060 306066
rect 321008 306002 321060 306008
rect 321388 305998 321416 310420
rect 321572 306270 321600 310420
rect 321756 306354 321784 310420
rect 321836 307012 321888 307018
rect 321836 306954 321888 306960
rect 321848 306456 321876 306954
rect 321940 306524 321968 310420
rect 322124 307018 322152 310420
rect 322112 307012 322164 307018
rect 322112 306954 322164 306960
rect 321940 306496 322152 306524
rect 321848 306428 321968 306456
rect 321664 306326 321784 306354
rect 321836 306332 321888 306338
rect 321560 306264 321612 306270
rect 321560 306206 321612 306212
rect 321560 306128 321612 306134
rect 321560 306070 321612 306076
rect 321376 305992 321428 305998
rect 321376 305934 321428 305940
rect 320744 296686 320864 296714
rect 320744 296138 320772 296686
rect 320732 296132 320784 296138
rect 320732 296074 320784 296080
rect 320640 290624 320692 290630
rect 320640 290566 320692 290572
rect 320548 280900 320600 280906
rect 320548 280842 320600 280848
rect 320456 279540 320508 279546
rect 320456 279482 320508 279488
rect 320364 269952 320416 269958
rect 320364 269894 320416 269900
rect 320272 256284 320324 256290
rect 320272 256226 320324 256232
rect 321572 252074 321600 306070
rect 321664 252142 321692 306326
rect 321836 306274 321888 306280
rect 321744 306196 321796 306202
rect 321744 306138 321796 306144
rect 321756 256222 321784 306138
rect 321848 278118 321876 306274
rect 321940 289270 321968 306428
rect 322020 306264 322072 306270
rect 322020 306206 322072 306212
rect 322032 296206 322060 306206
rect 322124 299474 322152 306496
rect 322308 306134 322336 310420
rect 322492 306202 322520 310420
rect 322676 306338 322704 310420
rect 322952 306354 322980 310420
rect 323136 306490 323164 310420
rect 323320 306610 323348 310420
rect 323308 306604 323360 306610
rect 323308 306546 323360 306552
rect 323136 306462 323348 306490
rect 322664 306332 322716 306338
rect 322952 306326 323164 306354
rect 322664 306274 322716 306280
rect 322940 306264 322992 306270
rect 322940 306206 322992 306212
rect 322480 306196 322532 306202
rect 322480 306138 322532 306144
rect 322296 306128 322348 306134
rect 322296 306070 322348 306076
rect 322124 299446 322244 299474
rect 322216 297702 322244 299446
rect 322204 297696 322256 297702
rect 322204 297638 322256 297644
rect 322020 296200 322072 296206
rect 322020 296142 322072 296148
rect 321928 289264 321980 289270
rect 321928 289206 321980 289212
rect 321836 278112 321888 278118
rect 321836 278054 321888 278060
rect 321744 256216 321796 256222
rect 321744 256158 321796 256164
rect 322952 253434 322980 306206
rect 323032 306196 323084 306202
rect 323032 306138 323084 306144
rect 323044 256154 323072 306138
rect 323136 258874 323164 306326
rect 323216 306332 323268 306338
rect 323216 306274 323268 306280
rect 323228 261730 323256 306274
rect 323320 263022 323348 306462
rect 323504 306338 323532 310420
rect 323492 306332 323544 306338
rect 323492 306274 323544 306280
rect 323400 306264 323452 306270
rect 323400 306206 323452 306212
rect 323308 263016 323360 263022
rect 323308 262958 323360 262964
rect 323412 262954 323440 306206
rect 323688 302234 323716 310420
rect 323872 306202 323900 310420
rect 324056 306270 324084 310420
rect 324044 306264 324096 306270
rect 324044 306206 324096 306212
rect 323860 306196 323912 306202
rect 323860 306138 323912 306144
rect 323504 302206 323716 302234
rect 323504 264382 323532 302206
rect 324240 296714 324268 310420
rect 324424 306542 324452 310420
rect 324412 306536 324464 306542
rect 324412 306478 324464 306484
rect 324608 306354 324636 310420
rect 324792 306474 324820 310420
rect 324780 306468 324832 306474
rect 324780 306410 324832 306416
rect 324976 306354 325004 310420
rect 323596 296686 324268 296714
rect 324332 306326 324636 306354
rect 324700 306326 325004 306354
rect 323492 264376 323544 264382
rect 323492 264318 323544 264324
rect 323596 264314 323624 296686
rect 323584 264308 323636 264314
rect 323584 264250 323636 264256
rect 323400 262948 323452 262954
rect 323400 262890 323452 262896
rect 323216 261724 323268 261730
rect 323216 261666 323268 261672
rect 323124 258868 323176 258874
rect 323124 258810 323176 258816
rect 323032 256148 323084 256154
rect 323032 256090 323084 256096
rect 322940 253428 322992 253434
rect 322940 253370 322992 253376
rect 321652 252136 321704 252142
rect 321652 252078 321704 252084
rect 321560 252068 321612 252074
rect 321560 252010 321612 252016
rect 320180 247920 320232 247926
rect 320180 247862 320232 247868
rect 324332 245206 324360 306326
rect 324412 306264 324464 306270
rect 324412 306206 324464 306212
rect 324504 306264 324556 306270
rect 324504 306206 324556 306212
rect 324424 254726 324452 306206
rect 324516 262886 324544 306206
rect 324596 306196 324648 306202
rect 324596 306138 324648 306144
rect 324608 274174 324636 306138
rect 324700 275466 324728 306326
rect 325160 305130 325188 310420
rect 325344 310406 325450 310434
rect 325240 306536 325292 306542
rect 325240 306478 325292 306484
rect 324792 305102 325188 305130
rect 324792 276758 324820 305102
rect 325252 302234 325280 306478
rect 325344 306270 325372 310406
rect 325332 306264 325384 306270
rect 325332 306206 325384 306212
rect 325620 306202 325648 310420
rect 325804 306610 325832 310420
rect 325792 306604 325844 306610
rect 325792 306546 325844 306552
rect 325988 306490 326016 310420
rect 326172 309058 326200 310420
rect 326160 309052 326212 309058
rect 326160 308994 326212 309000
rect 325712 306462 326016 306490
rect 325608 306196 325660 306202
rect 325608 306138 325660 306144
rect 325068 302206 325280 302234
rect 325068 296714 325096 302206
rect 324884 296686 325096 296714
rect 324884 283762 324912 296686
rect 324872 283756 324924 283762
rect 324872 283698 324924 283704
rect 324780 276752 324832 276758
rect 324780 276694 324832 276700
rect 324688 275460 324740 275466
rect 324688 275402 324740 275408
rect 324596 274168 324648 274174
rect 324596 274110 324648 274116
rect 324504 262880 324556 262886
rect 324504 262822 324556 262828
rect 325712 256086 325740 306462
rect 325792 306400 325844 306406
rect 326356 306354 326384 310420
rect 326436 306604 326488 306610
rect 326436 306546 326488 306552
rect 325792 306342 325844 306348
rect 325804 274038 325832 306342
rect 325884 306332 325936 306338
rect 325884 306274 325936 306280
rect 325988 306326 326384 306354
rect 325896 276826 325924 306274
rect 325988 286482 326016 306326
rect 326448 304434 326476 306546
rect 326540 306338 326568 310420
rect 326528 306332 326580 306338
rect 326528 306274 326580 306280
rect 326436 304428 326488 304434
rect 326436 304370 326488 304376
rect 326724 302234 326752 310420
rect 326908 306406 326936 310420
rect 326896 306400 326948 306406
rect 326896 306342 326948 306348
rect 327092 306354 327120 310420
rect 327276 306490 327304 310420
rect 327276 306462 327396 306490
rect 327092 306326 327304 306354
rect 327080 306264 327132 306270
rect 327080 306206 327132 306212
rect 326080 302206 326752 302234
rect 326080 294710 326108 302206
rect 326068 294704 326120 294710
rect 326068 294646 326120 294652
rect 325976 286476 326028 286482
rect 325976 286418 326028 286424
rect 325884 276820 325936 276826
rect 325884 276762 325936 276768
rect 325792 274032 325844 274038
rect 325792 273974 325844 273980
rect 325700 256080 325752 256086
rect 325700 256022 325752 256028
rect 324412 254720 324464 254726
rect 324412 254662 324464 254668
rect 327092 249286 327120 306206
rect 327172 302864 327224 302870
rect 327172 302806 327224 302812
rect 327184 252006 327212 302806
rect 327276 274106 327304 306326
rect 327368 306218 327396 306462
rect 327460 306338 327488 310420
rect 327644 306490 327672 310420
rect 327644 306462 327764 306490
rect 327448 306332 327500 306338
rect 327448 306274 327500 306280
rect 327632 306332 327684 306338
rect 327632 306274 327684 306280
rect 327368 306190 327580 306218
rect 327356 305992 327408 305998
rect 327356 305934 327408 305940
rect 327368 282266 327396 305934
rect 327448 305924 327500 305930
rect 327448 305866 327500 305872
rect 327460 286414 327488 305866
rect 327552 287910 327580 306190
rect 327644 300286 327672 306274
rect 327736 305930 327764 306462
rect 327828 305998 327856 310420
rect 327920 310406 328118 310434
rect 327816 305992 327868 305998
rect 327816 305934 327868 305940
rect 327724 305924 327776 305930
rect 327724 305866 327776 305872
rect 327920 302870 327948 310406
rect 328288 306270 328316 310420
rect 328472 306610 328500 310420
rect 328656 306678 328684 310420
rect 328644 306672 328696 306678
rect 328644 306614 328696 306620
rect 328460 306604 328512 306610
rect 328460 306546 328512 306552
rect 328840 306490 328868 310420
rect 328920 306672 328972 306678
rect 328920 306614 328972 306620
rect 328472 306462 328868 306490
rect 328276 306264 328328 306270
rect 328276 306206 328328 306212
rect 327908 302864 327960 302870
rect 327908 302806 327960 302812
rect 327632 300280 327684 300286
rect 327632 300222 327684 300228
rect 327540 287904 327592 287910
rect 327540 287846 327592 287852
rect 327448 286408 327500 286414
rect 327448 286350 327500 286356
rect 327356 282260 327408 282266
rect 327356 282202 327408 282208
rect 327264 274100 327316 274106
rect 327264 274042 327316 274048
rect 327172 252000 327224 252006
rect 327172 251942 327224 251948
rect 327080 249280 327132 249286
rect 327080 249222 327132 249228
rect 328472 246702 328500 306462
rect 328552 306332 328604 306338
rect 328552 306274 328604 306280
rect 328564 249218 328592 306274
rect 328736 306264 328788 306270
rect 328736 306206 328788 306212
rect 328644 306128 328696 306134
rect 328644 306070 328696 306076
rect 328656 268462 328684 306070
rect 328644 268456 328696 268462
rect 328644 268398 328696 268404
rect 328748 268394 328776 306206
rect 328828 306196 328880 306202
rect 328828 306138 328880 306144
rect 328840 272542 328868 306138
rect 328932 275398 328960 306614
rect 329024 285054 329052 310420
rect 329104 306604 329156 306610
rect 329104 306546 329156 306552
rect 329116 293418 329144 306546
rect 329208 306134 329236 310420
rect 329392 306270 329420 310420
rect 329380 306264 329432 306270
rect 329380 306206 329432 306212
rect 329576 306202 329604 310420
rect 329760 306338 329788 310420
rect 329944 308417 329972 310420
rect 329930 308408 329986 308417
rect 329930 308343 329986 308352
rect 330128 306882 330156 310420
rect 330116 306876 330168 306882
rect 330116 306818 330168 306824
rect 330116 306672 330168 306678
rect 330116 306614 330168 306620
rect 329748 306332 329800 306338
rect 329748 306274 329800 306280
rect 329840 306332 329892 306338
rect 329840 306274 329892 306280
rect 329564 306196 329616 306202
rect 329564 306138 329616 306144
rect 329196 306128 329248 306134
rect 329196 306070 329248 306076
rect 329104 293412 329156 293418
rect 329104 293354 329156 293360
rect 329012 285048 329064 285054
rect 329012 284990 329064 284996
rect 328920 275392 328972 275398
rect 328920 275334 328972 275340
rect 328828 272536 328880 272542
rect 328828 272478 328880 272484
rect 328736 268388 328788 268394
rect 328736 268330 328788 268336
rect 328552 249212 328604 249218
rect 328552 249154 328604 249160
rect 328460 246696 328512 246702
rect 328460 246638 328512 246644
rect 324320 245200 324372 245206
rect 324320 245142 324372 245148
rect 329852 245070 329880 306274
rect 330024 306264 330076 306270
rect 330024 306206 330076 306212
rect 329932 302660 329984 302666
rect 329932 302602 329984 302608
rect 329944 245138 329972 302602
rect 330036 246498 330064 306206
rect 330128 246634 330156 306614
rect 330312 302666 330340 310420
rect 330404 310406 330602 310434
rect 330404 306338 330432 310406
rect 330392 306332 330444 306338
rect 330392 306274 330444 306280
rect 330300 302660 330352 302666
rect 330300 302602 330352 302608
rect 330772 302234 330800 310420
rect 330220 302206 330800 302234
rect 330116 246628 330168 246634
rect 330116 246570 330168 246576
rect 330220 246566 330248 302206
rect 330956 296714 330984 310420
rect 331140 306270 331168 310420
rect 331220 308372 331272 308378
rect 331220 308314 331272 308320
rect 331128 306264 331180 306270
rect 331128 306206 331180 306212
rect 330312 296686 330984 296714
rect 330312 250646 330340 296686
rect 330300 250640 330352 250646
rect 330300 250582 330352 250588
rect 330208 246560 330260 246566
rect 330208 246502 330260 246508
rect 330024 246492 330076 246498
rect 330024 246434 330076 246440
rect 331232 246430 331260 308314
rect 331324 308310 331352 310420
rect 331508 308394 331536 310420
rect 331692 308530 331720 310420
rect 331416 308366 331536 308394
rect 331600 308502 331720 308530
rect 331312 308304 331364 308310
rect 331312 308246 331364 308252
rect 331312 308168 331364 308174
rect 331312 308110 331364 308116
rect 331324 265810 331352 308110
rect 331416 269890 331444 308366
rect 331600 308258 331628 308502
rect 331876 308394 331904 310420
rect 331508 308230 331628 308258
rect 331692 308366 331904 308394
rect 331508 289202 331536 308230
rect 331588 307692 331640 307698
rect 331588 307634 331640 307640
rect 331600 301578 331628 307634
rect 331692 303113 331720 308366
rect 331772 308304 331824 308310
rect 331772 308246 331824 308252
rect 331784 304366 331812 308246
rect 332060 308174 332088 310420
rect 332244 308378 332272 310420
rect 332232 308372 332284 308378
rect 332232 308314 332284 308320
rect 332048 308168 332100 308174
rect 332048 308110 332100 308116
rect 332428 307698 332456 310420
rect 332612 308394 332640 310420
rect 332796 308666 332824 310420
rect 332994 310406 333192 310434
rect 332796 308638 333008 308666
rect 332520 308366 332640 308394
rect 332520 308174 332548 308366
rect 332692 308304 332744 308310
rect 332980 308258 333008 308638
rect 333060 308372 333112 308378
rect 333060 308314 333112 308320
rect 332692 308246 332744 308252
rect 332600 308236 332652 308242
rect 332600 308178 332652 308184
rect 332508 308168 332560 308174
rect 332508 308110 332560 308116
rect 332416 307692 332468 307698
rect 332416 307634 332468 307640
rect 331772 304360 331824 304366
rect 331772 304302 331824 304308
rect 331678 303104 331734 303113
rect 331678 303039 331734 303048
rect 331588 301572 331640 301578
rect 331588 301514 331640 301520
rect 331496 289196 331548 289202
rect 331496 289138 331548 289144
rect 331404 269884 331456 269890
rect 331404 269826 331456 269832
rect 331312 265804 331364 265810
rect 331312 265746 331364 265752
rect 332612 247858 332640 308178
rect 332704 253298 332732 308246
rect 332796 308230 333008 308258
rect 332796 253366 332824 308230
rect 332876 308168 332928 308174
rect 332876 308110 332928 308116
rect 332888 267170 332916 308110
rect 332968 307352 333020 307358
rect 332968 307294 333020 307300
rect 332980 279478 333008 307294
rect 333072 298926 333100 308314
rect 333164 300218 333192 310406
rect 333256 307358 333284 310420
rect 333440 308310 333468 310420
rect 333624 308378 333652 310420
rect 333612 308372 333664 308378
rect 333612 308314 333664 308320
rect 333428 308304 333480 308310
rect 333428 308246 333480 308252
rect 333808 308242 333836 310420
rect 333992 308990 334020 310420
rect 333980 308984 334032 308990
rect 333980 308926 334032 308932
rect 334176 308394 334204 310420
rect 334256 308984 334308 308990
rect 334256 308926 334308 308932
rect 333992 308366 334204 308394
rect 333796 308236 333848 308242
rect 333796 308178 333848 308184
rect 333244 307352 333296 307358
rect 333244 307294 333296 307300
rect 333152 300212 333204 300218
rect 333152 300154 333204 300160
rect 333060 298920 333112 298926
rect 333060 298862 333112 298868
rect 332968 279472 333020 279478
rect 332968 279414 333020 279420
rect 332876 267164 332928 267170
rect 332876 267106 332928 267112
rect 332784 253360 332836 253366
rect 332784 253302 332836 253308
rect 332692 253292 332744 253298
rect 332692 253234 332744 253240
rect 332600 247852 332652 247858
rect 332600 247794 332652 247800
rect 333992 247790 334020 308366
rect 334072 308236 334124 308242
rect 334072 308178 334124 308184
rect 333980 247784 334032 247790
rect 333980 247726 334032 247732
rect 334084 247722 334112 308178
rect 334164 308168 334216 308174
rect 334164 308110 334216 308116
rect 334176 249150 334204 308110
rect 334268 250578 334296 308926
rect 334360 256018 334388 310420
rect 334544 308394 334572 310420
rect 334440 308372 334492 308378
rect 334544 308366 334664 308394
rect 334440 308314 334492 308320
rect 334452 257514 334480 308314
rect 334532 308304 334584 308310
rect 334532 308246 334584 308252
rect 334544 261594 334572 308246
rect 334636 261662 334664 308366
rect 334728 308242 334756 310420
rect 334912 308378 334940 310420
rect 334900 308372 334952 308378
rect 334900 308314 334952 308320
rect 335096 308310 335124 310420
rect 335084 308304 335136 308310
rect 335084 308246 335136 308252
rect 334716 308236 334768 308242
rect 334716 308178 334768 308184
rect 335280 308174 335308 310420
rect 335478 310406 335676 310434
rect 335544 308304 335596 308310
rect 335544 308246 335596 308252
rect 335360 308236 335412 308242
rect 335360 308178 335412 308184
rect 335268 308168 335320 308174
rect 335268 308110 335320 308116
rect 334624 261656 334676 261662
rect 334624 261598 334676 261604
rect 334532 261588 334584 261594
rect 334532 261530 334584 261536
rect 334440 257508 334492 257514
rect 334440 257450 334492 257456
rect 334348 256012 334400 256018
rect 334348 255954 334400 255960
rect 334256 250572 334308 250578
rect 334256 250514 334308 250520
rect 334164 249144 334216 249150
rect 334164 249086 334216 249092
rect 334072 247716 334124 247722
rect 334072 247658 334124 247664
rect 331220 246424 331272 246430
rect 331220 246366 331272 246372
rect 335372 246362 335400 308178
rect 335452 308168 335504 308174
rect 335452 308110 335504 308116
rect 335464 249082 335492 308110
rect 335556 271182 335584 308246
rect 335648 276690 335676 310406
rect 335740 293350 335768 310420
rect 335820 308372 335872 308378
rect 335820 308314 335872 308320
rect 335832 296070 335860 308314
rect 335924 304298 335952 310420
rect 336108 308242 336136 310420
rect 336292 308310 336320 310420
rect 336476 308378 336504 310420
rect 336464 308372 336516 308378
rect 336464 308314 336516 308320
rect 336280 308304 336332 308310
rect 336280 308246 336332 308252
rect 336096 308236 336148 308242
rect 336096 308178 336148 308184
rect 336660 308174 336688 310420
rect 336740 308984 336792 308990
rect 336740 308926 336792 308932
rect 336648 308168 336700 308174
rect 336648 308110 336700 308116
rect 335912 304292 335964 304298
rect 335912 304234 335964 304240
rect 335820 296064 335872 296070
rect 335820 296006 335872 296012
rect 335728 293344 335780 293350
rect 335728 293286 335780 293292
rect 335636 276684 335688 276690
rect 335636 276626 335688 276632
rect 335544 271176 335596 271182
rect 335544 271118 335596 271124
rect 335452 249076 335504 249082
rect 335452 249018 335504 249024
rect 336752 247625 336780 308926
rect 336844 308310 336872 310420
rect 337028 308530 337056 310420
rect 336936 308502 337056 308530
rect 336832 308304 336884 308310
rect 336832 308246 336884 308252
rect 336936 308174 336964 308502
rect 337212 308394 337240 310420
rect 337396 308990 337424 310420
rect 337384 308984 337436 308990
rect 337384 308926 337436 308932
rect 337028 308366 337240 308394
rect 336924 308168 336976 308174
rect 336924 308110 336976 308116
rect 336924 307896 336976 307902
rect 336924 307838 336976 307844
rect 336832 307828 336884 307834
rect 336832 307770 336884 307776
rect 336844 253230 336872 307770
rect 336936 275330 336964 307838
rect 337028 283694 337056 308366
rect 337108 308304 337160 308310
rect 337580 308292 337608 310420
rect 337108 308246 337160 308252
rect 337212 308264 337608 308292
rect 337120 287774 337148 308246
rect 337212 294642 337240 308264
rect 337292 308168 337344 308174
rect 337292 308110 337344 308116
rect 337304 302977 337332 308110
rect 337764 307902 337792 310420
rect 337752 307896 337804 307902
rect 337752 307838 337804 307844
rect 337948 307834 337976 310420
rect 338146 310406 338252 310434
rect 338224 308310 338252 310406
rect 338316 310406 338422 310434
rect 338212 308304 338264 308310
rect 338212 308246 338264 308252
rect 338120 308236 338172 308242
rect 338120 308178 338172 308184
rect 337936 307828 337988 307834
rect 337936 307770 337988 307776
rect 337290 302968 337346 302977
rect 337290 302903 337346 302912
rect 337200 294636 337252 294642
rect 337200 294578 337252 294584
rect 337108 287768 337160 287774
rect 337108 287710 337160 287716
rect 337016 283688 337068 283694
rect 337016 283630 337068 283636
rect 336924 275324 336976 275330
rect 336924 275266 336976 275272
rect 336832 253224 336884 253230
rect 336832 253166 336884 253172
rect 336738 247616 336794 247625
rect 336738 247551 336794 247560
rect 335360 246356 335412 246362
rect 335360 246298 335412 246304
rect 329932 245132 329984 245138
rect 329932 245074 329984 245080
rect 329840 245064 329892 245070
rect 329840 245006 329892 245012
rect 338132 245002 338160 308178
rect 338212 308168 338264 308174
rect 338212 308110 338264 308116
rect 338224 265742 338252 308110
rect 338316 273970 338344 310406
rect 338592 308530 338620 310420
rect 338408 308502 338620 308530
rect 338408 283626 338436 308502
rect 338776 308394 338804 310420
rect 338488 308372 338540 308378
rect 338488 308314 338540 308320
rect 338592 308366 338804 308394
rect 338500 291854 338528 308314
rect 338592 293282 338620 308366
rect 338672 308304 338724 308310
rect 338672 308246 338724 308252
rect 338684 301510 338712 308246
rect 338960 308242 338988 310420
rect 338948 308236 339000 308242
rect 338948 308178 339000 308184
rect 339144 308174 339172 310420
rect 339328 308378 339356 310420
rect 339316 308372 339368 308378
rect 339316 308314 339368 308320
rect 339132 308168 339184 308174
rect 339132 308110 339184 308116
rect 338672 301504 338724 301510
rect 338672 301446 338724 301452
rect 338580 293276 338632 293282
rect 338580 293218 338632 293224
rect 338488 291848 338540 291854
rect 338488 291790 338540 291796
rect 338396 283620 338448 283626
rect 338396 283562 338448 283568
rect 338304 273964 338356 273970
rect 338304 273906 338356 273912
rect 338212 265736 338264 265742
rect 338212 265678 338264 265684
rect 339512 251938 339540 310420
rect 339696 308394 339724 310420
rect 339880 308394 339908 310420
rect 339696 308366 339816 308394
rect 339880 308366 340000 308394
rect 339684 308236 339736 308242
rect 339684 308178 339736 308184
rect 339592 307284 339644 307290
rect 339592 307226 339644 307232
rect 339604 257378 339632 307226
rect 339696 257446 339724 308178
rect 339788 258738 339816 308366
rect 339868 308304 339920 308310
rect 339868 308246 339920 308252
rect 339880 260234 339908 308246
rect 339972 300150 340000 308366
rect 340064 308242 340092 310420
rect 340144 309052 340196 309058
rect 340144 308994 340196 309000
rect 340052 308236 340104 308242
rect 340052 308178 340104 308184
rect 339960 300144 340012 300150
rect 339960 300086 340012 300092
rect 339868 260228 339920 260234
rect 339868 260170 339920 260176
rect 339776 258732 339828 258738
rect 339776 258674 339828 258680
rect 339684 257440 339736 257446
rect 339684 257382 339736 257388
rect 339592 257372 339644 257378
rect 339592 257314 339644 257320
rect 339500 251932 339552 251938
rect 339500 251874 339552 251880
rect 340156 249422 340184 308994
rect 340248 308310 340276 310420
rect 340236 308304 340288 308310
rect 340236 308246 340288 308252
rect 340432 307086 340460 310420
rect 340616 307290 340644 310420
rect 340604 307284 340656 307290
rect 340604 307226 340656 307232
rect 340420 307080 340472 307086
rect 340420 307022 340472 307028
rect 340892 306542 340920 310420
rect 340880 306536 340932 306542
rect 340880 306478 340932 306484
rect 340880 306400 340932 306406
rect 340880 306342 340932 306348
rect 340892 267102 340920 306342
rect 340972 306264 341024 306270
rect 340972 306206 341024 306212
rect 340984 269822 341012 306206
rect 341076 306134 341104 310420
rect 341260 306354 341288 310420
rect 341444 306406 341472 310420
rect 341432 306400 341484 306406
rect 341156 306332 341208 306338
rect 341260 306326 341380 306354
rect 341432 306342 341484 306348
rect 341156 306274 341208 306280
rect 341064 306128 341116 306134
rect 341064 306070 341116 306076
rect 341064 305992 341116 305998
rect 341064 305934 341116 305940
rect 341076 278050 341104 305934
rect 341168 289134 341196 306274
rect 341248 306196 341300 306202
rect 341248 306138 341300 306144
rect 341260 290494 341288 306138
rect 341352 290562 341380 306326
rect 341628 306202 341656 310420
rect 341708 306536 341760 306542
rect 341708 306478 341760 306484
rect 341616 306196 341668 306202
rect 341616 306138 341668 306144
rect 341432 306128 341484 306134
rect 341432 306070 341484 306076
rect 341444 298858 341472 306070
rect 341720 302841 341748 306478
rect 341812 306270 341840 310420
rect 341800 306264 341852 306270
rect 341800 306206 341852 306212
rect 341996 305998 342024 310420
rect 342180 306338 342208 310420
rect 342364 306354 342392 310420
rect 342548 306626 342576 310420
rect 342732 306746 342760 310420
rect 342720 306740 342772 306746
rect 342720 306682 342772 306688
rect 342548 306598 342852 306626
rect 342720 306468 342772 306474
rect 342720 306410 342772 306416
rect 342168 306332 342220 306338
rect 342364 306326 342576 306354
rect 342168 306274 342220 306280
rect 342352 306264 342404 306270
rect 342352 306206 342404 306212
rect 341984 305992 342036 305998
rect 341984 305934 342036 305940
rect 342260 305788 342312 305794
rect 342260 305730 342312 305736
rect 341706 302832 341762 302841
rect 341706 302767 341762 302776
rect 341432 298852 341484 298858
rect 341432 298794 341484 298800
rect 341340 290556 341392 290562
rect 341340 290498 341392 290504
rect 341248 290488 341300 290494
rect 341248 290430 341300 290436
rect 341156 289128 341208 289134
rect 341156 289070 341208 289076
rect 341064 278044 341116 278050
rect 341064 277986 341116 277992
rect 340972 269816 341024 269822
rect 340972 269758 341024 269764
rect 340880 267096 340932 267102
rect 340880 267038 340932 267044
rect 340144 249416 340196 249422
rect 340144 249358 340196 249364
rect 338120 244996 338172 245002
rect 338120 244938 338172 244944
rect 342272 244934 342300 305730
rect 342364 260166 342392 306206
rect 342444 303748 342496 303754
rect 342444 303690 342496 303696
rect 342456 265674 342484 303690
rect 342548 282198 342576 306326
rect 342628 306332 342680 306338
rect 342628 306274 342680 306280
rect 342640 287706 342668 306274
rect 342732 297430 342760 306410
rect 342824 297498 342852 306598
rect 342916 306270 342944 310420
rect 342904 306264 342956 306270
rect 342904 306206 342956 306212
rect 343100 305794 343128 310420
rect 343284 306338 343312 310420
rect 343376 310406 343574 310434
rect 343272 306332 343324 306338
rect 343272 306274 343324 306280
rect 343088 305788 343140 305794
rect 343088 305730 343140 305736
rect 343376 303754 343404 310406
rect 343744 306354 343772 310420
rect 343652 306326 343772 306354
rect 343824 306332 343876 306338
rect 343364 303748 343416 303754
rect 343364 303690 343416 303696
rect 342812 297492 342864 297498
rect 342812 297434 342864 297440
rect 342720 297424 342772 297430
rect 342720 297366 342772 297372
rect 342628 287700 342680 287706
rect 342628 287642 342680 287648
rect 342536 282192 342588 282198
rect 342536 282134 342588 282140
rect 342444 265668 342496 265674
rect 342444 265610 342496 265616
rect 342352 260160 342404 260166
rect 342352 260102 342404 260108
rect 343652 254658 343680 306326
rect 343824 306274 343876 306280
rect 343732 306264 343784 306270
rect 343732 306206 343784 306212
rect 343640 254652 343692 254658
rect 343640 254594 343692 254600
rect 343744 254590 343772 306206
rect 343836 261526 343864 306274
rect 343928 306066 343956 310420
rect 344112 309134 344140 310420
rect 344020 309106 344140 309134
rect 343916 306060 343968 306066
rect 343916 306002 343968 306008
rect 344020 304042 344048 309106
rect 344296 306270 344324 310420
rect 344284 306264 344336 306270
rect 344284 306206 344336 306212
rect 344100 305856 344152 305862
rect 344100 305798 344152 305804
rect 343928 304014 344048 304042
rect 343928 267034 343956 304014
rect 344008 303612 344060 303618
rect 344008 303554 344060 303560
rect 344020 286346 344048 303554
rect 344112 296002 344140 305798
rect 344480 303618 344508 310420
rect 344664 306338 344692 310420
rect 344652 306332 344704 306338
rect 344652 306274 344704 306280
rect 344468 303612 344520 303618
rect 344468 303554 344520 303560
rect 344848 298790 344876 310420
rect 345032 306490 345060 310420
rect 345032 306462 345152 306490
rect 345020 306332 345072 306338
rect 345020 306274 345072 306280
rect 344836 298784 344888 298790
rect 344836 298726 344888 298732
rect 344100 295996 344152 296002
rect 344100 295938 344152 295944
rect 344008 286340 344060 286346
rect 344008 286282 344060 286288
rect 343916 267028 343968 267034
rect 343916 266970 343968 266976
rect 343824 261520 343876 261526
rect 343824 261462 343876 261468
rect 343732 254584 343784 254590
rect 343732 254526 343784 254532
rect 345032 250510 345060 306274
rect 345124 305697 345152 306462
rect 345216 306270 345244 310420
rect 345400 306354 345428 310420
rect 345308 306326 345428 306354
rect 345204 306264 345256 306270
rect 345204 306206 345256 306212
rect 345204 306128 345256 306134
rect 345204 306070 345256 306076
rect 345110 305688 345166 305697
rect 345110 305623 345166 305632
rect 345112 302388 345164 302394
rect 345112 302330 345164 302336
rect 345124 251870 345152 302330
rect 345216 254862 345244 306070
rect 345308 264246 345336 306326
rect 345388 306264 345440 306270
rect 345388 306206 345440 306212
rect 345400 280838 345428 306206
rect 345584 302234 345612 310420
rect 345768 306338 345796 310420
rect 345860 310406 346058 310434
rect 345756 306332 345808 306338
rect 345756 306274 345808 306280
rect 345860 302394 345888 310406
rect 346228 306134 346256 310420
rect 346216 306128 346268 306134
rect 346216 306070 346268 306076
rect 345848 302388 345900 302394
rect 345848 302330 345900 302336
rect 345492 302206 345612 302234
rect 345492 284986 345520 302206
rect 345480 284980 345532 284986
rect 345480 284922 345532 284928
rect 345388 280832 345440 280838
rect 345388 280774 345440 280780
rect 345296 264240 345348 264246
rect 345296 264182 345348 264188
rect 345204 254856 345256 254862
rect 345204 254798 345256 254804
rect 345112 251864 345164 251870
rect 345112 251806 345164 251812
rect 345020 250504 345072 250510
rect 345020 250446 345072 250452
rect 346412 249354 346440 310420
rect 346596 306354 346624 310420
rect 346780 308281 346808 310420
rect 346964 309097 346992 310420
rect 346950 309088 347006 309097
rect 346950 309023 347006 309032
rect 346766 308272 346822 308281
rect 346766 308207 346822 308216
rect 346504 306326 346624 306354
rect 346504 258806 346532 306326
rect 347148 305726 347176 310420
rect 347136 305720 347188 305726
rect 347136 305662 347188 305668
rect 347332 302234 347360 310420
rect 347516 308961 347544 310420
rect 347700 309126 347728 310420
rect 347688 309120 347740 309126
rect 347688 309062 347740 309068
rect 347502 308952 347558 308961
rect 347502 308887 347558 308896
rect 347884 306490 347912 310420
rect 347884 306462 348004 306490
rect 347780 306400 347832 306406
rect 347780 306342 347832 306348
rect 346596 302206 347360 302234
rect 346596 297566 346624 302206
rect 346584 297560 346636 297566
rect 346584 297502 346636 297508
rect 346492 258800 346544 258806
rect 346492 258742 346544 258748
rect 347792 253502 347820 306342
rect 347872 306332 347924 306338
rect 347872 306274 347924 306280
rect 347884 300082 347912 306274
rect 347976 303142 348004 306462
rect 347964 303136 348016 303142
rect 347964 303078 348016 303084
rect 348068 302234 348096 310420
rect 348252 306338 348280 310420
rect 348436 308825 348464 310420
rect 348422 308816 348478 308825
rect 348422 308751 348478 308760
rect 348424 307828 348476 307834
rect 348424 307770 348476 307776
rect 348240 306332 348292 306338
rect 348240 306274 348292 306280
rect 347976 302206 348096 302234
rect 347976 301646 348004 302206
rect 347964 301640 348016 301646
rect 347964 301582 348016 301588
rect 347872 300076 347924 300082
rect 347872 300018 347924 300024
rect 348436 256358 348464 307770
rect 348712 303346 348740 310420
rect 348700 303340 348752 303346
rect 348700 303282 348752 303288
rect 348896 303074 348924 310420
rect 348976 309052 349028 309058
rect 348976 308994 349028 309000
rect 348884 303068 348936 303074
rect 348884 303010 348936 303016
rect 348988 299946 349016 308994
rect 349080 306406 349108 310420
rect 349264 308689 349292 310420
rect 349250 308680 349306 308689
rect 349250 308615 349306 308624
rect 349068 306400 349120 306406
rect 349068 306342 349120 306348
rect 349448 302870 349476 310420
rect 349632 303210 349660 310420
rect 349620 303204 349672 303210
rect 349620 303146 349672 303152
rect 349436 302864 349488 302870
rect 349436 302806 349488 302812
rect 349816 301714 349844 310420
rect 350000 306241 350028 310420
rect 349986 306232 350042 306241
rect 349986 306167 350042 306176
rect 350184 302734 350212 310420
rect 350368 307834 350396 310420
rect 350552 308310 350580 310420
rect 350632 308984 350684 308990
rect 350632 308926 350684 308932
rect 350540 308304 350592 308310
rect 350540 308246 350592 308252
rect 350356 307828 350408 307834
rect 350356 307770 350408 307776
rect 350644 303278 350672 308926
rect 350736 303550 350764 310420
rect 350920 309058 350948 310420
rect 351012 310406 351210 310434
rect 350908 309052 350960 309058
rect 350908 308994 350960 309000
rect 351012 308394 351040 310406
rect 351380 308990 351408 310420
rect 351368 308984 351420 308990
rect 351368 308926 351420 308932
rect 351564 308394 351592 310420
rect 350828 308366 351040 308394
rect 351104 308366 351592 308394
rect 350828 305862 350856 308366
rect 351000 308304 351052 308310
rect 351000 308246 351052 308252
rect 350908 308236 350960 308242
rect 350908 308178 350960 308184
rect 350816 305856 350868 305862
rect 350816 305798 350868 305804
rect 350920 305454 350948 308178
rect 351012 306377 351040 308246
rect 350998 306368 351054 306377
rect 350998 306303 351054 306312
rect 350908 305448 350960 305454
rect 350908 305390 350960 305396
rect 350724 303544 350776 303550
rect 350724 303486 350776 303492
rect 350632 303272 350684 303278
rect 350632 303214 350684 303220
rect 350172 302728 350224 302734
rect 350172 302670 350224 302676
rect 349804 301708 349856 301714
rect 349804 301650 349856 301656
rect 348976 299940 349028 299946
rect 348976 299882 349028 299888
rect 351104 267238 351132 308366
rect 351184 308304 351236 308310
rect 351184 308246 351236 308252
rect 351196 287842 351224 308246
rect 351748 308242 351776 310420
rect 351736 308236 351788 308242
rect 351736 308178 351788 308184
rect 351932 308038 351960 310420
rect 352116 308530 352144 310420
rect 352024 308502 352144 308530
rect 352024 308310 352052 308502
rect 352104 308372 352156 308378
rect 352104 308314 352156 308320
rect 352012 308304 352064 308310
rect 352012 308246 352064 308252
rect 352012 308168 352064 308174
rect 352012 308110 352064 308116
rect 351920 308032 351972 308038
rect 351920 307974 351972 307980
rect 352024 303482 352052 308110
rect 352012 303476 352064 303482
rect 352012 303418 352064 303424
rect 352116 303414 352144 308314
rect 352196 308304 352248 308310
rect 352196 308246 352248 308252
rect 352208 306202 352236 308246
rect 352196 306196 352248 306202
rect 352196 306138 352248 306144
rect 352300 305930 352328 310420
rect 352484 308378 352512 310420
rect 352472 308372 352524 308378
rect 352472 308314 352524 308320
rect 352668 308310 352696 310420
rect 352656 308304 352708 308310
rect 352656 308246 352708 308252
rect 352852 308242 352880 310420
rect 353036 308242 353064 310420
rect 352840 308236 352892 308242
rect 352840 308178 352892 308184
rect 353024 308236 353076 308242
rect 353024 308178 353076 308184
rect 353220 308122 353248 310420
rect 353404 308530 353432 310420
rect 353404 308502 353524 308530
rect 353392 308372 353444 308378
rect 353392 308314 353444 308320
rect 353300 308304 353352 308310
rect 353300 308246 353352 308252
rect 352392 308094 353248 308122
rect 352392 306270 352420 308094
rect 352564 308032 352616 308038
rect 352564 307974 352616 307980
rect 352380 306264 352432 306270
rect 352380 306206 352432 306212
rect 352288 305924 352340 305930
rect 352288 305866 352340 305872
rect 352104 303408 352156 303414
rect 352104 303350 352156 303356
rect 352576 302802 352604 307974
rect 353312 305658 353340 308246
rect 353404 305794 353432 308314
rect 353496 308038 353524 308502
rect 353484 308032 353536 308038
rect 353484 307974 353536 307980
rect 353392 305788 353444 305794
rect 353392 305730 353444 305736
rect 353300 305652 353352 305658
rect 353300 305594 353352 305600
rect 353588 305590 353616 310420
rect 353864 308242 353892 310420
rect 354048 308378 354076 310420
rect 354232 309126 354260 310420
rect 354220 309120 354272 309126
rect 354220 309062 354272 309068
rect 354036 308372 354088 308378
rect 354036 308314 354088 308320
rect 354416 308310 354444 310420
rect 354600 309058 354628 310420
rect 354588 309052 354640 309058
rect 354588 308994 354640 309000
rect 354680 308440 354732 308446
rect 354680 308382 354732 308388
rect 354404 308304 354456 308310
rect 354404 308246 354456 308252
rect 353852 308236 353904 308242
rect 353852 308178 353904 308184
rect 354692 308106 354720 308382
rect 354680 308100 354732 308106
rect 354680 308042 354732 308048
rect 354784 307714 354812 310420
rect 354864 308440 354916 308446
rect 354864 308382 354916 308388
rect 354692 307686 354812 307714
rect 354692 305998 354720 307686
rect 354772 307624 354824 307630
rect 354772 307566 354824 307572
rect 354784 306134 354812 307566
rect 354876 306338 354904 308382
rect 354968 307902 354996 310420
rect 355048 308576 355100 308582
rect 355048 308518 355100 308524
rect 354956 307896 355008 307902
rect 354956 307838 355008 307844
rect 354956 307760 355008 307766
rect 354956 307702 355008 307708
rect 354864 306332 354916 306338
rect 354864 306274 354916 306280
rect 354772 306128 354824 306134
rect 354772 306070 354824 306076
rect 354968 306066 354996 307702
rect 355060 307170 355088 308518
rect 355152 307766 355180 310420
rect 355336 308922 355364 310420
rect 355232 308916 355284 308922
rect 355232 308858 355284 308864
rect 355324 308916 355376 308922
rect 355324 308858 355376 308864
rect 355140 307760 355192 307766
rect 355140 307702 355192 307708
rect 355244 307306 355272 308858
rect 355416 308712 355468 308718
rect 355416 308654 355468 308660
rect 355428 307442 355456 308654
rect 355520 307630 355548 310420
rect 355704 308802 355732 310420
rect 355600 308780 355652 308786
rect 355704 308774 355824 308802
rect 355600 308722 355652 308728
rect 355508 307624 355560 307630
rect 355508 307566 355560 307572
rect 355428 307414 355548 307442
rect 355244 307278 355456 307306
rect 355060 307142 355272 307170
rect 355244 306374 355272 307142
rect 355244 306346 355364 306374
rect 354956 306060 355008 306066
rect 354956 306002 355008 306008
rect 354680 305992 354732 305998
rect 354680 305934 354732 305940
rect 353576 305584 353628 305590
rect 353576 305526 353628 305532
rect 352564 302796 352616 302802
rect 352564 302738 352616 302744
rect 351184 287836 351236 287842
rect 351184 287778 351236 287784
rect 351092 267232 351144 267238
rect 351092 267174 351144 267180
rect 348424 256352 348476 256358
rect 348424 256294 348476 256300
rect 347780 253496 347832 253502
rect 347780 253438 347832 253444
rect 346400 249348 346452 249354
rect 346400 249290 346452 249296
rect 342260 244928 342312 244934
rect 342260 244870 342312 244876
rect 355336 244866 355364 306346
rect 355428 245614 355456 307278
rect 355416 245608 355468 245614
rect 355416 245550 355468 245556
rect 355324 244860 355376 244866
rect 355324 244802 355376 244808
rect 310518 244760 310574 244769
rect 310518 244695 310574 244704
rect 355520 244662 355548 307414
rect 355612 244798 355640 308722
rect 355692 308644 355744 308650
rect 355692 308586 355744 308592
rect 355704 247518 355732 308586
rect 355796 308174 355824 308774
rect 355888 308446 355916 310420
rect 356072 308786 356100 310420
rect 356164 310406 356362 310434
rect 356060 308780 356112 308786
rect 356060 308722 356112 308728
rect 355876 308440 355928 308446
rect 355876 308382 355928 308388
rect 355784 308168 355836 308174
rect 355784 308110 355836 308116
rect 356060 306876 356112 306882
rect 356060 306818 356112 306824
rect 356072 303618 356100 306818
rect 356164 305522 356192 310406
rect 356532 308718 356560 310420
rect 356520 308712 356572 308718
rect 356520 308654 356572 308660
rect 356716 307970 356744 310420
rect 356900 308938 356928 310420
rect 356900 308910 357020 308938
rect 356888 308848 356940 308854
rect 356888 308790 356940 308796
rect 356796 308508 356848 308514
rect 356796 308450 356848 308456
rect 356704 307964 356756 307970
rect 356704 307906 356756 307912
rect 356152 305516 356204 305522
rect 356152 305458 356204 305464
rect 356060 303612 356112 303618
rect 356060 303554 356112 303560
rect 356704 247580 356756 247586
rect 356704 247522 356756 247528
rect 355692 247512 355744 247518
rect 355692 247454 355744 247460
rect 355600 244792 355652 244798
rect 355600 244734 355652 244740
rect 355508 244656 355560 244662
rect 355508 244598 355560 244604
rect 303618 243672 303674 243681
rect 300952 243636 301004 243642
rect 303618 243607 303674 243616
rect 300952 243578 301004 243584
rect 299572 243568 299624 243574
rect 297272 243510 297324 243516
rect 298650 243536 298706 243545
rect 299572 243510 299624 243516
rect 298650 243471 298706 243480
rect 258538 159896 258594 159905
rect 258538 159831 258594 159840
rect 275834 159896 275890 159905
rect 275834 159831 275890 159840
rect 277030 159896 277086 159905
rect 277030 159831 277086 159840
rect 278134 159896 278190 159905
rect 278134 159831 278190 159840
rect 279238 159896 279294 159905
rect 279238 159831 279294 159840
rect 256700 159656 256752 159662
rect 255962 159624 256018 159633
rect 256700 159598 256752 159604
rect 255962 159559 256018 159568
rect 239588 158772 239640 158778
rect 239588 158714 239640 158720
rect 238116 158704 238168 158710
rect 220818 158672 220874 158681
rect 238114 158672 238116 158681
rect 239600 158681 239628 158714
rect 238168 158672 238170 158681
rect 220818 158607 220874 158616
rect 230480 158636 230532 158642
rect 219438 158264 219494 158273
rect 219438 158199 219494 158208
rect 219452 16574 219480 158199
rect 220832 16574 220860 158607
rect 238114 158607 238170 158616
rect 239586 158672 239642 158681
rect 239586 158607 239642 158616
rect 240690 158672 240746 158681
rect 240690 158607 240746 158616
rect 248326 158672 248382 158681
rect 248326 158607 248382 158616
rect 250166 158672 250222 158681
rect 250166 158607 250222 158616
rect 230480 158578 230532 158584
rect 224958 158536 225014 158545
rect 224958 158471 225014 158480
rect 223578 157856 223634 157865
rect 223578 157791 223634 157800
rect 219452 16546 220032 16574
rect 220832 16546 221136 16574
rect 219348 3936 219400 3942
rect 219348 3878 219400 3884
rect 218060 3528 218112 3534
rect 216862 3496 216918 3505
rect 216588 3460 216640 3466
rect 218060 3470 218112 3476
rect 219164 3528 219216 3534
rect 219164 3470 219216 3476
rect 219254 3496 219310 3505
rect 216862 3431 216918 3440
rect 216588 3402 216640 3408
rect 216496 3188 216548 3194
rect 216496 3130 216548 3136
rect 216876 480 216904 3431
rect 218072 480 218100 3470
rect 219254 3431 219310 3440
rect 219268 480 219296 3431
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 16546
rect 222750 3360 222806 3369
rect 222750 3295 222806 3304
rect 222764 480 222792 3295
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 157791
rect 224972 16574 225000 158471
rect 227718 158400 227774 158409
rect 227718 158335 227774 158344
rect 227732 16574 227760 158335
rect 229100 157820 229152 157826
rect 229100 157762 229152 157768
rect 229112 16574 229140 157762
rect 230492 16574 230520 158578
rect 236000 158568 236052 158574
rect 236000 158510 236052 158516
rect 234712 158500 234764 158506
rect 234712 158442 234764 158448
rect 231858 158128 231914 158137
rect 231858 158063 231914 158072
rect 224972 16546 225184 16574
rect 227732 16546 228312 16574
rect 229112 16546 229416 16574
rect 230492 16546 231072 16574
rect 225156 480 225184 16546
rect 226340 3324 226392 3330
rect 226340 3266 226392 3272
rect 226352 480 226380 3266
rect 227536 3188 227588 3194
rect 227536 3130 227588 3136
rect 227548 480 227576 3130
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 16546
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 16546
rect 231044 480 231072 16546
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 231872 354 231900 158063
rect 233240 157956 233292 157962
rect 233240 157898 233292 157904
rect 233252 16574 233280 157898
rect 234620 157888 234672 157894
rect 234620 157830 234672 157836
rect 233252 16546 233464 16574
rect 233436 480 233464 16546
rect 234632 11762 234660 157830
rect 234620 11756 234672 11762
rect 234620 11698 234672 11704
rect 234724 6914 234752 158442
rect 236012 16574 236040 158510
rect 238758 157992 238814 158001
rect 238758 157927 238814 157936
rect 237380 155848 237432 155854
rect 237380 155790 237432 155796
rect 237392 16574 237420 155790
rect 238772 16574 238800 157927
rect 240704 157758 240732 158607
rect 242992 158432 243044 158438
rect 242992 158374 243044 158380
rect 242900 158364 242952 158370
rect 242900 158306 242952 158312
rect 240692 157752 240744 157758
rect 240692 157694 240744 157700
rect 241520 155780 241572 155786
rect 241520 155722 241572 155728
rect 241532 16574 241560 155722
rect 236012 16546 236592 16574
rect 237392 16546 237696 16574
rect 238772 16546 239352 16574
rect 241532 16546 241744 16574
rect 235816 11756 235868 11762
rect 235816 11698 235868 11704
rect 234632 6886 234752 6914
rect 234632 480 234660 6886
rect 235828 480 235856 11698
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 16546
rect 239324 480 239352 16546
rect 240508 3392 240560 3398
rect 240508 3334 240560 3340
rect 240520 480 240548 3334
rect 241716 480 241744 16546
rect 242912 11762 242940 158306
rect 242900 11756 242952 11762
rect 242900 11698 242952 11704
rect 243004 6914 243032 158374
rect 245660 158296 245712 158302
rect 245382 158264 245438 158273
rect 245660 158238 245712 158244
rect 245382 158199 245438 158208
rect 245396 155922 245424 158199
rect 245384 155916 245436 155922
rect 245384 155858 245436 155864
rect 245672 16574 245700 158238
rect 247040 158228 247092 158234
rect 247040 158170 247092 158176
rect 246854 158128 246910 158137
rect 246854 158063 246910 158072
rect 246868 155961 246896 158063
rect 246854 155952 246910 155961
rect 246854 155887 246910 155896
rect 247052 16574 247080 158170
rect 248340 157282 248368 158607
rect 249800 158092 249852 158098
rect 249800 158034 249852 158040
rect 248694 157992 248750 158001
rect 248694 157927 248750 157936
rect 248328 157276 248380 157282
rect 248328 157218 248380 157224
rect 248708 155825 248736 157927
rect 248694 155816 248750 155825
rect 248694 155751 248750 155760
rect 248420 155712 248472 155718
rect 248420 155654 248472 155660
rect 245672 16546 245976 16574
rect 247052 16546 247632 16574
rect 244096 11756 244148 11762
rect 244096 11698 244148 11704
rect 242912 6886 243032 6914
rect 242912 480 242940 6886
rect 244108 480 244136 11698
rect 245200 4140 245252 4146
rect 245200 4082 245252 4088
rect 245212 480 245240 4082
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 16546
rect 247604 480 247632 16546
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248432 354 248460 155654
rect 249812 16574 249840 158034
rect 250180 157350 250208 158607
rect 252374 158536 252430 158545
rect 252374 158471 252430 158480
rect 251180 158160 251232 158166
rect 251180 158102 251232 158108
rect 250168 157344 250220 157350
rect 250168 157286 250220 157292
rect 249812 16546 250024 16574
rect 249996 480 250024 16546
rect 251192 480 251220 158102
rect 252098 157992 252154 158001
rect 252098 157927 252154 157936
rect 252112 155786 252140 157927
rect 252388 156777 252416 158471
rect 252560 158024 252612 158030
rect 252560 157966 252612 157972
rect 253570 157992 253626 158001
rect 252374 156768 252430 156777
rect 252374 156703 252430 156712
rect 252100 155780 252152 155786
rect 252100 155722 252152 155728
rect 251270 155408 251326 155417
rect 251270 155343 251326 155352
rect 251284 16574 251312 155343
rect 252572 16574 252600 157966
rect 253570 157927 253626 157936
rect 253202 157312 253258 157321
rect 253202 157247 253258 157256
rect 253216 156913 253244 157247
rect 253202 156904 253258 156913
rect 253202 156839 253258 156848
rect 253584 155854 253612 157927
rect 253662 157448 253718 157457
rect 253662 157383 253718 157392
rect 253572 155848 253624 155854
rect 253572 155790 253624 155796
rect 253676 154562 253704 157383
rect 255976 157146 256004 159559
rect 256606 158672 256662 158681
rect 256606 158607 256662 158616
rect 256620 157690 256648 158607
rect 256608 157684 256660 157690
rect 256608 157626 256660 157632
rect 255964 157140 256016 157146
rect 255964 157082 256016 157088
rect 253940 155576 253992 155582
rect 253940 155518 253992 155524
rect 253664 154556 253716 154562
rect 253664 154498 253716 154504
rect 253952 16574 253980 155518
rect 255320 155440 255372 155446
rect 255320 155382 255372 155388
rect 255332 16574 255360 155382
rect 251284 16546 252416 16574
rect 252572 16546 253520 16574
rect 253952 16546 254256 16574
rect 255332 16546 255912 16574
rect 252388 480 252416 16546
rect 253492 480 253520 16546
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 16546
rect 255884 480 255912 16546
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 256712 354 256740 159598
rect 258552 158778 258580 159831
rect 271050 159624 271106 159633
rect 260840 159588 260892 159594
rect 271050 159559 271106 159568
rect 274454 159624 274510 159633
rect 274454 159559 274510 159568
rect 260840 159530 260892 159536
rect 259460 159452 259512 159458
rect 259460 159394 259512 159400
rect 258540 158772 258592 158778
rect 258540 158714 258592 158720
rect 257158 158672 257214 158681
rect 257158 158607 257214 158616
rect 258630 158672 258686 158681
rect 258630 158607 258686 158616
rect 257172 157214 257200 158607
rect 257160 157208 257212 157214
rect 257160 157150 257212 157156
rect 258644 157078 258672 158607
rect 258632 157072 258684 157078
rect 258632 157014 258684 157020
rect 259472 151814 259500 159394
rect 259550 158672 259606 158681
rect 259550 158607 259606 158616
rect 259564 158574 259592 158607
rect 259552 158568 259604 158574
rect 259552 158510 259604 158516
rect 260654 158536 260710 158545
rect 260654 158471 260710 158480
rect 260668 157010 260696 158471
rect 260656 157004 260708 157010
rect 260656 156946 260708 156952
rect 259472 151786 259592 151814
rect 259564 6914 259592 151786
rect 260852 16574 260880 159530
rect 264980 159520 265032 159526
rect 264980 159462 265032 159468
rect 262864 158840 262916 158846
rect 262864 158782 262916 158788
rect 262876 158681 262904 158782
rect 261758 158672 261814 158681
rect 261758 158607 261814 158616
rect 262862 158672 262918 158681
rect 262862 158607 262918 158616
rect 261772 157418 261800 158607
rect 261942 157992 261998 158001
rect 261942 157927 261998 157936
rect 261760 157412 261812 157418
rect 261760 157354 261812 157360
rect 261956 155718 261984 157927
rect 264426 157720 264482 157729
rect 264426 157655 264482 157664
rect 263966 157448 264022 157457
rect 263966 157383 264022 157392
rect 261944 155712 261996 155718
rect 261944 155654 261996 155660
rect 263600 155372 263652 155378
rect 263600 155314 263652 155320
rect 263612 16574 263640 155314
rect 263980 154494 264008 157383
rect 264440 155378 264468 157655
rect 264428 155372 264480 155378
rect 264428 155314 264480 155320
rect 263968 154488 264020 154494
rect 263968 154430 264020 154436
rect 260852 16546 261800 16574
rect 263612 16546 264192 16574
rect 259472 6886 259592 6914
rect 258264 4072 258316 4078
rect 258264 4014 258316 4020
rect 258276 480 258304 4014
rect 259472 480 259500 6886
rect 260656 4004 260708 4010
rect 260656 3946 260708 3952
rect 260668 480 260696 3946
rect 261772 480 261800 16546
rect 262956 3868 263008 3874
rect 262956 3810 263008 3816
rect 262968 480 262996 3810
rect 264164 480 264192 16546
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 264992 354 265020 159462
rect 267648 158908 267700 158914
rect 267648 158850 267700 158856
rect 267660 158681 267688 158850
rect 265990 158672 266046 158681
rect 265990 158607 266046 158616
rect 267646 158672 267702 158681
rect 267646 158607 267702 158616
rect 268750 158672 268806 158681
rect 268750 158607 268806 158616
rect 270222 158672 270278 158681
rect 270222 158607 270278 158616
rect 266004 158506 266032 158607
rect 265992 158500 266044 158506
rect 265992 158442 266044 158448
rect 268764 158438 268792 158607
rect 268752 158432 268804 158438
rect 268752 158374 268804 158380
rect 270236 158370 270264 158607
rect 270224 158364 270276 158370
rect 270224 158306 270276 158312
rect 266726 157992 266782 158001
rect 266726 157927 266782 157936
rect 268934 157992 268990 158001
rect 268934 157927 268990 157936
rect 265990 157720 266046 157729
rect 265990 157655 266046 157664
rect 266004 155446 266032 157655
rect 266740 155582 266768 157927
rect 268948 155650 268976 157927
rect 267832 155644 267884 155650
rect 267832 155586 267884 155592
rect 268936 155644 268988 155650
rect 268936 155586 268988 155592
rect 266728 155576 266780 155582
rect 266728 155518 266780 155524
rect 265992 155440 266044 155446
rect 265992 155382 266044 155388
rect 267844 6914 267872 155586
rect 271064 155514 271092 159559
rect 274468 158982 274496 159559
rect 275848 159118 275876 159831
rect 275836 159112 275888 159118
rect 275836 159054 275888 159060
rect 277044 159050 277072 159831
rect 278148 159186 278176 159831
rect 279252 159254 279280 159831
rect 300950 159760 301006 159769
rect 300950 159695 301006 159704
rect 282920 159384 282972 159390
rect 282920 159326 282972 159332
rect 296718 159352 296774 159361
rect 279240 159248 279292 159254
rect 279240 159190 279292 159196
rect 278136 159180 278188 159186
rect 278136 159122 278188 159128
rect 277032 159044 277084 159050
rect 277032 158986 277084 158992
rect 274456 158976 274508 158982
rect 274456 158918 274508 158924
rect 271142 158672 271198 158681
rect 271142 158607 271198 158616
rect 272246 158672 272302 158681
rect 272246 158607 272302 158616
rect 271156 158302 271184 158607
rect 271144 158296 271196 158302
rect 271144 158238 271196 158244
rect 272260 157894 272288 158607
rect 276110 158536 276166 158545
rect 276110 158471 276166 158480
rect 281354 158536 281410 158545
rect 281354 158471 281410 158480
rect 273350 158400 273406 158409
rect 273350 158335 273406 158344
rect 272248 157888 272300 157894
rect 272248 157830 272300 157836
rect 273364 156738 273392 158335
rect 274454 157720 274510 157729
rect 274454 157655 274510 157664
rect 273352 156732 273404 156738
rect 273352 156674 273404 156680
rect 270500 155508 270552 155514
rect 270500 155450 270552 155456
rect 271052 155508 271104 155514
rect 271052 155450 271104 155456
rect 269118 155272 269174 155281
rect 269118 155207 269174 155216
rect 269132 16574 269160 155207
rect 270512 16574 270540 155450
rect 274468 155310 274496 157655
rect 276124 156942 276152 158471
rect 278686 157720 278742 157729
rect 278686 157655 278742 157664
rect 276112 156936 276164 156942
rect 276112 156878 276164 156884
rect 273260 155304 273312 155310
rect 273260 155246 273312 155252
rect 274456 155304 274508 155310
rect 274456 155246 274508 155252
rect 269132 16546 270080 16574
rect 270512 16546 270816 16574
rect 267752 6886 267872 6914
rect 266544 3936 266596 3942
rect 266544 3878 266596 3884
rect 266556 480 266584 3878
rect 267752 480 267780 6886
rect 268844 3732 268896 3738
rect 268844 3674 268896 3680
rect 268856 480 268884 3674
rect 270052 480 270080 16546
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 270788 354 270816 16546
rect 272432 3596 272484 3602
rect 272432 3538 272484 3544
rect 272444 480 272472 3538
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273272 354 273300 155246
rect 278700 155242 278728 157655
rect 281368 156874 281396 158471
rect 281356 156868 281408 156874
rect 281356 156810 281408 156816
rect 274640 155236 274692 155242
rect 274640 155178 274692 155184
rect 278688 155236 278740 155242
rect 278688 155178 278740 155184
rect 274652 16574 274680 155178
rect 278780 155168 278832 155174
rect 278780 155110 278832 155116
rect 277400 155032 277452 155038
rect 277400 154974 277452 154980
rect 277412 16574 277440 154974
rect 278792 16574 278820 155110
rect 282932 16574 282960 159326
rect 300964 159322 300992 159695
rect 322940 159588 322992 159594
rect 322940 159530 322992 159536
rect 320088 159520 320140 159526
rect 320088 159462 320140 159468
rect 314660 159452 314712 159458
rect 314660 159394 314712 159400
rect 310428 159384 310480 159390
rect 310428 159326 310480 159332
rect 296718 159287 296774 159296
rect 300952 159316 301004 159322
rect 286230 158536 286286 158545
rect 286230 158471 286286 158480
rect 284114 157720 284170 157729
rect 284114 157655 284170 157664
rect 284128 155174 284156 157655
rect 286244 156806 286272 158471
rect 291014 158400 291070 158409
rect 291014 158335 291070 158344
rect 296258 158400 296314 158409
rect 296258 158335 296314 158344
rect 288254 157584 288310 157593
rect 288254 157519 288310 157528
rect 286232 156800 286284 156806
rect 286232 156742 286284 156748
rect 284116 155168 284168 155174
rect 284116 155110 284168 155116
rect 288268 155106 288296 157519
rect 291028 156670 291056 158335
rect 293590 157584 293646 157593
rect 293590 157519 293646 157528
rect 291016 156664 291068 156670
rect 291016 156606 291068 156612
rect 292578 155408 292634 155417
rect 292578 155343 292634 155352
rect 291198 155272 291254 155281
rect 291198 155207 291254 155216
rect 287060 155100 287112 155106
rect 287060 155042 287112 155048
rect 288256 155100 288308 155106
rect 288256 155042 288308 155048
rect 287072 16574 287100 155042
rect 288440 153876 288492 153882
rect 288440 153818 288492 153824
rect 288452 16574 288480 153818
rect 291212 16574 291240 155207
rect 292592 16574 292620 155343
rect 293604 155038 293632 157519
rect 296272 156602 296300 158335
rect 296260 156596 296312 156602
rect 296260 156538 296312 156544
rect 293958 155544 294014 155553
rect 293958 155479 294014 155488
rect 293592 155032 293644 155038
rect 293592 154974 293644 154980
rect 293972 16574 294000 155479
rect 295340 153944 295392 153950
rect 295340 153886 295392 153892
rect 295352 16574 295380 153886
rect 296732 16574 296760 159287
rect 300952 159258 301004 159264
rect 308680 158704 308732 158710
rect 298926 158672 298982 158681
rect 298926 158607 298982 158616
rect 303526 158672 303582 158681
rect 303526 158607 303582 158616
rect 306102 158672 306158 158681
rect 306102 158607 306104 158616
rect 298940 158234 298968 158607
rect 298928 158228 298980 158234
rect 298928 158170 298980 158176
rect 303540 158166 303568 158607
rect 306156 158607 306158 158616
rect 308678 158672 308680 158681
rect 308732 158672 308734 158681
rect 308678 158607 308734 158616
rect 306104 158578 306156 158584
rect 310440 158166 310468 159326
rect 313462 158672 313518 158681
rect 314672 158642 314700 159394
rect 320100 158710 320128 159462
rect 320088 158704 320140 158710
rect 315854 158672 315910 158681
rect 313462 158607 313518 158616
rect 314660 158636 314712 158642
rect 311254 158264 311310 158273
rect 311254 158199 311310 158208
rect 303528 158160 303580 158166
rect 303528 158102 303580 158108
rect 310428 158160 310480 158166
rect 310428 158102 310480 158108
rect 311268 156466 311296 158199
rect 313476 158098 313504 158607
rect 315854 158607 315910 158616
rect 318614 158672 318670 158681
rect 320088 158646 320140 158652
rect 321190 158672 321246 158681
rect 318614 158607 318670 158616
rect 321190 158607 321246 158616
rect 314660 158578 314712 158584
rect 313464 158092 313516 158098
rect 313464 158034 313516 158040
rect 315868 158030 315896 158607
rect 315856 158024 315908 158030
rect 315856 157966 315908 157972
rect 318628 157962 318656 158607
rect 321204 158166 321232 158607
rect 321192 158160 321244 158166
rect 321192 158102 321244 158108
rect 318616 157956 318668 157962
rect 318616 157898 318668 157904
rect 322952 157894 322980 159530
rect 323398 158672 323454 158681
rect 323398 158607 323454 158616
rect 325974 158672 326030 158681
rect 325974 158607 326030 158616
rect 323412 157894 323440 158607
rect 322940 157888 322992 157894
rect 322940 157830 322992 157836
rect 323400 157888 323452 157894
rect 323400 157830 323452 157836
rect 325988 157826 326016 158607
rect 353942 158536 353998 158545
rect 353942 158471 353998 158480
rect 348422 158264 348478 158273
rect 348422 158199 348478 158208
rect 345662 157992 345718 158001
rect 345662 157927 345718 157936
rect 325976 157820 326028 157826
rect 325976 157762 326028 157768
rect 317052 157412 317104 157418
rect 317052 157354 317104 157360
rect 317064 156534 317092 157354
rect 317052 156528 317104 156534
rect 317052 156470 317104 156476
rect 311256 156460 311308 156466
rect 311256 156402 311308 156408
rect 299480 154012 299532 154018
rect 299480 153954 299532 153960
rect 299492 16574 299520 153954
rect 300860 152516 300912 152522
rect 300860 152458 300912 152464
rect 300872 16574 300900 152458
rect 274652 16546 274864 16574
rect 277412 16546 278360 16574
rect 278792 16546 279096 16574
rect 282932 16546 283144 16574
rect 287072 16546 287376 16574
rect 288452 16546 289032 16574
rect 291212 16546 291424 16574
rect 292592 16546 293264 16574
rect 293972 16546 294920 16574
rect 295352 16546 295656 16574
rect 296732 16546 297312 16574
rect 299492 16546 299704 16574
rect 300872 16546 301544 16574
rect 274836 480 274864 16546
rect 277124 3800 277176 3806
rect 277124 3742 277176 3748
rect 276020 3664 276072 3670
rect 276020 3606 276072 3612
rect 276032 480 276060 3606
rect 277136 480 277164 3742
rect 278332 480 278360 16546
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 280712 3528 280764 3534
rect 280712 3470 280764 3476
rect 281908 3528 281960 3534
rect 281908 3470 281960 3476
rect 280724 480 280752 3470
rect 281920 480 281948 3470
rect 283116 480 283144 16546
rect 285404 3596 285456 3602
rect 285404 3538 285456 3544
rect 284300 3460 284352 3466
rect 284300 3402 284352 3408
rect 284312 480 284340 3402
rect 285416 480 285444 3538
rect 286600 3460 286652 3466
rect 286600 3402 286652 3408
rect 286612 480 286640 3402
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 289004 480 289032 16546
rect 290188 3664 290240 3670
rect 290188 3606 290240 3612
rect 290200 480 290228 3606
rect 291396 480 291424 16546
rect 292580 3732 292632 3738
rect 292580 3674 292632 3680
rect 292592 480 292620 3674
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 294892 480 294920 16546
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 295628 354 295656 16546
rect 297284 480 297312 16546
rect 298468 3868 298520 3874
rect 298468 3810 298520 3816
rect 298480 480 298508 3810
rect 299676 480 299704 16546
rect 300768 3800 300820 3806
rect 300768 3742 300820 3748
rect 300780 480 300808 3742
rect 296046 354 296158 480
rect 295628 326 296158 354
rect 296046 -960 296158 326
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 16546
rect 316224 9308 316276 9314
rect 316224 9250 316276 9256
rect 312636 9172 312688 9178
rect 312636 9114 312688 9120
rect 305552 9104 305604 9110
rect 305552 9046 305604 9052
rect 303160 9036 303212 9042
rect 303160 8978 303212 8984
rect 303172 480 303200 8978
rect 304356 8968 304408 8974
rect 304356 8910 304408 8916
rect 304368 480 304396 8910
rect 305564 480 305592 9046
rect 311440 6452 311492 6458
rect 311440 6394 311492 6400
rect 310244 6384 310296 6390
rect 310244 6326 310296 6332
rect 307944 6316 307996 6322
rect 307944 6258 307996 6264
rect 306748 6248 306800 6254
rect 306748 6190 306800 6196
rect 306760 480 306788 6190
rect 307956 480 307984 6258
rect 309048 6180 309100 6186
rect 309048 6122 309100 6128
rect 309060 480 309088 6122
rect 310256 480 310284 6326
rect 311452 480 311480 6394
rect 312648 480 312676 9114
rect 315028 6724 315080 6730
rect 315028 6666 315080 6672
rect 313832 6656 313884 6662
rect 313832 6598 313884 6604
rect 313844 480 313872 6598
rect 315040 480 315068 6666
rect 316236 480 316264 9250
rect 319720 9240 319772 9246
rect 319720 9182 319772 9188
rect 318524 6588 318576 6594
rect 318524 6530 318576 6536
rect 317328 6520 317380 6526
rect 317328 6462 317380 6468
rect 317340 480 317368 6462
rect 318536 480 318564 6530
rect 319732 480 319760 9182
rect 330392 6860 330444 6866
rect 330392 6802 330444 6808
rect 326804 6792 326856 6798
rect 326804 6734 326856 6740
rect 323306 6352 323362 6361
rect 323306 6287 323362 6296
rect 320914 6216 320970 6225
rect 320914 6151 320970 6160
rect 320928 480 320956 6151
rect 322112 3936 322164 3942
rect 322112 3878 322164 3884
rect 322124 480 322152 3878
rect 323320 480 323348 6287
rect 325606 3496 325662 3505
rect 325606 3431 325662 3440
rect 324410 3360 324466 3369
rect 324410 3295 324466 3304
rect 324424 480 324452 3295
rect 325620 480 325648 3431
rect 326816 480 326844 6734
rect 329196 4004 329248 4010
rect 329196 3946 329248 3952
rect 327998 3632 328054 3641
rect 327998 3567 328054 3576
rect 328012 480 328040 3567
rect 329208 480 329236 3946
rect 330404 480 330432 6802
rect 344558 6488 344614 6497
rect 344558 6423 344614 6432
rect 333888 6112 333940 6118
rect 333888 6054 333940 6060
rect 332692 4072 332744 4078
rect 332692 4014 332744 4020
rect 331586 3768 331642 3777
rect 331586 3703 331642 3712
rect 331600 480 331628 3703
rect 332704 480 332732 4014
rect 333900 480 333928 6054
rect 337476 6044 337528 6050
rect 337476 5986 337528 5992
rect 336280 4140 336332 4146
rect 336280 4082 336332 4088
rect 335082 3904 335138 3913
rect 335082 3839 335138 3848
rect 335096 480 335124 3839
rect 336292 480 336320 4082
rect 337488 480 337516 5986
rect 340972 5976 341024 5982
rect 340972 5918 341024 5924
rect 339868 3392 339920 3398
rect 339868 3334 339920 3340
rect 338672 3324 338724 3330
rect 338672 3266 338724 3272
rect 338684 480 338712 3266
rect 339880 480 339908 3334
rect 340984 480 341012 5918
rect 343362 4040 343418 4049
rect 343362 3975 343418 3984
rect 342168 3256 342220 3262
rect 342168 3198 342220 3204
rect 342180 480 342208 3198
rect 343376 480 343404 3975
rect 344572 480 344600 6423
rect 345676 3602 345704 157927
rect 345756 152584 345808 152590
rect 345756 152526 345808 152532
rect 345768 3874 345796 152526
rect 348054 6624 348110 6633
rect 348054 6559 348110 6568
rect 345756 3868 345808 3874
rect 345756 3810 345808 3816
rect 345664 3596 345716 3602
rect 345664 3538 345716 3544
rect 346950 3224 347006 3233
rect 345756 3188 345808 3194
rect 346950 3159 347006 3168
rect 345756 3130 345808 3136
rect 345768 480 345796 3130
rect 346964 480 346992 3159
rect 348068 480 348096 6559
rect 348436 3738 348464 158199
rect 351182 158128 351238 158137
rect 351182 158063 351238 158072
rect 350446 6896 350502 6905
rect 350446 6831 350502 6840
rect 348424 3732 348476 3738
rect 348424 3674 348476 3680
rect 349252 3596 349304 3602
rect 349252 3538 349304 3544
rect 349264 480 349292 3538
rect 350460 480 350488 6831
rect 351196 3670 351224 158063
rect 351642 6760 351698 6769
rect 351642 6695 351698 6704
rect 351184 3664 351236 3670
rect 351184 3606 351236 3612
rect 351656 480 351684 6695
rect 352840 3732 352892 3738
rect 352840 3674 352892 3680
rect 352852 480 352880 3674
rect 353956 3534 353984 158471
rect 354126 158400 354182 158409
rect 354126 158335 354182 158344
rect 354140 3806 354168 158335
rect 356426 4040 356482 4049
rect 356426 3975 356482 3984
rect 356610 4040 356666 4049
rect 356610 3975 356666 3984
rect 354128 3800 354180 3806
rect 354128 3742 354180 3748
rect 355140 3800 355192 3806
rect 355140 3742 355192 3748
rect 354036 3664 354088 3670
rect 354036 3606 354088 3612
rect 353944 3528 353996 3534
rect 353944 3470 353996 3476
rect 354048 480 354076 3606
rect 355152 3602 355180 3742
rect 355140 3596 355192 3602
rect 355140 3538 355192 3544
rect 355232 3596 355284 3602
rect 355232 3538 355284 3544
rect 355244 480 355272 3538
rect 356336 3528 356388 3534
rect 356336 3470 356388 3476
rect 356348 480 356376 3470
rect 356440 2961 356468 3975
rect 356624 3777 356652 3975
rect 356716 3942 356744 247522
rect 356808 242214 356836 308450
rect 356900 243545 356928 308790
rect 356992 308650 357020 308910
rect 356980 308644 357032 308650
rect 356980 308586 357032 308592
rect 356980 308100 357032 308106
rect 356980 308042 357032 308048
rect 356992 243982 357020 308042
rect 357084 306882 357112 310420
rect 357268 308582 357296 310420
rect 357256 308576 357308 308582
rect 357452 308530 357480 310420
rect 357256 308518 357308 308524
rect 357360 308502 357480 308530
rect 357360 308242 357388 308502
rect 357636 308292 357664 310420
rect 357820 308394 357848 310420
rect 357452 308264 357664 308292
rect 357728 308366 357848 308394
rect 357348 308236 357400 308242
rect 357348 308178 357400 308184
rect 357072 306876 357124 306882
rect 357072 306818 357124 306824
rect 356980 243976 357032 243982
rect 356980 243918 357032 243924
rect 356886 243536 356942 243545
rect 356886 243471 356942 243480
rect 356796 242208 356848 242214
rect 356796 242150 356848 242156
rect 357346 159488 357402 159497
rect 357346 159423 357402 159432
rect 357360 158817 357388 159423
rect 357346 158808 357402 158817
rect 357346 158743 357402 158752
rect 357452 158438 357480 308264
rect 357624 308100 357676 308106
rect 357624 308042 357676 308048
rect 357532 306876 357584 306882
rect 357532 306818 357584 306824
rect 357440 158432 357492 158438
rect 357440 158374 357492 158380
rect 357544 158302 357572 306818
rect 357636 158370 357664 308042
rect 357728 159390 357756 308366
rect 357808 308236 357860 308242
rect 357808 308178 357860 308184
rect 357716 159384 357768 159390
rect 357716 159326 357768 159332
rect 357820 159322 357848 308178
rect 358004 308106 358032 310420
rect 357992 308100 358044 308106
rect 357992 308042 358044 308048
rect 358188 307986 358216 310420
rect 357912 307958 358216 307986
rect 357912 159458 357940 307958
rect 358372 306882 358400 310420
rect 358360 306876 358412 306882
rect 358360 306818 358412 306824
rect 358556 306762 358584 310420
rect 358004 306734 358584 306762
rect 358004 159526 358032 306734
rect 358740 306374 358768 310420
rect 358924 310406 359030 310434
rect 358820 308848 358872 308854
rect 358820 308790 358872 308796
rect 358096 306346 358768 306374
rect 358096 159594 358124 306346
rect 358266 305960 358322 305969
rect 358266 305895 358322 305904
rect 358176 244656 358228 244662
rect 358176 244598 358228 244604
rect 358084 159588 358136 159594
rect 358084 159530 358136 159536
rect 357992 159520 358044 159526
rect 357992 159462 358044 159468
rect 357900 159452 357952 159458
rect 357900 159394 357952 159400
rect 357808 159316 357860 159322
rect 357808 159258 357860 159264
rect 358082 158808 358138 158817
rect 358082 158743 358138 158752
rect 357624 158364 357676 158370
rect 357624 158306 357676 158312
rect 357532 158296 357584 158302
rect 357532 158238 357584 158244
rect 356704 3936 356756 3942
rect 356704 3878 356756 3884
rect 356610 3768 356666 3777
rect 356610 3703 356666 3712
rect 356702 3632 356758 3641
rect 356702 3567 356758 3576
rect 357530 3632 357586 3641
rect 357530 3567 357586 3576
rect 356716 3233 356744 3567
rect 356702 3224 356758 3233
rect 356702 3159 356758 3168
rect 356426 2952 356482 2961
rect 356426 2887 356482 2896
rect 357544 480 357572 3567
rect 358096 3534 358124 158743
rect 358188 6390 358216 244598
rect 358280 158545 358308 305895
rect 358266 158536 358322 158545
rect 358266 158471 358322 158480
rect 358832 156738 358860 308790
rect 358820 156732 358872 156738
rect 358820 156674 358872 156680
rect 358924 156466 358952 310406
rect 359200 308854 359228 310420
rect 359188 308848 359240 308854
rect 359188 308790 359240 308796
rect 359384 308530 359412 310420
rect 359016 308502 359412 308530
rect 359016 158098 359044 308502
rect 359280 308440 359332 308446
rect 359568 308394 359596 310420
rect 359280 308382 359332 308388
rect 359096 308236 359148 308242
rect 359096 308178 359148 308184
rect 359004 158092 359056 158098
rect 359004 158034 359056 158040
rect 359108 158030 359136 308178
rect 359188 308168 359240 308174
rect 359188 308110 359240 308116
rect 359096 158024 359148 158030
rect 359096 157966 359148 157972
rect 359200 157962 359228 308110
rect 359292 159118 359320 308382
rect 359384 308366 359596 308394
rect 359280 159112 359332 159118
rect 359280 159054 359332 159060
rect 359384 158982 359412 308366
rect 359752 308242 359780 310420
rect 359936 308446 359964 310420
rect 359924 308440 359976 308446
rect 359924 308382 359976 308388
rect 359740 308236 359792 308242
rect 359740 308178 359792 308184
rect 360120 308174 360148 310420
rect 360108 308168 360160 308174
rect 360108 308110 360160 308116
rect 359556 307964 359608 307970
rect 359556 307906 359608 307912
rect 359464 248328 359516 248334
rect 359464 248270 359516 248276
rect 359372 158976 359424 158982
rect 359372 158918 359424 158924
rect 359188 157956 359240 157962
rect 359188 157898 359240 157904
rect 358912 156460 358964 156466
rect 358912 156402 358964 156408
rect 359476 6458 359504 248270
rect 359568 156602 359596 307906
rect 360304 306270 360332 310420
rect 360488 306354 360516 310420
rect 360672 306746 360700 310420
rect 360660 306740 360712 306746
rect 360660 306682 360712 306688
rect 360856 306626 360884 310420
rect 360396 306326 360516 306354
rect 360580 306598 360884 306626
rect 360200 306264 360252 306270
rect 360200 306206 360252 306212
rect 360292 306264 360344 306270
rect 360292 306206 360344 306212
rect 360212 305318 360240 306206
rect 360292 305856 360344 305862
rect 360292 305798 360344 305804
rect 360304 305386 360332 305798
rect 360292 305380 360344 305386
rect 360292 305322 360344 305328
rect 360200 305312 360252 305318
rect 360200 305254 360252 305260
rect 360292 253836 360344 253842
rect 360292 253778 360344 253784
rect 360200 250368 360252 250374
rect 360200 250310 360252 250316
rect 359646 243672 359702 243681
rect 359646 243607 359702 243616
rect 359660 158001 359688 243607
rect 359646 157992 359702 158001
rect 359646 157927 359702 157936
rect 359556 156596 359608 156602
rect 359556 156538 359608 156544
rect 360212 6798 360240 250310
rect 360304 9178 360332 253778
rect 360396 158166 360424 306326
rect 360580 306218 360608 306598
rect 360660 306468 360712 306474
rect 360660 306410 360712 306416
rect 360488 306190 360608 306218
rect 360384 158160 360436 158166
rect 360384 158102 360436 158108
rect 360488 157894 360516 306190
rect 360568 305856 360620 305862
rect 360568 305798 360620 305804
rect 360476 157888 360528 157894
rect 360476 157830 360528 157836
rect 360580 157826 360608 305798
rect 360672 159186 360700 306410
rect 361040 306354 361068 310420
rect 360764 306326 361068 306354
rect 360764 159254 360792 306326
rect 360844 306264 360896 306270
rect 360844 306206 360896 306212
rect 360752 159248 360804 159254
rect 360752 159190 360804 159196
rect 360660 159180 360712 159186
rect 360660 159122 360712 159128
rect 360856 159050 360884 306206
rect 361224 305862 361252 310420
rect 362130 308272 362186 308281
rect 362130 308207 362186 308216
rect 361212 305856 361264 305862
rect 361212 305798 361264 305804
rect 362040 305448 362092 305454
rect 362040 305390 362092 305396
rect 361948 248056 362000 248062
rect 361948 247998 362000 248004
rect 361580 245540 361632 245546
rect 361580 245482 361632 245488
rect 360936 245268 360988 245274
rect 360936 245210 360988 245216
rect 360844 159044 360896 159050
rect 360844 158986 360896 158992
rect 360568 157820 360620 157826
rect 360568 157762 360620 157768
rect 360292 9172 360344 9178
rect 360292 9114 360344 9120
rect 360200 6792 360252 6798
rect 360200 6734 360252 6740
rect 360948 6662 360976 245210
rect 361028 243772 361080 243778
rect 361028 243714 361080 243720
rect 361040 153882 361068 243714
rect 361118 158808 361174 158817
rect 361118 158743 361174 158752
rect 361028 153876 361080 153882
rect 361028 153818 361080 153824
rect 361132 6914 361160 158743
rect 361040 6886 361160 6914
rect 360936 6656 360988 6662
rect 360936 6598 360988 6604
rect 359464 6452 359516 6458
rect 359464 6394 359516 6400
rect 358176 6384 358228 6390
rect 358176 6326 358228 6332
rect 361040 3738 361068 6886
rect 361592 3806 361620 245482
rect 361764 245472 361816 245478
rect 361764 245414 361816 245420
rect 361672 245336 361724 245342
rect 361672 245278 361724 245284
rect 361580 3800 361632 3806
rect 361580 3742 361632 3748
rect 361028 3732 361080 3738
rect 361028 3674 361080 3680
rect 358084 3528 358136 3534
rect 358084 3470 358136 3476
rect 358726 3496 358782 3505
rect 358726 3431 358782 3440
rect 359922 3496 359978 3505
rect 359922 3431 359978 3440
rect 361118 3496 361174 3505
rect 361118 3431 361174 3440
rect 358740 480 358768 3431
rect 359936 480 359964 3431
rect 361132 480 361160 3431
rect 361684 3330 361712 245278
rect 361672 3324 361724 3330
rect 361672 3266 361724 3272
rect 361776 3262 361804 245414
rect 361856 245404 361908 245410
rect 361856 245346 361908 245352
rect 361764 3256 361816 3262
rect 361764 3198 361816 3204
rect 361868 3194 361896 245346
rect 361960 6730 361988 247998
rect 362052 155786 362080 305390
rect 362144 159497 362172 308207
rect 362236 259418 362264 444110
rect 362500 443148 362552 443154
rect 362500 443090 362552 443096
rect 362408 442060 362460 442066
rect 362408 442002 362460 442008
rect 362316 441992 362368 441998
rect 362316 441934 362368 441940
rect 362328 325650 362356 441934
rect 362420 379506 362448 442002
rect 362512 405686 362540 443090
rect 363604 440564 363656 440570
rect 363604 440506 363656 440512
rect 363616 419490 363644 440506
rect 371976 440428 372028 440434
rect 371976 440370 372028 440376
rect 363604 419484 363656 419490
rect 363604 419426 363656 419432
rect 362500 405680 362552 405686
rect 362500 405622 362552 405628
rect 362408 379500 362460 379506
rect 362408 379442 362460 379448
rect 362316 325644 362368 325650
rect 362316 325586 362368 325592
rect 367560 309120 367612 309126
rect 366454 309088 366510 309097
rect 367560 309062 367612 309068
rect 366454 309023 366510 309032
rect 366180 308984 366232 308990
rect 366180 308926 366232 308932
rect 366270 308952 366326 308961
rect 363512 308780 363564 308786
rect 363512 308722 363564 308728
rect 362316 300484 362368 300490
rect 362316 300426 362368 300432
rect 362224 259412 362276 259418
rect 362224 259354 362276 259360
rect 362224 243840 362276 243846
rect 362224 243782 362276 243788
rect 362130 159488 362186 159497
rect 362130 159423 362186 159432
rect 362040 155780 362092 155786
rect 362040 155722 362092 155728
rect 362236 153950 362264 243782
rect 362328 155553 362356 300426
rect 363236 251116 363288 251122
rect 363236 251058 363288 251064
rect 362960 248396 363012 248402
rect 362960 248338 363012 248344
rect 362408 243908 362460 243914
rect 362408 243850 362460 243856
rect 362420 158273 362448 243850
rect 362406 158264 362462 158273
rect 362406 158199 362462 158208
rect 362314 155544 362370 155553
rect 362314 155479 362370 155488
rect 362224 153944 362276 153950
rect 362224 153886 362276 153892
rect 361948 6724 362000 6730
rect 361948 6666 362000 6672
rect 362972 4146 363000 248338
rect 363052 248192 363104 248198
rect 363052 248134 363104 248140
rect 362960 4140 363012 4146
rect 362960 4082 363012 4088
rect 363064 4010 363092 248134
rect 363144 247648 363196 247654
rect 363144 247590 363196 247596
rect 363052 4004 363104 4010
rect 363052 3946 363104 3952
rect 362316 3596 362368 3602
rect 362316 3538 362368 3544
rect 361856 3188 361908 3194
rect 361856 3130 361908 3136
rect 362328 480 362356 3538
rect 363156 2961 363184 247590
rect 363248 6050 363276 251058
rect 363328 250912 363380 250918
rect 363328 250854 363380 250860
rect 363340 6866 363368 250854
rect 363418 243808 363474 243817
rect 363418 243743 363474 243752
rect 363432 9314 363460 243743
rect 363524 155378 363552 308722
rect 365076 308304 365128 308310
rect 365076 308246 365128 308252
rect 364892 308032 364944 308038
rect 364892 307974 364944 307980
rect 363604 303000 363656 303006
rect 363604 302942 363656 302948
rect 363512 155372 363564 155378
rect 363512 155314 363564 155320
rect 363616 154018 363644 302942
rect 363696 302728 363748 302734
rect 363696 302670 363748 302676
rect 363708 158778 363736 302670
rect 364524 253700 364576 253706
rect 364524 253642 364576 253648
rect 364432 248260 364484 248266
rect 364432 248202 364484 248208
rect 364340 248124 364392 248130
rect 364340 248066 364392 248072
rect 363788 243704 363840 243710
rect 363788 243646 363840 243652
rect 363696 158772 363748 158778
rect 363696 158714 363748 158720
rect 363800 158409 363828 243646
rect 363786 158400 363842 158409
rect 363786 158335 363842 158344
rect 363604 154012 363656 154018
rect 363604 153954 363656 153960
rect 363420 9308 363472 9314
rect 363420 9250 363472 9256
rect 363328 6860 363380 6866
rect 363328 6802 363380 6808
rect 363236 6044 363288 6050
rect 363236 5986 363288 5992
rect 364352 4078 364380 248066
rect 364340 4072 364392 4078
rect 364340 4014 364392 4020
rect 363510 3496 363566 3505
rect 363510 3431 363566 3440
rect 363142 2952 363198 2961
rect 363142 2887 363198 2896
rect 363524 480 363552 3431
rect 364444 3398 364472 248202
rect 364536 9042 364564 253642
rect 364616 251048 364668 251054
rect 364616 250990 364668 250996
rect 364524 9036 364576 9042
rect 364524 8978 364576 8984
rect 364628 5982 364656 250990
rect 364708 250980 364760 250986
rect 364708 250922 364760 250928
rect 364720 6118 364748 250922
rect 364800 244792 364852 244798
rect 364800 244734 364852 244740
rect 364812 6526 364840 244734
rect 364904 157146 364932 307974
rect 364984 305720 365036 305726
rect 364984 305662 365036 305668
rect 364996 157282 365024 305662
rect 365088 159225 365116 308246
rect 365168 302932 365220 302938
rect 365168 302874 365220 302880
rect 365074 159216 365130 159225
rect 365074 159151 365130 159160
rect 365180 158137 365208 302874
rect 365812 251184 365864 251190
rect 365812 251126 365864 251132
rect 365720 250436 365772 250442
rect 365720 250378 365772 250384
rect 365258 158808 365314 158817
rect 365258 158743 365314 158752
rect 365166 158128 365222 158137
rect 365166 158063 365222 158072
rect 364984 157276 365036 157282
rect 364984 157218 365036 157224
rect 364892 157140 364944 157146
rect 364892 157082 364944 157088
rect 364800 6520 364852 6526
rect 364800 6462 364852 6468
rect 364708 6112 364760 6118
rect 364708 6054 364760 6060
rect 364616 5976 364668 5982
rect 364616 5918 364668 5924
rect 365272 3670 365300 158743
rect 365260 3664 365312 3670
rect 365260 3606 365312 3612
rect 365732 3534 365760 250378
rect 365824 6769 365852 251126
rect 365904 250776 365956 250782
rect 365904 250718 365956 250724
rect 365810 6760 365866 6769
rect 365810 6695 365866 6704
rect 365916 6594 365944 250718
rect 365996 244860 366048 244866
rect 365996 244802 366048 244808
rect 366008 8974 366036 244802
rect 366088 243636 366140 243642
rect 366088 243578 366140 243584
rect 366100 9110 366128 243578
rect 366192 155922 366220 308926
rect 366270 308887 366326 308896
rect 366284 157865 366312 308887
rect 366364 308100 366416 308106
rect 366364 308042 366416 308048
rect 366376 158846 366404 308042
rect 366468 158953 366496 309023
rect 367376 308916 367428 308922
rect 367376 308858 367428 308864
rect 367284 308712 367336 308718
rect 367284 308654 367336 308660
rect 367098 303376 367154 303385
rect 367098 303311 367154 303320
rect 366548 302864 366600 302870
rect 366548 302806 366600 302812
rect 366454 158944 366510 158953
rect 366454 158879 366510 158888
rect 366364 158840 366416 158846
rect 366364 158782 366416 158788
rect 366270 157856 366326 157865
rect 366270 157791 366326 157800
rect 366560 157690 366588 302806
rect 366548 157684 366600 157690
rect 366548 157626 366600 157632
rect 366180 155916 366232 155922
rect 366180 155858 366232 155864
rect 366088 9104 366140 9110
rect 366088 9046 366140 9052
rect 365996 8968 366048 8974
rect 365996 8910 366048 8916
rect 365904 6588 365956 6594
rect 365904 6530 365956 6536
rect 365810 3632 365866 3641
rect 365810 3567 365866 3576
rect 365720 3528 365772 3534
rect 364614 3496 364670 3505
rect 365720 3470 365772 3476
rect 364614 3431 364670 3440
rect 364432 3392 364484 3398
rect 364432 3334 364484 3340
rect 364628 480 364656 3431
rect 365824 480 365852 3567
rect 367006 3496 367062 3505
rect 367112 3466 367140 303311
rect 367192 253768 367244 253774
rect 367192 253710 367244 253716
rect 367204 9246 367232 253710
rect 367296 155446 367324 308654
rect 367388 155718 367416 308858
rect 367468 307896 367520 307902
rect 367468 307838 367520 307844
rect 367480 157010 367508 307838
rect 367572 157078 367600 309062
rect 367836 309052 367888 309058
rect 367836 308994 367888 309000
rect 367652 308372 367704 308378
rect 367652 308314 367704 308320
rect 367664 157214 367692 308314
rect 367744 305516 367796 305522
rect 367744 305458 367796 305464
rect 367652 157208 367704 157214
rect 367652 157150 367704 157156
rect 367560 157072 367612 157078
rect 367560 157014 367612 157020
rect 367468 157004 367520 157010
rect 367468 156946 367520 156952
rect 367376 155712 367428 155718
rect 367376 155654 367428 155660
rect 367284 155440 367336 155446
rect 367284 155382 367336 155388
rect 367756 155038 367784 305458
rect 367848 158574 367876 308994
rect 368570 308816 368626 308825
rect 368570 308751 368626 308760
rect 368480 253632 368532 253638
rect 368480 253574 368532 253580
rect 367928 243976 367980 243982
rect 367928 243918 367980 243924
rect 367836 158568 367888 158574
rect 367836 158510 367888 158516
rect 367940 155281 367968 243918
rect 367926 155272 367982 155281
rect 367926 155207 367982 155216
rect 367744 155032 367796 155038
rect 367744 154974 367796 154980
rect 367192 9240 367244 9246
rect 367192 9182 367244 9188
rect 368492 6254 368520 253574
rect 368584 157185 368612 308751
rect 370042 308680 370098 308689
rect 369952 308644 370004 308650
rect 370042 308615 370098 308624
rect 369952 308586 370004 308592
rect 369030 306232 369086 306241
rect 368664 306196 368716 306202
rect 369030 306167 369086 306176
rect 368664 306138 368716 306144
rect 368570 157176 368626 157185
rect 368570 157111 368626 157120
rect 368676 155854 368704 306138
rect 368940 305584 368992 305590
rect 368940 305526 368992 305532
rect 368848 305380 368900 305386
rect 368848 305322 368900 305328
rect 368756 305312 368808 305318
rect 368756 305254 368808 305260
rect 368664 155848 368716 155854
rect 368664 155790 368716 155796
rect 368768 155310 368796 305254
rect 368860 157350 368888 305322
rect 368848 157344 368900 157350
rect 368848 157286 368900 157292
rect 368952 156942 368980 305526
rect 369044 157049 369072 306167
rect 369124 302796 369176 302802
rect 369124 302738 369176 302744
rect 369136 158506 369164 302738
rect 369860 247512 369912 247518
rect 369860 247454 369912 247460
rect 369308 243568 369360 243574
rect 369308 243510 369360 243516
rect 369216 242208 369268 242214
rect 369216 242150 369268 242156
rect 369124 158500 369176 158506
rect 369124 158442 369176 158448
rect 369030 157040 369086 157049
rect 369030 156975 369086 156984
rect 368940 156936 368992 156942
rect 368940 156878 368992 156884
rect 368756 155304 368808 155310
rect 368756 155246 368808 155252
rect 369228 152590 369256 242150
rect 369320 159361 369348 243510
rect 369306 159352 369362 159361
rect 369306 159287 369362 159296
rect 369216 152584 369268 152590
rect 369216 152526 369268 152532
rect 369872 6322 369900 247454
rect 369964 155582 369992 308586
rect 370056 155961 370084 308615
rect 370504 308576 370556 308582
rect 370504 308518 370556 308524
rect 371330 308544 371386 308553
rect 370134 306368 370190 306377
rect 370134 306303 370190 306312
rect 370412 306332 370464 306338
rect 370042 155952 370098 155961
rect 370042 155887 370098 155896
rect 370148 155825 370176 306303
rect 370412 306274 370464 306280
rect 370320 305924 370372 305930
rect 370320 305866 370372 305872
rect 370228 303340 370280 303346
rect 370228 303282 370280 303288
rect 370134 155816 370190 155825
rect 370134 155751 370190 155760
rect 369952 155576 370004 155582
rect 369952 155518 370004 155524
rect 370240 154562 370268 303282
rect 370332 156913 370360 305866
rect 370318 156904 370374 156913
rect 370318 156839 370374 156848
rect 370424 156670 370452 306274
rect 370516 158914 370544 308518
rect 371330 308479 371386 308488
rect 370688 303544 370740 303550
rect 370688 303486 370740 303492
rect 370596 300348 370648 300354
rect 370596 300290 370648 300296
rect 370504 158908 370556 158914
rect 370504 158850 370556 158856
rect 370412 156664 370464 156670
rect 370412 156606 370464 156612
rect 370228 154556 370280 154562
rect 370228 154498 370280 154504
rect 370608 152522 370636 300290
rect 370700 156534 370728 303486
rect 371240 250844 371292 250850
rect 371240 250786 371292 250792
rect 370688 156528 370740 156534
rect 370688 156470 370740 156476
rect 370596 152516 370648 152522
rect 370596 152458 370648 152464
rect 369860 6316 369912 6322
rect 369860 6258 369912 6264
rect 368480 6248 368532 6254
rect 368480 6190 368532 6196
rect 369400 3596 369452 3602
rect 369400 3538 369452 3544
rect 368202 3496 368258 3505
rect 367006 3431 367062 3440
rect 367100 3460 367152 3466
rect 367020 480 367048 3431
rect 368202 3431 368258 3440
rect 367100 3402 367152 3408
rect 368216 480 368244 3431
rect 369412 480 369440 3538
rect 370594 3496 370650 3505
rect 370594 3431 370650 3440
rect 370608 480 370636 3431
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371252 354 371280 250786
rect 371344 3670 371372 308479
rect 371424 306128 371476 306134
rect 371424 306070 371476 306076
rect 371436 155106 371464 306070
rect 371700 306060 371752 306066
rect 371700 306002 371752 306008
rect 371516 305992 371568 305998
rect 371516 305934 371568 305940
rect 371528 155174 371556 305934
rect 371608 305788 371660 305794
rect 371608 305730 371660 305736
rect 371620 155242 371648 305730
rect 371712 156806 371740 306002
rect 371792 305652 371844 305658
rect 371792 305594 371844 305600
rect 371804 156874 371832 305594
rect 371884 285116 371936 285122
rect 371884 285058 371936 285064
rect 371792 156868 371844 156874
rect 371792 156810 371844 156816
rect 371700 156800 371752 156806
rect 371700 156742 371752 156748
rect 371608 155236 371660 155242
rect 371608 155178 371660 155184
rect 371516 155168 371568 155174
rect 371516 155110 371568 155116
rect 371424 155100 371476 155106
rect 371424 155042 371476 155048
rect 371896 3942 371924 285058
rect 371988 167006 372016 440370
rect 372988 303476 373040 303482
rect 372988 303418 373040 303424
rect 372896 303272 372948 303278
rect 372896 303214 372948 303220
rect 372068 303136 372120 303142
rect 372068 303078 372120 303084
rect 371976 167000 372028 167006
rect 371976 166942 372028 166948
rect 372080 159089 372108 303078
rect 372620 296268 372672 296274
rect 372620 296210 372672 296216
rect 372066 159080 372122 159089
rect 372066 159015 372122 159024
rect 371884 3936 371936 3942
rect 371884 3878 371936 3884
rect 371332 3664 371384 3670
rect 371332 3606 371384 3612
rect 372632 3482 372660 296210
rect 372712 247988 372764 247994
rect 372712 247930 372764 247936
rect 372724 6186 372752 247930
rect 372804 245608 372856 245614
rect 372804 245550 372856 245556
rect 372712 6180 372764 6186
rect 372712 6122 372764 6128
rect 372816 3602 372844 245550
rect 372908 154494 372936 303214
rect 373000 155514 373028 303418
rect 373080 303408 373132 303414
rect 373080 303350 373132 303356
rect 373092 155650 373120 303350
rect 373172 303204 373224 303210
rect 373172 303146 373224 303152
rect 373184 157321 373212 303146
rect 373170 157312 373226 157321
rect 373170 157247 373226 157256
rect 373080 155644 373132 155650
rect 373080 155586 373132 155592
rect 372988 155508 373040 155514
rect 372988 155450 373040 155456
rect 372896 154488 372948 154494
rect 372896 154430 372948 154436
rect 373276 60722 373304 445810
rect 378784 444712 378836 444718
rect 378784 444654 378836 444660
rect 374736 441924 374788 441930
rect 374736 441866 374788 441872
rect 373448 303612 373500 303618
rect 373448 303554 373500 303560
rect 373356 303068 373408 303074
rect 373356 303010 373408 303016
rect 373368 157758 373396 303010
rect 373460 158234 373488 303554
rect 374092 301776 374144 301782
rect 374092 301718 374144 301724
rect 373448 158228 373500 158234
rect 373448 158170 373500 158176
rect 373356 157752 373408 157758
rect 373356 157694 373408 157700
rect 373264 60716 373316 60722
rect 373264 60658 373316 60664
rect 372804 3596 372856 3602
rect 372804 3538 372856 3544
rect 372632 3454 372936 3482
rect 372908 480 372936 3454
rect 374104 480 374132 301718
rect 374644 282396 374696 282402
rect 374644 282338 374696 282344
rect 374656 3058 374684 282338
rect 374748 179382 374776 441866
rect 377404 440496 377456 440502
rect 377404 440438 377456 440444
rect 377416 313274 377444 440438
rect 378796 365702 378824 444654
rect 578884 444440 578936 444446
rect 578884 444382 578936 444388
rect 388444 443216 388496 443222
rect 388444 443158 388496 443164
rect 378784 365696 378836 365702
rect 378784 365638 378836 365644
rect 377404 313268 377456 313274
rect 377404 313210 377456 313216
rect 378784 307216 378836 307222
rect 378784 307158 378836 307164
rect 377402 306096 377458 306105
rect 377402 306031 377458 306040
rect 376760 300416 376812 300422
rect 376760 300358 376812 300364
rect 374736 179376 374788 179382
rect 374736 179318 374788 179324
rect 376772 16574 376800 300358
rect 376772 16546 377352 16574
rect 375288 3936 375340 3942
rect 375288 3878 375340 3884
rect 374644 3052 374696 3058
rect 374644 2994 374696 3000
rect 375300 480 375328 3878
rect 377324 3482 377352 16546
rect 377416 3670 377444 306031
rect 378140 299056 378192 299062
rect 378140 298998 378192 299004
rect 378152 16574 378180 298998
rect 378152 16546 378456 16574
rect 377404 3664 377456 3670
rect 377404 3606 377456 3612
rect 377324 3454 377720 3482
rect 376484 3052 376536 3058
rect 376484 2994 376536 3000
rect 376496 480 376524 2994
rect 377692 480 377720 3454
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378428 354 378456 16546
rect 378796 2990 378824 307158
rect 385038 305824 385094 305833
rect 385038 305759 385094 305768
rect 381544 298988 381596 298994
rect 381544 298930 381596 298936
rect 381556 3602 381584 298930
rect 381636 297696 381688 297702
rect 381636 297638 381688 297644
rect 381544 3596 381596 3602
rect 381544 3538 381596 3544
rect 381648 3534 381676 297638
rect 382280 287972 382332 287978
rect 382280 287914 382332 287920
rect 381636 3528 381688 3534
rect 381636 3470 381688 3476
rect 379978 3360 380034 3369
rect 382292 3346 382320 287914
rect 382372 265872 382424 265878
rect 382372 265814 382424 265820
rect 382384 3466 382412 265814
rect 385052 16574 385080 305759
rect 387064 294772 387116 294778
rect 387064 294714 387116 294720
rect 386420 271244 386472 271250
rect 386420 271186 386472 271192
rect 386432 16574 386460 271186
rect 385052 16546 386000 16574
rect 386432 16546 386736 16574
rect 384764 3596 384816 3602
rect 384764 3538 384816 3544
rect 382372 3460 382424 3466
rect 382372 3402 382424 3408
rect 383568 3460 383620 3466
rect 383568 3402 383620 3408
rect 382292 3318 382412 3346
rect 379978 3295 380034 3304
rect 378784 2984 378836 2990
rect 378784 2926 378836 2932
rect 379992 480 380020 3295
rect 381176 2984 381228 2990
rect 381176 2926 381228 2932
rect 381188 480 381216 2926
rect 382384 480 382412 3318
rect 383580 480 383608 3402
rect 384776 480 384804 3538
rect 385972 480 386000 16546
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 378846 -960 378958 326
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 386708 354 386736 16546
rect 387076 3466 387104 294714
rect 387064 3460 387116 3466
rect 387064 3402 387116 3408
rect 388260 3460 388312 3466
rect 388260 3402 388312 3408
rect 388272 480 388300 3402
rect 388456 3398 388484 443158
rect 577596 441788 577648 441794
rect 577596 441730 577648 441736
rect 577504 441652 577556 441658
rect 577504 441594 577556 441600
rect 462962 308408 463018 308417
rect 462962 308343 463018 308352
rect 402980 307148 403032 307154
rect 402980 307090 403032 307096
rect 396722 303240 396778 303249
rect 396722 303175 396778 303184
rect 390560 283824 390612 283830
rect 390560 283766 390612 283772
rect 389180 264444 389232 264450
rect 389180 264386 389232 264392
rect 389192 16574 389220 264386
rect 389192 16546 389496 16574
rect 388444 3392 388496 3398
rect 388444 3334 388496 3340
rect 389468 480 389496 16546
rect 390572 3466 390600 283766
rect 393320 263152 393372 263158
rect 393320 263094 393372 263100
rect 390652 261860 390704 261866
rect 390652 261802 390704 261808
rect 390560 3460 390612 3466
rect 390560 3402 390612 3408
rect 390664 480 390692 261802
rect 391940 260364 391992 260370
rect 391940 260306 391992 260312
rect 391952 16574 391980 260306
rect 393332 16574 393360 263094
rect 396080 260296 396132 260302
rect 396080 260238 396132 260244
rect 394700 253564 394752 253570
rect 394700 253506 394752 253512
rect 394712 16574 394740 253506
rect 391952 16546 392624 16574
rect 393332 16546 394280 16574
rect 394712 16546 395384 16574
rect 391848 3460 391900 3466
rect 391848 3402 391900 3408
rect 391860 480 391888 3402
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387126 -960 387238 326
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 394252 480 394280 16546
rect 395356 480 395384 16546
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 260238
rect 396736 2990 396764 303175
rect 400220 270020 400272 270026
rect 400220 269962 400272 269968
rect 397460 263084 397512 263090
rect 397460 263026 397512 263032
rect 397472 16574 397500 263026
rect 398840 261792 398892 261798
rect 398840 261734 398892 261740
rect 397472 16546 397776 16574
rect 396724 2984 396776 2990
rect 396724 2926 396776 2932
rect 397748 480 397776 16546
rect 398852 3602 398880 261734
rect 398932 254788 398984 254794
rect 398932 254730 398984 254736
rect 398840 3596 398892 3602
rect 398840 3538 398892 3544
rect 398944 480 398972 254730
rect 400232 16574 400260 269962
rect 402992 16574 403020 307090
rect 452660 304428 452712 304434
rect 452660 304370 452712 304376
rect 412640 297628 412692 297634
rect 412640 297570 412692 297576
rect 405740 291916 405792 291922
rect 405740 291858 405792 291864
rect 404360 275528 404412 275534
rect 404360 275470 404412 275476
rect 400232 16546 400904 16574
rect 402992 16546 403664 16574
rect 400128 3596 400180 3602
rect 400128 3538 400180 3544
rect 400140 480 400168 3538
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 16546
rect 402520 2984 402572 2990
rect 402520 2926 402572 2932
rect 402532 480 402560 2926
rect 403636 480 403664 16546
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 275470
rect 405752 16574 405780 291858
rect 408500 290692 408552 290698
rect 408500 290634 408552 290640
rect 407120 279608 407172 279614
rect 407120 279550 407172 279556
rect 405752 16546 406056 16574
rect 406028 480 406056 16546
rect 407132 3482 407160 279550
rect 407212 267300 407264 267306
rect 407212 267242 407264 267248
rect 407224 3602 407252 267242
rect 408512 16574 408540 290634
rect 409880 278180 409932 278186
rect 409880 278122 409932 278128
rect 409892 16574 409920 278122
rect 408512 16546 409184 16574
rect 409892 16546 410840 16574
rect 407212 3596 407264 3602
rect 407212 3538 407264 3544
rect 408408 3596 408460 3602
rect 408408 3538 408460 3544
rect 407132 3454 407252 3482
rect 407224 480 407252 3454
rect 408420 480 408448 3538
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 410812 480 410840 16546
rect 411904 3664 411956 3670
rect 411904 3606 411956 3612
rect 411916 480 411944 3606
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 297570
rect 421564 296200 421616 296206
rect 421564 296142 421616 296148
rect 418160 290624 418212 290630
rect 418160 290566 418212 290572
rect 414664 282328 414716 282334
rect 414664 282270 414716 282276
rect 413284 256420 413336 256426
rect 413284 256362 413336 256368
rect 413296 3058 413324 256362
rect 414020 249484 414072 249490
rect 414020 249426 414072 249432
rect 414032 16574 414060 249426
rect 414032 16546 414336 16574
rect 413284 3052 413336 3058
rect 413284 2994 413336 3000
rect 414308 480 414336 16546
rect 414676 3466 414704 282270
rect 417424 280900 417476 280906
rect 417424 280842 417476 280848
rect 416780 250708 416832 250714
rect 416780 250650 416832 250656
rect 416792 6914 416820 250650
rect 417436 16574 417464 280842
rect 418172 16574 418200 290566
rect 420920 269952 420972 269958
rect 420920 269894 420972 269900
rect 417436 16546 417556 16574
rect 418172 16546 418568 16574
rect 416792 6886 417464 6914
rect 414664 3460 414716 3466
rect 414664 3402 414716 3408
rect 416688 3460 416740 3466
rect 416688 3402 416740 3408
rect 415492 3052 415544 3058
rect 415492 2994 415544 3000
rect 415504 480 415532 2994
rect 416700 480 416728 3402
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 6886
rect 417528 3058 417556 16546
rect 417516 3052 417568 3058
rect 417516 2994 417568 3000
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 418540 354 418568 16546
rect 420184 3052 420236 3058
rect 420184 2994 420236 3000
rect 420196 480 420224 2994
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 269894
rect 421576 3602 421604 296142
rect 422300 296132 422352 296138
rect 422300 296074 422352 296080
rect 422312 16574 422340 296074
rect 430580 289264 430632 289270
rect 430580 289206 430632 289212
rect 423680 279540 423732 279546
rect 423680 279482 423732 279488
rect 422312 16546 422616 16574
rect 421564 3596 421616 3602
rect 421564 3538 421616 3544
rect 422588 480 422616 16546
rect 423692 3346 423720 279482
rect 428464 278112 428516 278118
rect 428464 278054 428516 278060
rect 425060 256284 425112 256290
rect 425060 256226 425112 256232
rect 423772 247920 423824 247926
rect 423772 247862 423824 247868
rect 423784 3534 423812 247862
rect 425072 16574 425100 256226
rect 427820 252136 427872 252142
rect 427820 252078 427872 252084
rect 425072 16546 425744 16574
rect 423772 3528 423824 3534
rect 423772 3470 423824 3476
rect 424968 3528 425020 3534
rect 424968 3470 425020 3476
rect 423692 3318 423812 3346
rect 423784 480 423812 3318
rect 424980 480 425008 3470
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 16546
rect 427832 6914 427860 252078
rect 428476 16574 428504 278054
rect 430592 16574 430620 289206
rect 442264 283756 442316 283762
rect 442264 283698 442316 283704
rect 440240 264376 440292 264382
rect 440240 264318 440292 264324
rect 436100 263016 436152 263022
rect 436100 262958 436152 262964
rect 434720 258868 434772 258874
rect 434720 258810 434772 258816
rect 431960 256216 432012 256222
rect 431960 256158 432012 256164
rect 428476 16546 428596 16574
rect 430592 16546 430896 16574
rect 427832 6886 428504 6914
rect 427268 3596 427320 3602
rect 427268 3538 427320 3544
rect 427280 480 427308 3538
rect 428476 480 428504 6886
rect 428568 3330 428596 16546
rect 429660 3528 429712 3534
rect 429660 3470 429712 3476
rect 428556 3324 428608 3330
rect 428556 3266 428608 3272
rect 429672 480 429700 3470
rect 430868 480 430896 16546
rect 431972 3534 432000 256158
rect 432052 252068 432104 252074
rect 432052 252010 432104 252016
rect 431960 3528 432012 3534
rect 431960 3470 432012 3476
rect 432064 480 432092 252010
rect 434732 16574 434760 258810
rect 436112 16574 436140 262958
rect 438860 261724 438912 261730
rect 438860 261666 438912 261672
rect 437480 253428 437532 253434
rect 437480 253370 437532 253376
rect 434732 16546 435128 16574
rect 436112 16546 436784 16574
rect 433248 3528 433300 3534
rect 433248 3470 433300 3476
rect 433260 480 433288 3470
rect 434444 3324 434496 3330
rect 434444 3266 434496 3272
rect 434456 480 434484 3266
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426134 -960 426246 326
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435100 354 435128 16546
rect 436756 480 436784 16546
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437492 354 437520 253370
rect 438872 16574 438900 261666
rect 438872 16546 439176 16574
rect 439148 480 439176 16546
rect 440252 3346 440280 264318
rect 441620 262948 441672 262954
rect 441620 262890 441672 262896
rect 440332 256148 440384 256154
rect 440332 256090 440384 256096
rect 440344 3534 440372 256090
rect 441632 16574 441660 262890
rect 441632 16546 442212 16574
rect 440332 3528 440384 3534
rect 440332 3470 440384 3476
rect 441528 3528 441580 3534
rect 441528 3470 441580 3476
rect 442184 3482 442212 16546
rect 442276 3602 442304 283698
rect 445024 276820 445076 276826
rect 445024 276762 445076 276768
rect 443000 264308 443052 264314
rect 443000 264250 443052 264256
rect 443012 16574 443040 264250
rect 443644 254720 443696 254726
rect 443644 254662 443696 254668
rect 443012 16546 443408 16574
rect 442264 3596 442316 3602
rect 442264 3538 442316 3544
rect 440252 3318 440372 3346
rect 440344 480 440372 3318
rect 441540 480 441568 3470
rect 442184 3454 442672 3482
rect 442644 480 442672 3454
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 354 443408 16546
rect 443656 3534 443684 254662
rect 445036 16574 445064 276762
rect 448520 276752 448572 276758
rect 448520 276694 448572 276700
rect 446404 274168 446456 274174
rect 446404 274110 446456 274116
rect 445760 245200 445812 245206
rect 445760 245142 445812 245148
rect 445036 16546 445156 16574
rect 445128 3602 445156 16546
rect 445024 3596 445076 3602
rect 445024 3538 445076 3544
rect 445116 3596 445168 3602
rect 445116 3538 445168 3544
rect 443644 3528 443696 3534
rect 443644 3470 443696 3476
rect 445036 480 445064 3538
rect 443798 354 443910 480
rect 443380 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 445772 354 445800 245142
rect 446416 3262 446444 274110
rect 448532 3534 448560 276694
rect 448612 275460 448664 275466
rect 448612 275402 448664 275408
rect 447416 3528 447468 3534
rect 447416 3470 447468 3476
rect 448520 3528 448572 3534
rect 448520 3470 448572 3476
rect 446404 3256 446456 3262
rect 446404 3198 446456 3204
rect 447428 480 447456 3470
rect 448624 480 448652 275402
rect 449900 262880 449952 262886
rect 449900 262822 449952 262828
rect 449912 16574 449940 262822
rect 452672 16574 452700 304370
rect 457444 294704 457496 294710
rect 457444 294646 457496 294652
rect 454684 286476 454736 286482
rect 454684 286418 454736 286424
rect 454040 256080 454092 256086
rect 454040 256022 454092 256028
rect 449912 16546 450952 16574
rect 452672 16546 453344 16574
rect 449808 3528 449860 3534
rect 449808 3470 449860 3476
rect 449820 480 449848 3470
rect 450924 480 450952 16546
rect 452108 3256 452160 3262
rect 452108 3198 452160 3204
rect 452120 480 452148 3198
rect 453316 480 453344 16546
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454052 354 454080 256022
rect 454696 3534 454724 286418
rect 455420 249416 455472 249422
rect 455420 249358 455472 249364
rect 455432 16574 455460 249358
rect 455432 16546 455736 16574
rect 454684 3528 454736 3534
rect 454684 3470 454736 3476
rect 455708 480 455736 16546
rect 456892 3528 456944 3534
rect 456892 3470 456944 3476
rect 456904 480 456932 3470
rect 457456 2990 457484 294646
rect 460204 287904 460256 287910
rect 460204 287846 460256 287852
rect 458824 286408 458876 286414
rect 458824 286350 458876 286356
rect 458836 3602 458864 286350
rect 459560 274032 459612 274038
rect 459560 273974 459612 273980
rect 459572 16574 459600 273974
rect 459572 16546 459968 16574
rect 458088 3596 458140 3602
rect 458088 3538 458140 3544
rect 458824 3596 458876 3602
rect 458824 3538 458876 3544
rect 457444 2984 457496 2990
rect 457444 2926 457496 2932
rect 458100 480 458128 3538
rect 459192 2984 459244 2990
rect 459192 2926 459244 2932
rect 459204 480 459232 2926
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 460216 4146 460244 287846
rect 460940 274100 460992 274106
rect 460940 274042 460992 274048
rect 460952 16574 460980 274042
rect 460952 16546 461624 16574
rect 460204 4140 460256 4146
rect 460204 4082 460256 4088
rect 461596 480 461624 16546
rect 462780 4140 462832 4146
rect 462780 4082 462832 4088
rect 462792 480 462820 4082
rect 462976 3534 463004 308343
rect 543740 307080 543792 307086
rect 543740 307022 543792 307028
rect 485044 304360 485096 304366
rect 485044 304302 485096 304308
rect 463700 300280 463752 300286
rect 463700 300222 463752 300228
rect 463712 16574 463740 300222
rect 467104 293412 467156 293418
rect 467104 293354 467156 293360
rect 464344 282260 464396 282266
rect 464344 282202 464396 282208
rect 463712 16546 464016 16574
rect 462964 3528 463016 3534
rect 462964 3470 463016 3476
rect 463988 480 464016 16546
rect 464356 3058 464384 282202
rect 466460 252000 466512 252006
rect 466460 251942 466512 251948
rect 466472 16574 466500 251942
rect 466472 16546 467052 16574
rect 465172 3596 465224 3602
rect 465172 3538 465224 3544
rect 464344 3052 464396 3058
rect 464344 2994 464396 3000
rect 465184 480 465212 3538
rect 467024 3482 467052 16546
rect 467116 3602 467144 293354
rect 471244 285048 471296 285054
rect 471244 284990 471296 284996
rect 468484 275392 468536 275398
rect 468484 275334 468536 275340
rect 467840 249280 467892 249286
rect 467840 249222 467892 249228
rect 467852 16574 467880 249222
rect 467852 16546 468248 16574
rect 467104 3596 467156 3602
rect 467104 3538 467156 3544
rect 467024 3454 467512 3482
rect 466276 3052 466328 3058
rect 466276 2994 466328 3000
rect 466288 480 466316 2994
rect 467484 480 467512 3454
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468220 354 468248 16546
rect 468496 4146 468524 275334
rect 468484 4140 468536 4146
rect 468484 4082 468536 4088
rect 471060 4140 471112 4146
rect 471060 4082 471112 4088
rect 469864 3596 469916 3602
rect 469864 3538 469916 3544
rect 469876 480 469904 3538
rect 471072 480 471100 4082
rect 471256 3534 471284 284990
rect 475384 272536 475436 272542
rect 475384 272478 475436 272484
rect 473452 268456 473504 268462
rect 473452 268398 473504 268404
rect 471980 246696 472032 246702
rect 471980 246638 472032 246644
rect 471992 16574 472020 246638
rect 473464 16574 473492 268398
rect 474740 268388 474792 268394
rect 474740 268330 474792 268336
rect 474752 16574 474780 268330
rect 471992 16546 472296 16574
rect 473464 16546 474136 16574
rect 474752 16546 475332 16574
rect 471244 3528 471296 3534
rect 471244 3470 471296 3476
rect 472268 480 472296 16546
rect 473452 3528 473504 3534
rect 473452 3470 473504 3476
rect 473464 480 473492 3470
rect 468638 354 468750 480
rect 468220 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 16546
rect 475304 3482 475332 16546
rect 475396 3602 475424 272478
rect 484400 250640 484452 250646
rect 484400 250582 484452 250588
rect 477500 249212 477552 249218
rect 477500 249154 477552 249160
rect 477512 16574 477540 249154
rect 480260 246628 480312 246634
rect 480260 246570 480312 246576
rect 480272 16574 480300 246570
rect 483020 246560 483072 246566
rect 483020 246502 483072 246508
rect 481732 245132 481784 245138
rect 481732 245074 481784 245080
rect 481640 245064 481692 245070
rect 481640 245006 481692 245012
rect 477512 16546 478184 16574
rect 480272 16546 480576 16574
rect 475384 3596 475436 3602
rect 475384 3538 475436 3544
rect 476948 3596 477000 3602
rect 476948 3538 477000 3544
rect 475304 3454 475792 3482
rect 475764 480 475792 3454
rect 476960 480 476988 3538
rect 478156 480 478184 16546
rect 479340 3528 479392 3534
rect 479340 3470 479392 3476
rect 479352 480 479380 3470
rect 480548 480 480576 16546
rect 481652 3534 481680 245006
rect 481640 3528 481692 3534
rect 481640 3470 481692 3476
rect 481744 480 481772 245074
rect 483032 16574 483060 246502
rect 484412 16574 484440 250582
rect 483032 16546 484072 16574
rect 484412 16546 484808 16574
rect 482468 3528 482520 3534
rect 482468 3470 482520 3476
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482480 354 482508 3470
rect 484044 480 484072 16546
rect 482806 354 482918 480
rect 482480 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 485056 3194 485084 304302
rect 514024 304292 514076 304298
rect 514024 304234 514076 304240
rect 489182 303104 489238 303113
rect 489182 303039 489238 303048
rect 486424 269884 486476 269890
rect 486424 269826 486476 269832
rect 485780 246492 485832 246498
rect 485780 246434 485832 246440
rect 485792 6914 485820 246434
rect 486436 16574 486464 269826
rect 486436 16546 486556 16574
rect 485792 6886 486464 6914
rect 485044 3188 485096 3194
rect 485044 3130 485096 3136
rect 486436 480 486464 6886
rect 486528 3058 486556 16546
rect 489196 3738 489224 303039
rect 494060 301572 494112 301578
rect 494060 301514 494112 301520
rect 490012 289196 490064 289202
rect 490012 289138 490064 289144
rect 490024 6914 490052 289138
rect 493324 279472 493376 279478
rect 493324 279414 493376 279420
rect 491300 265804 491352 265810
rect 491300 265746 491352 265752
rect 491312 16574 491340 265746
rect 492680 246424 492732 246430
rect 492680 246366 492732 246372
rect 492692 16574 492720 246366
rect 491312 16546 492352 16574
rect 492692 16546 493088 16574
rect 489932 6886 490052 6914
rect 489184 3732 489236 3738
rect 489184 3674 489236 3680
rect 487620 3188 487672 3194
rect 487620 3130 487672 3136
rect 486516 3052 486568 3058
rect 486516 2994 486568 3000
rect 487632 480 487660 3130
rect 488816 3052 488868 3058
rect 488816 2994 488868 3000
rect 488828 480 488856 2994
rect 489932 480 489960 6886
rect 491116 3732 491168 3738
rect 491116 3674 491168 3680
rect 491128 480 491156 3674
rect 492324 480 492352 16546
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 493336 3398 493364 279414
rect 494072 16574 494100 301514
rect 498292 300212 498344 300218
rect 498292 300154 498344 300160
rect 495440 267164 495492 267170
rect 495440 267106 495492 267112
rect 494072 16546 494744 16574
rect 493324 3392 493376 3398
rect 493324 3334 493376 3340
rect 494716 480 494744 16546
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 267106
rect 496084 253360 496136 253366
rect 496084 253302 496136 253308
rect 496096 3534 496124 253302
rect 498304 6914 498332 300154
rect 500224 298920 500276 298926
rect 500224 298862 500276 298868
rect 499580 253292 499632 253298
rect 499580 253234 499632 253240
rect 499592 16574 499620 253234
rect 499592 16546 500172 16574
rect 498212 6886 498332 6914
rect 496084 3528 496136 3534
rect 496084 3470 496136 3476
rect 497096 3528 497148 3534
rect 497096 3470 497148 3476
rect 497108 480 497136 3470
rect 498212 480 498240 6886
rect 500144 3482 500172 16546
rect 500236 3602 500264 298862
rect 509884 293344 509936 293350
rect 509884 293286 509936 293292
rect 506480 261656 506532 261662
rect 506480 261598 506532 261604
rect 503720 250572 503772 250578
rect 503720 250514 503772 250520
rect 502340 247852 502392 247858
rect 502340 247794 502392 247800
rect 502352 16574 502380 247794
rect 502352 16546 503024 16574
rect 500224 3596 500276 3602
rect 500224 3538 500276 3544
rect 501788 3596 501840 3602
rect 501788 3538 501840 3544
rect 500144 3454 500632 3482
rect 499396 3392 499448 3398
rect 499396 3334 499448 3340
rect 499408 480 499436 3334
rect 500604 480 500632 3454
rect 501800 480 501828 3538
rect 502996 480 503024 16546
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503732 354 503760 250514
rect 505100 247784 505152 247790
rect 505100 247726 505152 247732
rect 505112 16574 505140 247726
rect 505112 16546 505416 16574
rect 505388 480 505416 16546
rect 506492 3534 506520 261598
rect 509240 257508 509292 257514
rect 509240 257450 509292 257456
rect 506572 256012 506624 256018
rect 506572 255954 506624 255960
rect 506480 3528 506532 3534
rect 506480 3470 506532 3476
rect 506584 3380 506612 255954
rect 507860 247716 507912 247722
rect 507860 247658 507912 247664
rect 507872 16574 507900 247658
rect 509252 16574 509280 257450
rect 507872 16546 508912 16574
rect 509252 16546 509648 16574
rect 507308 3528 507360 3534
rect 507308 3470 507360 3476
rect 506492 3352 506612 3380
rect 506492 480 506520 3352
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507320 354 507348 3470
rect 508884 480 508912 16546
rect 507646 354 507758 480
rect 507320 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 509896 3330 509924 293286
rect 511264 276684 511316 276690
rect 511264 276626 511316 276632
rect 510620 261588 510672 261594
rect 510620 261530 510672 261536
rect 510632 16574 510660 261530
rect 510632 16546 511212 16574
rect 511184 3482 511212 16546
rect 511276 3602 511304 276626
rect 512000 249144 512052 249150
rect 512000 249086 512052 249092
rect 511264 3596 511316 3602
rect 511264 3538 511316 3544
rect 511184 3454 511304 3482
rect 509884 3324 509936 3330
rect 509884 3266 509936 3272
rect 511276 480 511304 3454
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 249086
rect 513564 3596 513616 3602
rect 513564 3538 513616 3544
rect 513576 480 513604 3538
rect 514036 3058 514064 304234
rect 520922 302968 520978 302977
rect 520922 302903 520978 302912
rect 516784 296064 516836 296070
rect 516784 296006 516836 296012
rect 516140 246356 516192 246362
rect 516140 246298 516192 246304
rect 516152 16574 516180 246298
rect 516152 16546 516732 16574
rect 516704 3482 516732 16546
rect 516796 3874 516824 296006
rect 518164 287768 518216 287774
rect 518164 287710 518216 287716
rect 517520 271176 517572 271182
rect 517520 271118 517572 271124
rect 517532 16574 517560 271118
rect 517532 16546 517928 16574
rect 516784 3868 516836 3874
rect 516784 3810 516836 3816
rect 516704 3454 517192 3482
rect 514760 3324 514812 3330
rect 514760 3266 514812 3272
rect 514024 3052 514076 3058
rect 514024 2994 514076 3000
rect 514772 480 514800 3266
rect 515956 3052 516008 3058
rect 515956 2994 516008 3000
rect 515968 480 515996 2994
rect 517164 480 517192 3454
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 512430 -960 512542 326
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 518176 3602 518204 287710
rect 520280 249076 520332 249082
rect 520280 249018 520332 249024
rect 519544 3868 519596 3874
rect 519544 3810 519596 3816
rect 518164 3596 518216 3602
rect 518164 3538 518216 3544
rect 519556 480 519584 3810
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 249018
rect 520936 3534 520964 302903
rect 529940 301504 529992 301510
rect 529940 301446 529992 301452
rect 525800 294636 525852 294642
rect 525800 294578 525852 294584
rect 522304 283688 522356 283694
rect 522304 283630 522356 283636
rect 521844 3596 521896 3602
rect 521844 3538 521896 3544
rect 520924 3528 520976 3534
rect 520924 3470 520976 3476
rect 521856 480 521884 3538
rect 522316 3058 522344 283630
rect 525064 275324 525116 275330
rect 525064 275266 525116 275272
rect 524418 247616 524474 247625
rect 524418 247551 524474 247560
rect 524432 16574 524460 247551
rect 524432 16546 525012 16574
rect 523040 3528 523092 3534
rect 523040 3470 523092 3476
rect 524984 3482 525012 16546
rect 525076 3602 525104 275266
rect 525812 16574 525840 294578
rect 527824 293276 527876 293282
rect 527824 293218 527876 293224
rect 525812 16546 526208 16574
rect 525064 3596 525116 3602
rect 525064 3538 525116 3544
rect 522304 3052 522356 3058
rect 522304 2994 522356 3000
rect 523052 480 523080 3470
rect 524984 3454 525472 3482
rect 524236 3052 524288 3058
rect 524236 2994 524288 3000
rect 524248 480 524276 2994
rect 525444 480 525472 3454
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 520710 -960 520822 326
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527732 3596 527784 3602
rect 527732 3538 527784 3544
rect 527744 3346 527772 3538
rect 527836 3534 527864 293218
rect 528560 253224 528612 253230
rect 528560 253166 528612 253172
rect 527824 3528 527876 3534
rect 527824 3470 527876 3476
rect 527744 3318 527864 3346
rect 527836 480 527864 3318
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 253166
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 301446
rect 538864 300144 538916 300150
rect 538864 300086 538916 300092
rect 534724 291848 534776 291854
rect 534724 291790 534776 291796
rect 531320 283620 531372 283626
rect 531320 283562 531372 283568
rect 531332 3534 531360 283562
rect 531412 273964 531464 273970
rect 531412 273906 531464 273912
rect 531320 3528 531372 3534
rect 531320 3470 531372 3476
rect 531424 3346 531452 273906
rect 534080 244996 534132 245002
rect 534080 244938 534132 244944
rect 534092 16574 534120 244938
rect 534092 16546 534488 16574
rect 533712 3596 533764 3602
rect 533712 3538 533764 3544
rect 532148 3528 532200 3534
rect 532148 3470 532200 3476
rect 531332 3318 531452 3346
rect 531332 480 531360 3318
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532160 354 532188 3470
rect 533724 480 533752 3538
rect 532486 354 532598 480
rect 532160 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 534736 3194 534764 291790
rect 535460 265736 535512 265742
rect 535460 265678 535512 265684
rect 535472 16574 535500 265678
rect 538220 251932 538272 251938
rect 538220 251874 538272 251880
rect 535472 16546 536144 16574
rect 534724 3188 534776 3194
rect 534724 3130 534776 3136
rect 536116 480 536144 16546
rect 537208 3188 537260 3194
rect 537208 3130 537260 3136
rect 537220 480 537248 3130
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 251874
rect 538876 3058 538904 300086
rect 543004 290556 543056 290562
rect 543004 290498 543056 290504
rect 542360 260228 542412 260234
rect 542360 260170 542412 260176
rect 539692 258732 539744 258738
rect 539692 258674 539744 258680
rect 539704 6914 539732 258674
rect 540980 257440 541032 257446
rect 540980 257382 541032 257388
rect 540992 16574 541020 257382
rect 542372 16574 542400 260170
rect 540992 16546 542032 16574
rect 542372 16546 542768 16574
rect 539612 6886 539732 6914
rect 538864 3052 538916 3058
rect 538864 2994 538916 3000
rect 539612 480 539640 6886
rect 540796 3052 540848 3058
rect 540796 2994 540848 3000
rect 540808 480 540836 2994
rect 542004 480 542032 16546
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 543016 3398 543044 290498
rect 543752 16574 543780 307022
rect 570602 305688 570658 305697
rect 570602 305623 570658 305632
rect 545762 302832 545818 302841
rect 545762 302767 545818 302776
rect 545120 257372 545172 257378
rect 545120 257314 545172 257320
rect 545132 16574 545160 257314
rect 543752 16546 544424 16574
rect 545132 16546 545528 16574
rect 543004 3392 543056 3398
rect 543004 3334 543056 3340
rect 544396 480 544424 16546
rect 545500 480 545528 16546
rect 545776 3534 545804 302767
rect 547972 298852 548024 298858
rect 547972 298794 548024 298800
rect 547984 6914 548012 298794
rect 567844 298784 567896 298790
rect 567844 298726 567896 298732
rect 556160 297492 556212 297498
rect 556160 297434 556212 297440
rect 549904 290488 549956 290494
rect 549904 290430 549956 290436
rect 549260 267096 549312 267102
rect 549260 267038 549312 267044
rect 549272 16574 549300 267038
rect 549272 16546 549852 16574
rect 547892 6886 548012 6914
rect 545764 3528 545816 3534
rect 545764 3470 545816 3476
rect 546684 3528 546736 3534
rect 546684 3470 546736 3476
rect 546696 480 546724 3470
rect 547892 480 547920 6886
rect 549824 3482 549852 16546
rect 549916 3602 549944 290430
rect 552664 289128 552716 289134
rect 552664 289070 552716 289076
rect 552020 269816 552072 269822
rect 552020 269758 552072 269764
rect 552032 6914 552060 269758
rect 552676 16574 552704 289070
rect 553400 278044 553452 278050
rect 553400 277986 553452 277992
rect 553412 16574 553440 277986
rect 552676 16546 552796 16574
rect 553412 16546 553808 16574
rect 552032 6886 552704 6914
rect 549904 3596 549956 3602
rect 549904 3538 549956 3544
rect 551468 3596 551520 3602
rect 551468 3538 551520 3544
rect 549824 3454 550312 3482
rect 549076 3392 549128 3398
rect 549076 3334 549128 3340
rect 549088 480 549116 3334
rect 550284 480 550312 3454
rect 551480 480 551508 3538
rect 552676 480 552704 6886
rect 552768 2990 552796 16546
rect 552756 2984 552808 2990
rect 552756 2926 552808 2932
rect 553780 480 553808 16546
rect 556172 3534 556200 297434
rect 557540 297424 557592 297430
rect 557540 297366 557592 297372
rect 556252 282192 556304 282198
rect 556252 282134 556304 282140
rect 556160 3528 556212 3534
rect 556160 3470 556212 3476
rect 556264 3346 556292 282134
rect 557552 16574 557580 297366
rect 563704 295996 563756 296002
rect 563704 295938 563756 295944
rect 561680 287700 561732 287706
rect 561680 287642 561732 287648
rect 560944 265668 560996 265674
rect 560944 265610 560996 265616
rect 558920 260160 558972 260166
rect 558920 260102 558972 260108
rect 558932 16574 558960 260102
rect 560300 244928 560352 244934
rect 560300 244870 560352 244876
rect 560312 16574 560340 244870
rect 557552 16546 558592 16574
rect 558932 16546 559328 16574
rect 560312 16546 560432 16574
rect 556988 3528 557040 3534
rect 556988 3470 557040 3476
rect 556172 3318 556292 3346
rect 554964 2984 555016 2990
rect 554964 2926 555016 2932
rect 554976 480 555004 2926
rect 556172 480 556200 3318
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557000 354 557028 3470
rect 558564 480 558592 16546
rect 557326 354 557438 480
rect 557000 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 16546
rect 560956 3194 560984 265610
rect 561692 16574 561720 287642
rect 561692 16546 562088 16574
rect 560944 3188 560996 3194
rect 560944 3130 560996 3136
rect 562060 480 562088 16546
rect 563244 3188 563296 3194
rect 563244 3130 563296 3136
rect 563256 480 563284 3130
rect 563716 3058 563744 295938
rect 566464 286340 566516 286346
rect 566464 286282 566516 286288
rect 565820 267028 565872 267034
rect 565820 266970 565872 266976
rect 564532 254652 564584 254658
rect 564532 254594 564584 254600
rect 564544 6914 564572 254594
rect 565832 16574 565860 266970
rect 565832 16546 566412 16574
rect 564452 6886 564572 6914
rect 563704 3052 563756 3058
rect 563704 2994 563756 3000
rect 564452 480 564480 6886
rect 566384 3482 566412 16546
rect 566476 3874 566504 286282
rect 567200 254584 567252 254590
rect 567200 254526 567252 254532
rect 567212 16574 567240 254526
rect 567212 16546 567608 16574
rect 566464 3868 566516 3874
rect 566464 3810 566516 3816
rect 566384 3454 566872 3482
rect 565636 3052 565688 3058
rect 565636 2994 565688 3000
rect 565648 480 565676 2994
rect 566844 480 566872 3454
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 567856 3602 567884 298726
rect 569960 261520 570012 261526
rect 569960 261462 570012 261468
rect 569972 16574 570000 261462
rect 569972 16546 570368 16574
rect 569132 3868 569184 3874
rect 569132 3810 569184 3816
rect 567844 3596 567896 3602
rect 567844 3538 567896 3544
rect 569144 480 569172 3810
rect 570340 480 570368 16546
rect 570616 3534 570644 305623
rect 575480 284980 575532 284986
rect 575480 284922 575532 284928
rect 571984 280832 572036 280838
rect 571984 280774 572036 280780
rect 571524 3596 571576 3602
rect 571524 3538 571576 3544
rect 570604 3528 570656 3534
rect 570604 3470 570656 3476
rect 571536 480 571564 3538
rect 571996 3058 572024 280774
rect 574100 264240 574152 264246
rect 574100 264182 574152 264188
rect 574112 16574 574140 264182
rect 575492 16574 575520 284922
rect 576860 250504 576912 250510
rect 576860 250446 576912 250452
rect 576872 16574 576900 250446
rect 577516 33114 577544 441594
rect 577608 206990 577636 441730
rect 578240 251864 578292 251870
rect 578240 251806 578292 251812
rect 577596 206984 577648 206990
rect 577596 206926 577648 206932
rect 577504 33108 577556 33114
rect 577504 33050 577556 33056
rect 578252 16574 578280 251806
rect 578896 245585 578924 444382
rect 580538 443184 580594 443193
rect 580538 443119 580594 443128
rect 580262 443048 580318 443057
rect 580262 442983 580318 442992
rect 580080 442264 580132 442270
rect 580080 442206 580132 442212
rect 580092 431633 580120 442206
rect 580172 440904 580224 440910
rect 580172 440846 580224 440852
rect 580078 431624 580134 431633
rect 580078 431559 580134 431568
rect 579988 419484 580040 419490
rect 579988 419426 580040 419432
rect 580000 418305 580028 419426
rect 579986 418296 580042 418305
rect 579986 418231 580042 418240
rect 579804 405680 579856 405686
rect 579804 405622 579856 405628
rect 579816 404977 579844 405622
rect 579802 404968 579858 404977
rect 579802 404903 579858 404912
rect 580080 379500 580132 379506
rect 580080 379442 580132 379448
rect 580092 378457 580120 379442
rect 580078 378448 580134 378457
rect 580078 378383 580134 378392
rect 580080 365696 580132 365702
rect 580080 365638 580132 365644
rect 580092 365129 580120 365638
rect 580078 365120 580134 365129
rect 580078 365055 580134 365064
rect 580184 351937 580212 440846
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 580172 325644 580224 325650
rect 580172 325586 580224 325592
rect 580184 325281 580212 325586
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 579804 259412 579856 259418
rect 579804 259354 579856 259360
rect 579816 258913 579844 259354
rect 579802 258904 579858 258913
rect 579802 258839 579858 258848
rect 578882 245576 578938 245585
rect 578882 245511 578938 245520
rect 579620 206984 579672 206990
rect 579620 206926 579672 206932
rect 579632 205737 579660 206926
rect 579618 205728 579674 205737
rect 579618 205663 579674 205672
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 579620 167000 579672 167006
rect 579620 166942 579672 166948
rect 579632 165889 579660 166942
rect 579618 165880 579674 165889
rect 579618 165815 579674 165824
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 579618 33144 579674 33153
rect 579618 33079 579620 33088
rect 579672 33079 579674 33088
rect 579620 33050 579672 33056
rect 574112 16546 575152 16574
rect 575492 16546 575888 16574
rect 576872 16546 576992 16574
rect 578252 16546 578648 16574
rect 572720 3528 572772 3534
rect 572720 3470 572772 3476
rect 571984 3052 572036 3058
rect 571984 2994 572036 3000
rect 572732 480 572760 3470
rect 573916 3052 573968 3058
rect 573916 2994 573968 3000
rect 573928 480 573956 2994
rect 575124 480 575152 16546
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 567998 -960 568110 326
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 575860 354 575888 16546
rect 576278 354 576390 480
rect 575860 326 576390 354
rect 576964 354 576992 16546
rect 578620 480 578648 16546
rect 580276 6633 580304 442983
rect 580354 442232 580410 442241
rect 580354 442167 580410 442176
rect 580368 19825 580396 442167
rect 580448 441720 580500 441726
rect 580448 441662 580500 441668
rect 580460 112849 580488 441662
rect 580552 139369 580580 443119
rect 581092 443080 581144 443086
rect 581092 443022 581144 443028
rect 580816 442468 580868 442474
rect 580816 442410 580868 442416
rect 580632 442400 580684 442406
rect 580632 442342 580684 442348
rect 580644 152697 580672 442342
rect 580724 442332 580776 442338
rect 580724 442274 580776 442280
rect 580736 192545 580764 442274
rect 580828 272241 580856 442410
rect 580908 440972 580960 440978
rect 580908 440914 580960 440920
rect 580920 298761 580948 440914
rect 580906 298752 580962 298761
rect 580906 298687 580962 298696
rect 580814 272232 580870 272241
rect 580814 272167 580870 272176
rect 580722 192536 580778 192545
rect 580722 192471 580778 192480
rect 580630 152688 580686 152697
rect 580630 152623 580686 152632
rect 580538 139360 580594 139369
rect 580538 139295 580594 139304
rect 580446 112840 580502 112849
rect 580446 112775 580502 112784
rect 580354 19816 580410 19825
rect 580354 19751 580410 19760
rect 581104 16574 581132 443022
rect 582380 443012 582432 443018
rect 582380 442954 582432 442960
rect 582392 16574 582420 442954
rect 581104 16546 581776 16574
rect 582392 16546 583432 16574
rect 580262 6624 580318 6633
rect 580262 6559 580318 6568
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 581012 480 581040 3402
rect 577382 354 577494 480
rect 576964 326 577494 354
rect 576278 -960 576390 326
rect 577382 -960 577494 326
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 581748 354 581776 16546
rect 583404 480 583432 16546
rect 582166 354 582278 480
rect 581748 326 582278 354
rect 582166 -960 582278 326
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 2778 632068 2780 632088
rect 2780 632068 2832 632088
rect 2832 632068 2834 632088
rect 2778 632032 2834 632068
rect 3146 619112 3202 619168
rect 3422 606076 3478 606112
rect 3422 606056 3424 606076
rect 3424 606056 3476 606076
rect 3476 606056 3478 606076
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3422 553832 3478 553888
rect 3422 527856 3478 527912
rect 3422 514820 3478 514856
rect 3422 514800 3424 514820
rect 3424 514800 3476 514820
rect 3476 514800 3478 514820
rect 3054 501744 3110 501800
rect 3422 475632 3478 475688
rect 3238 462576 3294 462632
rect 217598 516840 217654 516896
rect 217506 513712 217562 513768
rect 217414 489912 217470 489968
rect 217322 488008 217378 488064
rect 4066 449520 4122 449576
rect 217690 515888 217746 515944
rect 3330 423580 3332 423600
rect 3332 423580 3384 423600
rect 3384 423580 3386 423600
rect 3330 423544 3386 423580
rect 2962 410488 3018 410544
rect 3054 397432 3110 397488
rect 3146 371320 3202 371376
rect 2962 319232 3018 319288
rect 3330 306176 3386 306232
rect 2962 267144 3018 267200
rect 3330 254088 3386 254144
rect 3054 201864 3110 201920
rect 3790 358400 3846 358456
rect 3698 345344 3754 345400
rect 3606 293120 3662 293176
rect 3514 241032 3570 241088
rect 3514 188808 3570 188864
rect 3514 149776 3570 149832
rect 3514 136720 3570 136776
rect 3422 110608 3478 110664
rect 3422 97552 3478 97608
rect 3146 84632 3202 84688
rect 3422 71576 3478 71632
rect 3054 58520 3110 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 20718 300056 20774 300112
rect 95882 440272 95938 440328
rect 97722 364656 97778 364712
rect 97630 361936 97686 361992
rect 97906 367376 97962 367432
rect 97906 356496 97962 356552
rect 97814 351056 97870 351112
rect 97814 348336 97870 348392
rect 97722 345616 97778 345672
rect 97630 340176 97686 340232
rect 97538 334736 97594 334792
rect 97446 332016 97502 332072
rect 97354 326576 97410 326632
rect 97446 299376 97502 299432
rect 155866 373224 155922 373280
rect 159914 374040 159970 374096
rect 124678 371612 124734 371648
rect 124678 371592 124680 371612
rect 124680 371592 124732 371612
rect 124732 371592 124734 371612
rect 135074 371592 135130 371648
rect 137926 371612 137982 371648
rect 137926 371592 137928 371612
rect 137928 371592 137980 371612
rect 137980 371592 137982 371612
rect 144182 371612 144238 371648
rect 144182 371592 144184 371612
rect 144184 371592 144236 371612
rect 144236 371592 144238 371612
rect 99838 370640 99894 370696
rect 99286 359216 99342 359272
rect 99194 353776 99250 353832
rect 99102 337456 99158 337512
rect 99010 329296 99066 329352
rect 98918 323856 98974 323912
rect 98826 318416 98882 318472
rect 98734 315696 98790 315752
rect 98642 310256 98698 310312
rect 97906 304816 97962 304872
rect 97538 299240 97594 299296
rect 97262 299104 97318 299160
rect 99378 342896 99434 342952
rect 99286 300736 99342 300792
rect 99470 321136 99526 321192
rect 99562 312976 99618 313032
rect 99838 307536 99894 307592
rect 99746 301552 99802 301608
rect 170586 309304 170642 309360
rect 171690 358536 171746 358592
rect 171138 350376 171194 350432
rect 170954 309440 171010 309496
rect 170770 309168 170826 309224
rect 164238 300328 164294 300384
rect 160098 300192 160154 300248
rect 101954 298016 102010 298072
rect 145746 297880 145802 297936
rect 170494 303048 170550 303104
rect 171322 323176 171378 323232
rect 171506 320456 171562 320512
rect 171506 317736 171562 317792
rect 172334 369416 172390 369472
rect 172426 366696 172482 366752
rect 172334 363976 172390 364032
rect 171874 361256 171930 361312
rect 171966 355816 172022 355872
rect 172426 353096 172482 353152
rect 172426 347656 172482 347712
rect 172058 344936 172114 344992
rect 172150 342216 172206 342272
rect 172058 310800 172114 310856
rect 172242 339496 172298 339552
rect 172426 336796 172482 336832
rect 172426 336776 172428 336796
rect 172428 336776 172480 336796
rect 172480 336776 172482 336796
rect 172426 334056 172482 334112
rect 172426 331336 172482 331392
rect 172334 328616 172390 328672
rect 172426 325896 172482 325952
rect 172426 315016 172482 315072
rect 172426 312296 172482 312352
rect 172242 309576 172298 309632
rect 173438 308896 173494 308952
rect 173254 308216 173310 308272
rect 171414 306856 171470 306912
rect 172334 304136 172390 304192
rect 172426 301416 172482 301472
rect 184938 302912 184994 302968
rect 182178 302776 182234 302832
rect 219070 512760 219126 512816
rect 218978 508136 219034 508192
rect 218886 488280 218942 488336
rect 219162 510992 219218 511048
rect 219254 509904 219310 509960
rect 238482 477264 238538 477320
rect 242806 477128 242862 477184
rect 253754 477128 253810 477184
rect 240046 476856 240102 476912
rect 241426 476876 241482 476912
rect 241426 476856 241428 476876
rect 241428 476856 241480 476876
rect 241480 476856 241482 476876
rect 237286 476740 237342 476776
rect 237286 476720 237288 476740
rect 237288 476720 237340 476740
rect 237340 476720 237342 476740
rect 237194 476176 237250 476232
rect 245566 476312 245622 476368
rect 248234 476312 248290 476368
rect 251086 476312 251142 476368
rect 252374 476312 252430 476368
rect 244186 476176 244242 476232
rect 245474 476176 245530 476232
rect 246946 476176 247002 476232
rect 248326 476176 248382 476232
rect 249706 476176 249762 476232
rect 250994 476176 251050 476232
rect 252466 476176 252522 476232
rect 243726 445848 243782 445904
rect 205086 3304 205142 3360
rect 214838 308352 214894 308408
rect 210790 155216 210846 155272
rect 211986 300464 212042 300520
rect 212078 297336 212134 297392
rect 213366 297608 213422 297664
rect 213550 297472 213606 297528
rect 214654 157800 214710 157856
rect 214470 3440 214526 3496
rect 215666 3440 215722 3496
rect 215206 3304 215262 3360
rect 217138 192752 217194 192808
rect 216678 188128 216734 188184
rect 217322 195880 217378 195936
rect 217230 168000 217286 168056
rect 217414 168272 217470 168328
rect 217690 196832 217746 196888
rect 217782 193704 217838 193760
rect 217598 169904 217654 169960
rect 218426 190984 218482 191040
rect 218610 193160 218666 193216
rect 218518 189896 218574 189952
rect 234618 444624 234674 444680
rect 232686 442992 232742 443048
rect 235262 443264 235318 443320
rect 237838 445712 237894 445768
rect 236550 444352 236606 444408
rect 238574 444488 238630 444544
rect 239862 443128 239918 443184
rect 243082 441632 243138 441688
rect 246946 442176 247002 442232
rect 256606 476992 256662 477048
rect 253846 476176 253902 476232
rect 255226 476176 255282 476232
rect 256514 476176 256570 476232
rect 259366 476720 259422 476776
rect 257986 476176 258042 476232
rect 259274 476176 259330 476232
rect 266266 476584 266322 476640
rect 262126 476448 262182 476504
rect 260654 476312 260710 476368
rect 264794 476312 264850 476368
rect 267646 476312 267702 476368
rect 260746 476176 260802 476232
rect 262034 476176 262090 476232
rect 263506 476176 263562 476232
rect 264886 476176 264942 476232
rect 266174 476176 266230 476232
rect 267554 476176 267610 476232
rect 268934 476312 268990 476368
rect 269026 476176 269082 476232
rect 270406 476176 270462 476232
rect 271786 476604 271842 476640
rect 271786 476584 271788 476604
rect 271788 476584 271840 476604
rect 271840 476584 271842 476604
rect 274546 476448 274602 476504
rect 274454 476312 274510 476368
rect 271694 476176 271750 476232
rect 273166 476176 273222 476232
rect 274362 476176 274418 476232
rect 277306 476312 277362 476368
rect 278594 476312 278650 476368
rect 275926 476176 275982 476232
rect 277214 476176 277270 476232
rect 278686 476176 278742 476232
rect 280066 476176 280122 476232
rect 281446 476176 281502 476232
rect 284206 476176 284262 476232
rect 286506 476176 286562 476232
rect 288346 476176 288402 476232
rect 291106 476176 291162 476232
rect 293866 476176 293922 476232
rect 296626 476176 296682 476232
rect 299386 476176 299442 476232
rect 302146 476176 302202 476232
rect 303526 476176 303582 476232
rect 306286 476176 306342 476232
rect 297454 444896 297510 444952
rect 299386 444760 299442 444816
rect 306010 441768 306066 441824
rect 309046 476720 309102 476776
rect 311806 476312 311862 476368
rect 321466 476992 321522 477048
rect 314566 476720 314622 476776
rect 315946 476196 316002 476232
rect 315946 476176 315948 476196
rect 315948 476176 316000 476196
rect 316000 476176 316002 476196
rect 318706 476468 318762 476504
rect 318706 476448 318708 476468
rect 318708 476448 318760 476468
rect 318760 476448 318762 476468
rect 324226 476448 324282 476504
rect 326986 476448 327042 476504
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580262 630808 580318 630864
rect 580170 617480 580226 617536
rect 580170 590960 580226 591016
rect 579894 564304 579950 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 580170 471416 580226 471472
rect 580170 458088 580226 458144
rect 580354 577632 580410 577688
rect 289818 441224 289874 441280
rect 290738 441124 290740 441144
rect 290740 441124 290792 441144
rect 290792 441124 290794 441144
rect 290738 441088 290794 441124
rect 293774 441224 293830 441280
rect 293682 441088 293738 441144
rect 304998 440952 305054 441008
rect 225786 310528 225842 310584
rect 228546 309576 228602 309632
rect 228638 308624 228694 308680
rect 231214 309848 231270 309904
rect 231306 309032 231362 309088
rect 231490 308760 231546 308816
rect 232226 311244 232228 311264
rect 232228 311244 232280 311264
rect 232280 311244 232282 311264
rect 232226 311208 232282 311244
rect 233698 310528 233754 310584
rect 234066 310528 234122 310584
rect 232410 310392 232466 310448
rect 232870 310256 232926 310312
rect 234526 308896 234582 308952
rect 234342 299240 234398 299296
rect 235722 309032 235778 309088
rect 236274 301552 236330 301608
rect 237562 299376 237618 299432
rect 240322 309848 240378 309904
rect 241242 309984 241298 310040
rect 244646 309304 244702 309360
rect 245658 300736 245714 300792
rect 247314 309712 247370 309768
rect 248142 309576 248198 309632
rect 248326 308760 248382 308816
rect 248602 301144 248658 301200
rect 250350 308216 250406 308272
rect 250994 308488 251050 308544
rect 251730 309168 251786 309224
rect 252650 308624 252706 308680
rect 255778 300056 255834 300112
rect 260102 303048 260158 303104
rect 278594 300192 278650 300248
rect 279330 300328 279386 300384
rect 282090 302776 282146 302832
rect 282642 302912 282698 302968
rect 285954 284824 286010 284880
rect 288346 306176 288402 306232
rect 287610 303320 287666 303376
rect 287518 303184 287574 303240
rect 288714 305904 288770 305960
rect 288898 306040 288954 306096
rect 290094 305768 290150 305824
rect 290002 300464 290058 300520
rect 290186 297608 290242 297664
rect 291566 297472 291622 297528
rect 290278 297336 290334 297392
rect 291750 305632 291806 305688
rect 293314 297744 293370 297800
rect 287150 255856 287206 255912
rect 287058 250416 287114 250472
rect 298282 308352 298338 308408
rect 298098 305904 298154 305960
rect 298834 303320 298890 303376
rect 299754 300056 299810 300112
rect 303986 250824 304042 250880
rect 303802 250416 303858 250472
rect 305274 248104 305330 248160
rect 308402 250688 308458 250744
rect 308218 250552 308274 250608
rect 308126 247696 308182 247752
rect 309230 247968 309286 248024
rect 309138 245520 309194 245576
rect 309414 247832 309470 247888
rect 309322 245384 309378 245440
rect 306470 245248 306526 245304
rect 305366 245112 305422 245168
rect 305182 244976 305238 245032
rect 304998 244840 305054 244896
rect 311070 308488 311126 308544
rect 310794 253136 310850 253192
rect 311070 258712 311126 258768
rect 310978 254632 311034 254688
rect 310886 251912 310942 251968
rect 310702 251776 310758 251832
rect 312358 303456 312414 303512
rect 312082 286320 312138 286376
rect 315394 305768 315450 305824
rect 313278 254496 313334 254552
rect 318246 303184 318302 303240
rect 319350 306040 319406 306096
rect 310610 248240 310666 248296
rect 329930 308352 329986 308408
rect 331678 303048 331734 303104
rect 337290 302912 337346 302968
rect 336738 247560 336794 247616
rect 341706 302776 341762 302832
rect 345110 305632 345166 305688
rect 346950 309032 347006 309088
rect 346766 308216 346822 308272
rect 347502 308896 347558 308952
rect 348422 308760 348478 308816
rect 349250 308624 349306 308680
rect 349986 306176 350042 306232
rect 350998 306312 351054 306368
rect 310518 244704 310574 244760
rect 303618 243616 303674 243672
rect 298650 243480 298706 243536
rect 258538 159840 258594 159896
rect 275834 159840 275890 159896
rect 277030 159840 277086 159896
rect 278134 159840 278190 159896
rect 279238 159840 279294 159896
rect 255962 159568 256018 159624
rect 220818 158616 220874 158672
rect 238114 158652 238116 158672
rect 238116 158652 238168 158672
rect 238168 158652 238170 158672
rect 219438 158208 219494 158264
rect 238114 158616 238170 158652
rect 239586 158616 239642 158672
rect 240690 158616 240746 158672
rect 248326 158616 248382 158672
rect 250166 158616 250222 158672
rect 224958 158480 225014 158536
rect 223578 157800 223634 157856
rect 216862 3440 216918 3496
rect 219254 3440 219310 3496
rect 222750 3304 222806 3360
rect 227718 158344 227774 158400
rect 231858 158072 231914 158128
rect 238758 157936 238814 157992
rect 245382 158208 245438 158264
rect 246854 158072 246910 158128
rect 246854 155896 246910 155952
rect 248694 157936 248750 157992
rect 248694 155760 248750 155816
rect 252374 158480 252430 158536
rect 252098 157936 252154 157992
rect 252374 156712 252430 156768
rect 251270 155352 251326 155408
rect 253570 157936 253626 157992
rect 253202 157256 253258 157312
rect 253202 156848 253258 156904
rect 253662 157392 253718 157448
rect 256606 158616 256662 158672
rect 271050 159568 271106 159624
rect 274454 159568 274510 159624
rect 257158 158616 257214 158672
rect 258630 158616 258686 158672
rect 259550 158616 259606 158672
rect 260654 158480 260710 158536
rect 261758 158616 261814 158672
rect 262862 158616 262918 158672
rect 261942 157936 261998 157992
rect 264426 157664 264482 157720
rect 263966 157392 264022 157448
rect 265990 158616 266046 158672
rect 267646 158616 267702 158672
rect 268750 158616 268806 158672
rect 270222 158616 270278 158672
rect 266726 157936 266782 157992
rect 268934 157936 268990 157992
rect 265990 157664 266046 157720
rect 300950 159704 301006 159760
rect 271142 158616 271198 158672
rect 272246 158616 272302 158672
rect 276110 158480 276166 158536
rect 281354 158480 281410 158536
rect 273350 158344 273406 158400
rect 274454 157664 274510 157720
rect 269118 155216 269174 155272
rect 278686 157664 278742 157720
rect 296718 159296 296774 159352
rect 286230 158480 286286 158536
rect 284114 157664 284170 157720
rect 291014 158344 291070 158400
rect 296258 158344 296314 158400
rect 288254 157528 288310 157584
rect 293590 157528 293646 157584
rect 292578 155352 292634 155408
rect 291198 155216 291254 155272
rect 293958 155488 294014 155544
rect 298926 158616 298982 158672
rect 303526 158616 303582 158672
rect 306102 158636 306158 158672
rect 306102 158616 306104 158636
rect 306104 158616 306156 158636
rect 306156 158616 306158 158636
rect 308678 158652 308680 158672
rect 308680 158652 308732 158672
rect 308732 158652 308734 158672
rect 308678 158616 308734 158652
rect 313462 158616 313518 158672
rect 311254 158208 311310 158264
rect 315854 158616 315910 158672
rect 318614 158616 318670 158672
rect 321190 158616 321246 158672
rect 323398 158616 323454 158672
rect 325974 158616 326030 158672
rect 353942 158480 353998 158536
rect 348422 158208 348478 158264
rect 345662 157936 345718 157992
rect 323306 6296 323362 6352
rect 320914 6160 320970 6216
rect 325606 3440 325662 3496
rect 324410 3304 324466 3360
rect 327998 3576 328054 3632
rect 344558 6432 344614 6488
rect 331586 3712 331642 3768
rect 335082 3848 335138 3904
rect 343362 3984 343418 4040
rect 348054 6568 348110 6624
rect 346950 3168 347006 3224
rect 351182 158072 351238 158128
rect 350446 6840 350502 6896
rect 351642 6704 351698 6760
rect 354126 158344 354182 158400
rect 356426 3984 356482 4040
rect 356610 3984 356666 4040
rect 356886 243480 356942 243536
rect 357346 159432 357402 159488
rect 357346 158752 357402 158808
rect 358266 305904 358322 305960
rect 358082 158752 358138 158808
rect 356610 3712 356666 3768
rect 356702 3576 356758 3632
rect 357530 3576 357586 3632
rect 356702 3168 356758 3224
rect 356426 2896 356482 2952
rect 358266 158480 358322 158536
rect 359646 243616 359702 243672
rect 359646 157936 359702 157992
rect 362130 308216 362186 308272
rect 361118 158752 361174 158808
rect 358726 3440 358782 3496
rect 359922 3440 359978 3496
rect 361118 3440 361174 3496
rect 366454 309032 366510 309088
rect 362130 159432 362186 159488
rect 362406 158208 362462 158264
rect 362314 155488 362370 155544
rect 363418 243752 363474 243808
rect 363786 158344 363842 158400
rect 363510 3440 363566 3496
rect 363142 2896 363198 2952
rect 365074 159160 365130 159216
rect 365258 158752 365314 158808
rect 365166 158072 365222 158128
rect 365810 6704 365866 6760
rect 366270 308896 366326 308952
rect 367098 303320 367154 303376
rect 366454 158888 366510 158944
rect 366270 157800 366326 157856
rect 365810 3576 365866 3632
rect 364614 3440 364670 3496
rect 367006 3440 367062 3496
rect 368570 308760 368626 308816
rect 367926 155216 367982 155272
rect 370042 308624 370098 308680
rect 369030 306176 369086 306232
rect 368570 157120 368626 157176
rect 369030 156984 369086 157040
rect 369306 159296 369362 159352
rect 370134 306312 370190 306368
rect 370042 155896 370098 155952
rect 370134 155760 370190 155816
rect 370318 156848 370374 156904
rect 371330 308488 371386 308544
rect 368202 3440 368258 3496
rect 370594 3440 370650 3496
rect 372066 159024 372122 159080
rect 373170 157256 373226 157312
rect 377402 306040 377458 306096
rect 385038 305768 385094 305824
rect 379978 3304 380034 3360
rect 462962 308352 463018 308408
rect 396722 303184 396778 303240
rect 489182 303048 489238 303104
rect 520922 302912 520978 302968
rect 524418 247560 524474 247616
rect 570602 305632 570658 305688
rect 545762 302776 545818 302832
rect 580538 443128 580594 443184
rect 580262 442992 580318 443048
rect 580078 431568 580134 431624
rect 579986 418240 580042 418296
rect 579802 404912 579858 404968
rect 580078 378392 580134 378448
rect 580078 365064 580134 365120
rect 580170 351872 580226 351928
rect 580170 325216 580226 325272
rect 580170 312024 580226 312080
rect 579802 258848 579858 258904
rect 578882 245520 578938 245576
rect 579618 205672 579674 205728
rect 580170 179152 580226 179208
rect 579618 165824 579674 165880
rect 580170 59608 580226 59664
rect 579618 33108 579674 33144
rect 579618 33088 579620 33108
rect 579620 33088 579672 33108
rect 579672 33088 579674 33108
rect 580354 442176 580410 442232
rect 580906 298696 580962 298752
rect 580814 272176 580870 272232
rect 580722 192480 580778 192536
rect 580630 152632 580686 152688
rect 580538 139304 580594 139360
rect 580446 112784 580502 112840
rect 580354 19760 580410 19816
rect 580262 6568 580318 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 2773 632090 2839 632093
rect -960 632088 2839 632090
rect -960 632032 2778 632088
rect 2834 632032 2839 632088
rect -960 632030 2839 632032
rect -960 631940 480 632030
rect 2773 632027 2839 632030
rect 580257 630866 580323 630869
rect 583520 630866 584960 630956
rect 580257 630864 584960 630866
rect 580257 630808 580262 630864
rect 580318 630808 584960 630864
rect 580257 630806 584960 630808
rect 580257 630803 580323 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3417 606114 3483 606117
rect -960 606112 3483 606114
rect -960 606056 3422 606112
rect 3478 606056 3483 606112
rect -960 606054 3483 606056
rect -960 605964 480 606054
rect 3417 606051 3483 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580349 577690 580415 577693
rect 583520 577690 584960 577780
rect 580349 577688 584960 577690
rect 580349 577632 580354 577688
rect 580410 577632 584960 577688
rect 580349 577630 584960 577632
rect 580349 577627 580415 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 579889 564362 579955 564365
rect 583520 564362 584960 564452
rect 579889 564360 584960 564362
rect 579889 564304 579894 564360
rect 579950 564304 584960 564360
rect 579889 564302 584960 564304
rect 579889 564299 579955 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect 217593 516898 217659 516901
rect 219390 516898 220064 516924
rect 217593 516896 220064 516898
rect 217593 516840 217598 516896
rect 217654 516864 220064 516896
rect 217654 516840 219450 516864
rect 217593 516838 219450 516840
rect 217593 516835 217659 516838
rect 217685 515946 217751 515949
rect 219390 515946 220064 515972
rect 217685 515944 220064 515946
rect 217685 515888 217690 515944
rect 217746 515912 220064 515944
rect 217746 515888 219450 515912
rect 217685 515886 219450 515888
rect 217685 515883 217751 515886
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 217501 513770 217567 513773
rect 219390 513770 220064 513796
rect 217501 513768 220064 513770
rect 217501 513712 217506 513768
rect 217562 513736 220064 513768
rect 217562 513712 219450 513736
rect 217501 513710 219450 513712
rect 217501 513707 217567 513710
rect 219065 512818 219131 512821
rect 219390 512818 220064 512844
rect 219065 512816 220064 512818
rect 219065 512760 219070 512816
rect 219126 512784 220064 512816
rect 219126 512760 219450 512784
rect 219065 512758 219450 512760
rect 219065 512755 219131 512758
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect 219157 511050 219223 511053
rect 219390 511050 220064 511076
rect 219157 511048 220064 511050
rect 219157 510992 219162 511048
rect 219218 511016 220064 511048
rect 219218 510992 219450 511016
rect 219157 510990 219450 510992
rect 219157 510987 219223 510990
rect 219249 509962 219315 509965
rect 219390 509962 220064 509988
rect 219249 509960 220064 509962
rect 219249 509904 219254 509960
rect 219310 509928 220064 509960
rect 219310 509904 219450 509928
rect 219249 509902 219450 509904
rect 219249 509899 219315 509902
rect 218973 508194 219039 508197
rect 219390 508194 220064 508220
rect 218973 508192 220064 508194
rect 218973 508136 218978 508192
rect 219034 508160 220064 508192
rect 219034 508136 219450 508160
rect 218973 508134 219450 508136
rect 218973 508131 219039 508134
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 583520 497844 584960 498084
rect 217409 489970 217475 489973
rect 219390 489970 220064 489996
rect 217409 489968 220064 489970
rect 217409 489912 217414 489968
rect 217470 489936 220064 489968
rect 217470 489912 219450 489936
rect 217409 489910 219450 489912
rect 217409 489907 217475 489910
rect -960 488596 480 488836
rect 218881 488338 218947 488341
rect 219390 488338 220064 488364
rect 218881 488336 220064 488338
rect 218881 488280 218886 488336
rect 218942 488304 220064 488336
rect 218942 488280 219450 488304
rect 218881 488278 219450 488280
rect 218881 488275 218947 488278
rect 217317 488066 217383 488069
rect 219390 488066 220064 488092
rect 217317 488064 220064 488066
rect 217317 488008 217322 488064
rect 217378 488032 220064 488064
rect 217378 488008 219450 488032
rect 217317 488006 219450 488008
rect 217317 488003 217383 488006
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect 238334 477260 238340 477324
rect 238404 477322 238410 477324
rect 238477 477322 238543 477325
rect 238404 477320 238543 477322
rect 238404 477264 238482 477320
rect 238538 477264 238543 477320
rect 238404 477262 238543 477264
rect 238404 477260 238410 477262
rect 238477 477259 238543 477262
rect 241830 477124 241836 477188
rect 241900 477186 241906 477188
rect 242801 477186 242867 477189
rect 241900 477184 242867 477186
rect 241900 477128 242806 477184
rect 242862 477128 242867 477184
rect 241900 477126 242867 477128
rect 241900 477124 241906 477126
rect 242801 477123 242867 477126
rect 253422 477124 253428 477188
rect 253492 477186 253498 477188
rect 253749 477186 253815 477189
rect 253492 477184 253815 477186
rect 253492 477128 253754 477184
rect 253810 477128 253815 477184
rect 253492 477126 253815 477128
rect 253492 477124 253498 477126
rect 253749 477123 253815 477126
rect 256182 476988 256188 477052
rect 256252 477050 256258 477052
rect 256601 477050 256667 477053
rect 256252 477048 256667 477050
rect 256252 476992 256606 477048
rect 256662 476992 256667 477048
rect 256252 476990 256667 476992
rect 256252 476988 256258 476990
rect 256601 476987 256667 476990
rect 320950 476988 320956 477052
rect 321020 477050 321026 477052
rect 321461 477050 321527 477053
rect 321020 477048 321527 477050
rect 321020 476992 321466 477048
rect 321522 476992 321527 477048
rect 321020 476990 321527 476992
rect 321020 476988 321026 476990
rect 321461 476987 321527 476990
rect 239622 476852 239628 476916
rect 239692 476914 239698 476916
rect 240041 476914 240107 476917
rect 239692 476912 240107 476914
rect 239692 476856 240046 476912
rect 240102 476856 240107 476912
rect 239692 476854 240107 476856
rect 239692 476852 239698 476854
rect 240041 476851 240107 476854
rect 240542 476852 240548 476916
rect 240612 476914 240618 476916
rect 241421 476914 241487 476917
rect 240612 476912 241487 476914
rect 240612 476856 241426 476912
rect 241482 476856 241487 476912
rect 240612 476854 241487 476856
rect 240612 476852 240618 476854
rect 241421 476851 241487 476854
rect 236126 476716 236132 476780
rect 236196 476778 236202 476780
rect 237281 476778 237347 476781
rect 236196 476776 237347 476778
rect 236196 476720 237286 476776
rect 237342 476720 237347 476776
rect 236196 476718 237347 476720
rect 236196 476716 236202 476718
rect 237281 476715 237347 476718
rect 258022 476716 258028 476780
rect 258092 476778 258098 476780
rect 259361 476778 259427 476781
rect 258092 476776 259427 476778
rect 258092 476720 259366 476776
rect 259422 476720 259427 476776
rect 258092 476718 259427 476720
rect 258092 476716 258098 476718
rect 259361 476715 259427 476718
rect 308622 476716 308628 476780
rect 308692 476778 308698 476780
rect 309041 476778 309107 476781
rect 308692 476776 309107 476778
rect 308692 476720 309046 476776
rect 309102 476720 309107 476776
rect 308692 476718 309107 476720
rect 308692 476716 308698 476718
rect 309041 476715 309107 476718
rect 313406 476716 313412 476780
rect 313476 476778 313482 476780
rect 314561 476778 314627 476781
rect 313476 476776 314627 476778
rect 313476 476720 314566 476776
rect 314622 476720 314627 476776
rect 313476 476718 314627 476720
rect 313476 476716 313482 476718
rect 314561 476715 314627 476718
rect 265934 476580 265940 476644
rect 266004 476642 266010 476644
rect 266261 476642 266327 476645
rect 266004 476640 266327 476642
rect 266004 476584 266266 476640
rect 266322 476584 266327 476640
rect 266004 476582 266327 476584
rect 266004 476580 266010 476582
rect 266261 476579 266327 476582
rect 270902 476580 270908 476644
rect 270972 476642 270978 476644
rect 271781 476642 271847 476645
rect 270972 476640 271847 476642
rect 270972 476584 271786 476640
rect 271842 476584 271847 476640
rect 270972 476582 271847 476584
rect 270972 476580 270978 476582
rect 271781 476579 271847 476582
rect 261150 476444 261156 476508
rect 261220 476506 261226 476508
rect 262121 476506 262187 476509
rect 261220 476504 262187 476506
rect 261220 476448 262126 476504
rect 262182 476448 262187 476504
rect 261220 476446 262187 476448
rect 261220 476444 261226 476446
rect 262121 476443 262187 476446
rect 273662 476444 273668 476508
rect 273732 476506 273738 476508
rect 274541 476506 274607 476509
rect 273732 476504 274607 476506
rect 273732 476448 274546 476504
rect 274602 476448 274607 476504
rect 273732 476446 274607 476448
rect 273732 476444 273738 476446
rect 274541 476443 274607 476446
rect 318558 476444 318564 476508
rect 318628 476506 318634 476508
rect 318701 476506 318767 476509
rect 318628 476504 318767 476506
rect 318628 476448 318706 476504
rect 318762 476448 318767 476504
rect 318628 476446 318767 476448
rect 318628 476444 318634 476446
rect 318701 476443 318767 476446
rect 323342 476444 323348 476508
rect 323412 476506 323418 476508
rect 324221 476506 324287 476509
rect 323412 476504 324287 476506
rect 323412 476448 324226 476504
rect 324282 476448 324287 476504
rect 323412 476446 324287 476448
rect 323412 476444 323418 476446
rect 324221 476443 324287 476446
rect 325918 476444 325924 476508
rect 325988 476506 325994 476508
rect 326981 476506 327047 476509
rect 325988 476504 327047 476506
rect 325988 476448 326986 476504
rect 327042 476448 327047 476504
rect 325988 476446 327047 476448
rect 325988 476444 325994 476446
rect 326981 476443 327047 476446
rect 244222 476308 244228 476372
rect 244292 476370 244298 476372
rect 245561 476370 245627 476373
rect 244292 476368 245627 476370
rect 244292 476312 245566 476368
rect 245622 476312 245627 476368
rect 244292 476310 245627 476312
rect 244292 476308 244298 476310
rect 245561 476307 245627 476310
rect 247718 476308 247724 476372
rect 247788 476370 247794 476372
rect 248229 476370 248295 476373
rect 247788 476368 248295 476370
rect 247788 476312 248234 476368
rect 248290 476312 248295 476368
rect 247788 476310 248295 476312
rect 247788 476308 247794 476310
rect 248229 476307 248295 476310
rect 250110 476308 250116 476372
rect 250180 476370 250186 476372
rect 251081 476370 251147 476373
rect 250180 476368 251147 476370
rect 250180 476312 251086 476368
rect 251142 476312 251147 476368
rect 250180 476310 251147 476312
rect 250180 476308 250186 476310
rect 251081 476307 251147 476310
rect 251398 476308 251404 476372
rect 251468 476370 251474 476372
rect 252369 476370 252435 476373
rect 251468 476368 252435 476370
rect 251468 476312 252374 476368
rect 252430 476312 252435 476368
rect 251468 476310 252435 476312
rect 251468 476308 251474 476310
rect 252369 476307 252435 476310
rect 259494 476308 259500 476372
rect 259564 476370 259570 476372
rect 260649 476370 260715 476373
rect 259564 476368 260715 476370
rect 259564 476312 260654 476368
rect 260710 476312 260715 476368
rect 259564 476310 260715 476312
rect 259564 476308 259570 476310
rect 260649 476307 260715 476310
rect 263542 476308 263548 476372
rect 263612 476370 263618 476372
rect 264789 476370 264855 476373
rect 263612 476368 264855 476370
rect 263612 476312 264794 476368
rect 264850 476312 264855 476368
rect 263612 476310 264855 476312
rect 263612 476308 263618 476310
rect 264789 476307 264855 476310
rect 266486 476308 266492 476372
rect 266556 476370 266562 476372
rect 267641 476370 267707 476373
rect 266556 476368 267707 476370
rect 266556 476312 267646 476368
rect 267702 476312 267707 476368
rect 266556 476310 267707 476312
rect 266556 476308 266562 476310
rect 267641 476307 267707 476310
rect 268326 476308 268332 476372
rect 268396 476370 268402 476372
rect 268929 476370 268995 476373
rect 268396 476368 268995 476370
rect 268396 476312 268934 476368
rect 268990 476312 268995 476368
rect 268396 476310 268995 476312
rect 268396 476308 268402 476310
rect 268929 476307 268995 476310
rect 273294 476308 273300 476372
rect 273364 476370 273370 476372
rect 274449 476370 274515 476373
rect 273364 476368 274515 476370
rect 273364 476312 274454 476368
rect 274510 476312 274515 476368
rect 273364 476310 274515 476312
rect 273364 476308 273370 476310
rect 274449 476307 274515 476310
rect 276054 476308 276060 476372
rect 276124 476370 276130 476372
rect 277301 476370 277367 476373
rect 276124 476368 277367 476370
rect 276124 476312 277306 476368
rect 277362 476312 277367 476368
rect 276124 476310 277367 476312
rect 276124 476308 276130 476310
rect 277301 476307 277367 476310
rect 278078 476308 278084 476372
rect 278148 476370 278154 476372
rect 278589 476370 278655 476373
rect 278148 476368 278655 476370
rect 278148 476312 278594 476368
rect 278650 476312 278655 476368
rect 278148 476310 278655 476312
rect 278148 476308 278154 476310
rect 278589 476307 278655 476310
rect 311014 476308 311020 476372
rect 311084 476370 311090 476372
rect 311801 476370 311867 476373
rect 311084 476368 311867 476370
rect 311084 476312 311806 476368
rect 311862 476312 311867 476368
rect 311084 476310 311867 476312
rect 311084 476308 311090 476310
rect 311801 476307 311867 476310
rect 237189 476236 237255 476237
rect 237189 476234 237236 476236
rect 237144 476232 237236 476234
rect 237144 476176 237194 476232
rect 237144 476174 237236 476176
rect 237189 476172 237236 476174
rect 237300 476172 237306 476236
rect 243118 476172 243124 476236
rect 243188 476234 243194 476236
rect 244181 476234 244247 476237
rect 245469 476236 245535 476237
rect 245469 476234 245516 476236
rect 243188 476232 244247 476234
rect 243188 476176 244186 476232
rect 244242 476176 244247 476232
rect 243188 476174 244247 476176
rect 245424 476232 245516 476234
rect 245424 476176 245474 476232
rect 245424 476174 245516 476176
rect 243188 476172 243194 476174
rect 237189 476171 237255 476172
rect 244181 476171 244247 476174
rect 245469 476172 245516 476174
rect 245580 476172 245586 476236
rect 246614 476172 246620 476236
rect 246684 476234 246690 476236
rect 246941 476234 247007 476237
rect 248321 476236 248387 476237
rect 248270 476234 248276 476236
rect 246684 476232 247007 476234
rect 246684 476176 246946 476232
rect 247002 476176 247007 476232
rect 246684 476174 247007 476176
rect 248230 476174 248276 476234
rect 248340 476232 248387 476236
rect 248382 476176 248387 476232
rect 246684 476172 246690 476174
rect 245469 476171 245535 476172
rect 246941 476171 247007 476174
rect 248270 476172 248276 476174
rect 248340 476172 248387 476176
rect 248638 476172 248644 476236
rect 248708 476234 248714 476236
rect 249701 476234 249767 476237
rect 248708 476232 249767 476234
rect 248708 476176 249706 476232
rect 249762 476176 249767 476232
rect 248708 476174 249767 476176
rect 248708 476172 248714 476174
rect 248321 476171 248387 476172
rect 249701 476171 249767 476174
rect 250846 476172 250852 476236
rect 250916 476234 250922 476236
rect 250989 476234 251055 476237
rect 250916 476232 251055 476234
rect 250916 476176 250994 476232
rect 251050 476176 251055 476232
rect 250916 476174 251055 476176
rect 250916 476172 250922 476174
rect 250989 476171 251055 476174
rect 252318 476172 252324 476236
rect 252388 476234 252394 476236
rect 252461 476234 252527 476237
rect 252388 476232 252527 476234
rect 252388 476176 252466 476232
rect 252522 476176 252527 476232
rect 252388 476174 252527 476176
rect 252388 476172 252394 476174
rect 252461 476171 252527 476174
rect 253606 476172 253612 476236
rect 253676 476234 253682 476236
rect 253841 476234 253907 476237
rect 253676 476232 253907 476234
rect 253676 476176 253846 476232
rect 253902 476176 253907 476232
rect 253676 476174 253907 476176
rect 253676 476172 253682 476174
rect 253841 476171 253907 476174
rect 254526 476172 254532 476236
rect 254596 476234 254602 476236
rect 255221 476234 255287 476237
rect 254596 476232 255287 476234
rect 254596 476176 255226 476232
rect 255282 476176 255287 476232
rect 254596 476174 255287 476176
rect 254596 476172 254602 476174
rect 255221 476171 255287 476174
rect 255814 476172 255820 476236
rect 255884 476234 255890 476236
rect 256509 476234 256575 476237
rect 255884 476232 256575 476234
rect 255884 476176 256514 476232
rect 256570 476176 256575 476232
rect 255884 476174 256575 476176
rect 255884 476172 255890 476174
rect 256509 476171 256575 476174
rect 257102 476172 257108 476236
rect 257172 476234 257178 476236
rect 257981 476234 258047 476237
rect 257172 476232 258047 476234
rect 257172 476176 257986 476232
rect 258042 476176 258047 476232
rect 257172 476174 258047 476176
rect 257172 476172 257178 476174
rect 257981 476171 258047 476174
rect 258574 476172 258580 476236
rect 258644 476234 258650 476236
rect 259269 476234 259335 476237
rect 258644 476232 259335 476234
rect 258644 476176 259274 476232
rect 259330 476176 259335 476232
rect 258644 476174 259335 476176
rect 258644 476172 258650 476174
rect 259269 476171 259335 476174
rect 260598 476172 260604 476236
rect 260668 476234 260674 476236
rect 260741 476234 260807 476237
rect 260668 476232 260807 476234
rect 260668 476176 260746 476232
rect 260802 476176 260807 476232
rect 260668 476174 260807 476176
rect 260668 476172 260674 476174
rect 260741 476171 260807 476174
rect 261702 476172 261708 476236
rect 261772 476234 261778 476236
rect 262029 476234 262095 476237
rect 261772 476232 262095 476234
rect 261772 476176 262034 476232
rect 262090 476176 262095 476232
rect 261772 476174 262095 476176
rect 261772 476172 261778 476174
rect 262029 476171 262095 476174
rect 262806 476172 262812 476236
rect 262876 476234 262882 476236
rect 263501 476234 263567 476237
rect 262876 476232 263567 476234
rect 262876 476176 263506 476232
rect 263562 476176 263567 476232
rect 262876 476174 263567 476176
rect 262876 476172 262882 476174
rect 263501 476171 263567 476174
rect 263910 476172 263916 476236
rect 263980 476234 263986 476236
rect 264881 476234 264947 476237
rect 263980 476232 264947 476234
rect 263980 476176 264886 476232
rect 264942 476176 264947 476232
rect 263980 476174 264947 476176
rect 263980 476172 263986 476174
rect 264881 476171 264947 476174
rect 265382 476172 265388 476236
rect 265452 476234 265458 476236
rect 266169 476234 266235 476237
rect 267549 476236 267615 476237
rect 267549 476234 267596 476236
rect 265452 476232 266235 476234
rect 265452 476176 266174 476232
rect 266230 476176 266235 476232
rect 265452 476174 266235 476176
rect 267504 476232 267596 476234
rect 267504 476176 267554 476232
rect 267504 476174 267596 476176
rect 265452 476172 265458 476174
rect 266169 476171 266235 476174
rect 267549 476172 267596 476174
rect 267660 476172 267666 476236
rect 268694 476172 268700 476236
rect 268764 476234 268770 476236
rect 269021 476234 269087 476237
rect 268764 476232 269087 476234
rect 268764 476176 269026 476232
rect 269082 476176 269087 476232
rect 268764 476174 269087 476176
rect 268764 476172 268770 476174
rect 267549 476171 267615 476172
rect 269021 476171 269087 476174
rect 269798 476172 269804 476236
rect 269868 476234 269874 476236
rect 270401 476234 270467 476237
rect 269868 476232 270467 476234
rect 269868 476176 270406 476232
rect 270462 476176 270467 476232
rect 269868 476174 270467 476176
rect 269868 476172 269874 476174
rect 270401 476171 270467 476174
rect 271270 476172 271276 476236
rect 271340 476234 271346 476236
rect 271689 476234 271755 476237
rect 271340 476232 271755 476234
rect 271340 476176 271694 476232
rect 271750 476176 271755 476232
rect 271340 476174 271755 476176
rect 271340 476172 271346 476174
rect 271689 476171 271755 476174
rect 272190 476172 272196 476236
rect 272260 476234 272266 476236
rect 273161 476234 273227 476237
rect 274357 476236 274423 476237
rect 275921 476236 275987 476237
rect 274357 476234 274404 476236
rect 272260 476232 273227 476234
rect 272260 476176 273166 476232
rect 273222 476176 273227 476232
rect 272260 476174 273227 476176
rect 274312 476232 274404 476234
rect 274312 476176 274362 476232
rect 274312 476174 274404 476176
rect 272260 476172 272266 476174
rect 273161 476171 273227 476174
rect 274357 476172 274404 476174
rect 274468 476172 274474 476236
rect 275870 476172 275876 476236
rect 275940 476234 275987 476236
rect 275940 476232 276032 476234
rect 275982 476176 276032 476232
rect 275940 476174 276032 476176
rect 275940 476172 275987 476174
rect 276974 476172 276980 476236
rect 277044 476234 277050 476236
rect 277209 476234 277275 476237
rect 277044 476232 277275 476234
rect 277044 476176 277214 476232
rect 277270 476176 277275 476232
rect 277044 476174 277275 476176
rect 277044 476172 277050 476174
rect 274357 476171 274423 476172
rect 275921 476171 275987 476172
rect 277209 476171 277275 476174
rect 278446 476172 278452 476236
rect 278516 476234 278522 476236
rect 278681 476234 278747 476237
rect 278516 476232 278747 476234
rect 278516 476176 278686 476232
rect 278742 476176 278747 476232
rect 278516 476174 278747 476176
rect 278516 476172 278522 476174
rect 278681 476171 278747 476174
rect 279182 476172 279188 476236
rect 279252 476234 279258 476236
rect 280061 476234 280127 476237
rect 279252 476232 280127 476234
rect 279252 476176 280066 476232
rect 280122 476176 280127 476232
rect 279252 476174 280127 476176
rect 279252 476172 279258 476174
rect 280061 476171 280127 476174
rect 281022 476172 281028 476236
rect 281092 476234 281098 476236
rect 281441 476234 281507 476237
rect 281092 476232 281507 476234
rect 281092 476176 281446 476232
rect 281502 476176 281507 476232
rect 281092 476174 281507 476176
rect 281092 476172 281098 476174
rect 281441 476171 281507 476174
rect 283598 476172 283604 476236
rect 283668 476234 283674 476236
rect 284201 476234 284267 476237
rect 283668 476232 284267 476234
rect 283668 476176 284206 476232
rect 284262 476176 284267 476232
rect 283668 476174 284267 476176
rect 283668 476172 283674 476174
rect 284201 476171 284267 476174
rect 285990 476172 285996 476236
rect 286060 476234 286066 476236
rect 286501 476234 286567 476237
rect 286060 476232 286567 476234
rect 286060 476176 286506 476232
rect 286562 476176 286567 476232
rect 286060 476174 286567 476176
rect 286060 476172 286066 476174
rect 286501 476171 286567 476174
rect 288198 476172 288204 476236
rect 288268 476234 288274 476236
rect 288341 476234 288407 476237
rect 288268 476232 288407 476234
rect 288268 476176 288346 476232
rect 288402 476176 288407 476232
rect 288268 476174 288407 476176
rect 288268 476172 288274 476174
rect 288341 476171 288407 476174
rect 290958 476172 290964 476236
rect 291028 476234 291034 476236
rect 291101 476234 291167 476237
rect 291028 476232 291167 476234
rect 291028 476176 291106 476232
rect 291162 476176 291167 476232
rect 291028 476174 291167 476176
rect 291028 476172 291034 476174
rect 291101 476171 291167 476174
rect 293534 476172 293540 476236
rect 293604 476234 293610 476236
rect 293861 476234 293927 476237
rect 293604 476232 293927 476234
rect 293604 476176 293866 476232
rect 293922 476176 293927 476232
rect 293604 476174 293927 476176
rect 293604 476172 293610 476174
rect 293861 476171 293927 476174
rect 295926 476172 295932 476236
rect 295996 476234 296002 476236
rect 296621 476234 296687 476237
rect 295996 476232 296687 476234
rect 295996 476176 296626 476232
rect 296682 476176 296687 476232
rect 295996 476174 296687 476176
rect 295996 476172 296002 476174
rect 296621 476171 296687 476174
rect 298502 476172 298508 476236
rect 298572 476234 298578 476236
rect 299381 476234 299447 476237
rect 298572 476232 299447 476234
rect 298572 476176 299386 476232
rect 299442 476176 299447 476232
rect 298572 476174 299447 476176
rect 298572 476172 298578 476174
rect 299381 476171 299447 476174
rect 300894 476172 300900 476236
rect 300964 476234 300970 476236
rect 302141 476234 302207 476237
rect 303521 476236 303587 476237
rect 300964 476232 302207 476234
rect 300964 476176 302146 476232
rect 302202 476176 302207 476232
rect 300964 476174 302207 476176
rect 300964 476172 300970 476174
rect 302141 476171 302207 476174
rect 303470 476172 303476 476236
rect 303540 476234 303587 476236
rect 303540 476232 303632 476234
rect 303582 476176 303632 476232
rect 303540 476174 303632 476176
rect 303540 476172 303587 476174
rect 306046 476172 306052 476236
rect 306116 476234 306122 476236
rect 306281 476234 306347 476237
rect 306116 476232 306347 476234
rect 306116 476176 306286 476232
rect 306342 476176 306347 476232
rect 306116 476174 306347 476176
rect 306116 476172 306122 476174
rect 303521 476171 303587 476172
rect 306281 476171 306347 476174
rect 315798 476172 315804 476236
rect 315868 476234 315874 476236
rect 315941 476234 316007 476237
rect 315868 476232 316007 476234
rect 315868 476176 315946 476232
rect 316002 476176 316007 476232
rect 315868 476174 316007 476176
rect 315868 476172 315874 476174
rect 315941 476171 316007 476174
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3233 462634 3299 462637
rect -960 462632 3299 462634
rect -960 462576 3238 462632
rect 3294 462576 3299 462632
rect -960 462574 3299 462576
rect -960 462484 480 462574
rect 3233 462571 3299 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 4061 449578 4127 449581
rect -960 449576 4127 449578
rect -960 449520 4066 449576
rect 4122 449520 4127 449576
rect -960 449518 4127 449520
rect -960 449428 480 449518
rect 4061 449515 4127 449518
rect 243721 445906 243787 445909
rect 369342 445906 369348 445908
rect 243721 445904 369348 445906
rect 243721 445848 243726 445904
rect 243782 445848 369348 445904
rect 243721 445846 369348 445848
rect 243721 445843 243787 445846
rect 369342 445844 369348 445846
rect 369412 445844 369418 445908
rect 237833 445770 237899 445773
rect 367870 445770 367876 445772
rect 237833 445768 367876 445770
rect 237833 445712 237838 445768
rect 237894 445712 367876 445768
rect 237833 445710 367876 445712
rect 237833 445707 237899 445710
rect 367870 445708 367876 445710
rect 367940 445708 367946 445772
rect 216070 444892 216076 444956
rect 216140 444954 216146 444956
rect 297449 444954 297515 444957
rect 216140 444952 297515 444954
rect 216140 444896 297454 444952
rect 297510 444896 297515 444952
rect 216140 444894 297515 444896
rect 216140 444892 216146 444894
rect 297449 444891 297515 444894
rect 214598 444756 214604 444820
rect 214668 444818 214674 444820
rect 299381 444818 299447 444821
rect 214668 444816 299447 444818
rect 214668 444760 299386 444816
rect 299442 444760 299447 444816
rect 214668 444758 299447 444760
rect 214668 444756 214674 444758
rect 299381 444755 299447 444758
rect 234613 444682 234679 444685
rect 364926 444682 364932 444684
rect 234613 444680 364932 444682
rect 234613 444624 234618 444680
rect 234674 444624 364932 444680
rect 234613 444622 364932 444624
rect 234613 444619 234679 444622
rect 364926 444620 364932 444622
rect 364996 444620 365002 444684
rect 583520 444668 584960 444908
rect 238569 444546 238635 444549
rect 368974 444546 368980 444548
rect 238569 444544 368980 444546
rect 238569 444488 238574 444544
rect 238630 444488 368980 444544
rect 238569 444486 368980 444488
rect 238569 444483 238635 444486
rect 368974 444484 368980 444486
rect 369044 444484 369050 444548
rect 236545 444410 236611 444413
rect 367686 444410 367692 444412
rect 236545 444408 367692 444410
rect 236545 444352 236550 444408
rect 236606 444352 367692 444408
rect 236545 444350 367692 444352
rect 236545 444347 236611 444350
rect 367686 444348 367692 444350
rect 367756 444348 367762 444412
rect 235257 443322 235323 443325
rect 362534 443322 362540 443324
rect 235257 443320 362540 443322
rect 235257 443264 235262 443320
rect 235318 443264 362540 443320
rect 235257 443262 362540 443264
rect 235257 443259 235323 443262
rect 362534 443260 362540 443262
rect 362604 443260 362610 443324
rect 239857 443186 239923 443189
rect 580533 443186 580599 443189
rect 239857 443184 580599 443186
rect 239857 443128 239862 443184
rect 239918 443128 580538 443184
rect 580594 443128 580599 443184
rect 239857 443126 580599 443128
rect 239857 443123 239923 443126
rect 580533 443123 580599 443126
rect 232681 443050 232747 443053
rect 580257 443050 580323 443053
rect 232681 443048 580323 443050
rect 232681 442992 232686 443048
rect 232742 442992 580262 443048
rect 580318 442992 580323 443048
rect 232681 442990 580323 442992
rect 232681 442987 232747 442990
rect 580257 442987 580323 442990
rect 246941 442234 247007 442237
rect 580349 442234 580415 442237
rect 246941 442232 580415 442234
rect 246941 442176 246946 442232
rect 247002 442176 580354 442232
rect 580410 442176 580415 442232
rect 246941 442174 580415 442176
rect 246941 442171 247007 442174
rect 580349 442171 580415 442174
rect 215886 441764 215892 441828
rect 215956 441826 215962 441828
rect 306005 441826 306071 441829
rect 215956 441824 306071 441826
rect 215956 441768 306010 441824
rect 306066 441768 306071 441824
rect 215956 441766 306071 441768
rect 215956 441764 215962 441766
rect 306005 441763 306071 441766
rect 243077 441690 243143 441693
rect 362718 441690 362724 441692
rect 243077 441688 362724 441690
rect 243077 441632 243082 441688
rect 243138 441632 362724 441688
rect 243077 441630 362724 441632
rect 243077 441627 243143 441630
rect 362718 441628 362724 441630
rect 362788 441628 362794 441692
rect 289813 441282 289879 441285
rect 293769 441282 293835 441285
rect 289813 441280 293835 441282
rect 289813 441224 289818 441280
rect 289874 441224 293774 441280
rect 293830 441224 293835 441280
rect 289813 441222 293835 441224
rect 289813 441219 289879 441222
rect 293769 441219 293835 441222
rect 290733 441146 290799 441149
rect 293677 441146 293743 441149
rect 290733 441144 293743 441146
rect 290733 441088 290738 441144
rect 290794 441088 293682 441144
rect 293738 441088 293743 441144
rect 290733 441086 293743 441088
rect 290733 441083 290799 441086
rect 293677 441083 293743 441086
rect 304993 441010 305059 441013
rect 292530 441008 305059 441010
rect 292530 440952 304998 441008
rect 305054 440952 305059 441008
rect 292530 440950 305059 440952
rect 95877 440330 95943 440333
rect 292530 440330 292590 440950
rect 304993 440947 305059 440950
rect 95877 440328 292590 440330
rect 95877 440272 95882 440328
rect 95938 440272 292590 440328
rect 95877 440270 292590 440272
rect 95877 440267 95943 440270
rect -960 436508 480 436748
rect 580073 431626 580139 431629
rect 583520 431626 584960 431716
rect 580073 431624 584960 431626
rect 580073 431568 580078 431624
rect 580134 431568 584960 431624
rect 580073 431566 584960 431568
rect 580073 431563 580139 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3325 423602 3391 423605
rect -960 423600 3391 423602
rect -960 423544 3330 423600
rect 3386 423544 3391 423600
rect -960 423542 3391 423544
rect -960 423452 480 423542
rect 3325 423539 3391 423542
rect 579981 418298 580047 418301
rect 583520 418298 584960 418388
rect 579981 418296 584960 418298
rect 579981 418240 579986 418296
rect 580042 418240 584960 418296
rect 579981 418238 584960 418240
rect 579981 418235 580047 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 2957 410546 3023 410549
rect -960 410544 3023 410546
rect -960 410488 2962 410544
rect 3018 410488 3023 410544
rect -960 410486 3023 410488
rect -960 410396 480 410486
rect 2957 410483 3023 410486
rect 579797 404970 579863 404973
rect 583520 404970 584960 405060
rect 579797 404968 584960 404970
rect 579797 404912 579802 404968
rect 579858 404912 584960 404968
rect 579797 404910 584960 404912
rect 579797 404907 579863 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3049 397490 3115 397493
rect -960 397488 3115 397490
rect -960 397432 3054 397488
rect 3110 397432 3115 397488
rect -960 397430 3115 397432
rect -960 397340 480 397430
rect 3049 397427 3115 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580073 378450 580139 378453
rect 583520 378450 584960 378540
rect 580073 378448 584960 378450
rect 580073 378392 580078 378448
rect 580134 378392 584960 378448
rect 580073 378390 584960 378392
rect 580073 378387 580139 378390
rect 583520 378300 584960 378390
rect 159909 374098 159975 374101
rect 232078 374098 232084 374100
rect 159909 374096 232084 374098
rect 159909 374040 159914 374096
rect 159970 374040 232084 374096
rect 159909 374038 232084 374040
rect 159909 374035 159975 374038
rect 232078 374036 232084 374038
rect 232148 374036 232154 374100
rect 155861 373282 155927 373285
rect 231894 373282 231900 373284
rect 155861 373280 231900 373282
rect 155861 373224 155866 373280
rect 155922 373224 231900 373280
rect 155861 373222 231900 373224
rect 155861 373219 155927 373222
rect 231894 373220 231900 373222
rect 231964 373220 231970 373284
rect 124673 371650 124739 371653
rect 135069 371650 135135 371653
rect 124673 371648 135135 371650
rect 124673 371592 124678 371648
rect 124734 371592 135074 371648
rect 135130 371592 135135 371648
rect 124673 371590 135135 371592
rect 124673 371587 124739 371590
rect 135069 371587 135135 371590
rect 137921 371650 137987 371653
rect 144177 371650 144243 371653
rect 137921 371648 144243 371650
rect 137921 371592 137926 371648
rect 137982 371592 144182 371648
rect 144238 371592 144243 371648
rect 137921 371590 144243 371592
rect 137921 371587 137987 371590
rect 144177 371587 144243 371590
rect -960 371378 480 371468
rect 3141 371378 3207 371381
rect -960 371376 3207 371378
rect -960 371320 3146 371376
rect 3202 371320 3207 371376
rect -960 371318 3207 371320
rect -960 371228 480 371318
rect 3141 371315 3207 371318
rect 99833 370698 99899 370701
rect 99833 370696 100218 370698
rect 99833 370640 99838 370696
rect 99894 370640 100218 370696
rect 99833 370638 100218 370640
rect 99833 370635 99899 370638
rect 100158 370124 100218 370638
rect 172329 369474 172395 369477
rect 169924 369472 172395 369474
rect 169924 369416 172334 369472
rect 172390 369416 172395 369472
rect 169924 369414 172395 369416
rect 172329 369411 172395 369414
rect 97901 367434 97967 367437
rect 97901 367432 100188 367434
rect 97901 367376 97906 367432
rect 97962 367376 100188 367432
rect 97901 367374 100188 367376
rect 97901 367371 97967 367374
rect 172421 366754 172487 366757
rect 169924 366752 172487 366754
rect 169924 366696 172426 366752
rect 172482 366696 172487 366752
rect 169924 366694 172487 366696
rect 172421 366691 172487 366694
rect 580073 365122 580139 365125
rect 583520 365122 584960 365212
rect 580073 365120 584960 365122
rect 580073 365064 580078 365120
rect 580134 365064 584960 365120
rect 580073 365062 584960 365064
rect 580073 365059 580139 365062
rect 583520 364972 584960 365062
rect 97717 364714 97783 364717
rect 97717 364712 100188 364714
rect 97717 364656 97722 364712
rect 97778 364656 100188 364712
rect 97717 364654 100188 364656
rect 97717 364651 97783 364654
rect 172329 364034 172395 364037
rect 169924 364032 172395 364034
rect 169924 363976 172334 364032
rect 172390 363976 172395 364032
rect 169924 363974 172395 363976
rect 172329 363971 172395 363974
rect 97625 361994 97691 361997
rect 97625 361992 100188 361994
rect 97625 361936 97630 361992
rect 97686 361936 100188 361992
rect 97625 361934 100188 361936
rect 97625 361931 97691 361934
rect 171869 361314 171935 361317
rect 169924 361312 171935 361314
rect 169924 361256 171874 361312
rect 171930 361256 171935 361312
rect 169924 361254 171935 361256
rect 171869 361251 171935 361254
rect 99281 359274 99347 359277
rect 99281 359272 100188 359274
rect 99281 359216 99286 359272
rect 99342 359216 100188 359272
rect 99281 359214 100188 359216
rect 99281 359211 99347 359214
rect 171685 358594 171751 358597
rect 169924 358592 171751 358594
rect -960 358458 480 358548
rect 169924 358536 171690 358592
rect 171746 358536 171751 358592
rect 169924 358534 171751 358536
rect 171685 358531 171751 358534
rect 3785 358458 3851 358461
rect -960 358456 3851 358458
rect -960 358400 3790 358456
rect 3846 358400 3851 358456
rect -960 358398 3851 358400
rect -960 358308 480 358398
rect 3785 358395 3851 358398
rect 97901 356554 97967 356557
rect 97901 356552 100188 356554
rect 97901 356496 97906 356552
rect 97962 356496 100188 356552
rect 97901 356494 100188 356496
rect 97901 356491 97967 356494
rect 171961 355874 172027 355877
rect 169924 355872 172027 355874
rect 169924 355816 171966 355872
rect 172022 355816 172027 355872
rect 169924 355814 172027 355816
rect 171961 355811 172027 355814
rect 99189 353834 99255 353837
rect 99189 353832 100188 353834
rect 99189 353776 99194 353832
rect 99250 353776 100188 353832
rect 99189 353774 100188 353776
rect 99189 353771 99255 353774
rect 172421 353154 172487 353157
rect 169924 353152 172487 353154
rect 169924 353096 172426 353152
rect 172482 353096 172487 353152
rect 169924 353094 172487 353096
rect 172421 353091 172487 353094
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect 97809 351114 97875 351117
rect 97809 351112 100188 351114
rect 97809 351056 97814 351112
rect 97870 351056 100188 351112
rect 97809 351054 100188 351056
rect 97809 351051 97875 351054
rect 171133 350434 171199 350437
rect 169924 350432 171199 350434
rect 169924 350376 171138 350432
rect 171194 350376 171199 350432
rect 169924 350374 171199 350376
rect 171133 350371 171199 350374
rect 97809 348394 97875 348397
rect 97809 348392 100188 348394
rect 97809 348336 97814 348392
rect 97870 348336 100188 348392
rect 97809 348334 100188 348336
rect 97809 348331 97875 348334
rect 172421 347714 172487 347717
rect 169924 347712 172487 347714
rect 169924 347656 172426 347712
rect 172482 347656 172487 347712
rect 169924 347654 172487 347656
rect 172421 347651 172487 347654
rect 97717 345674 97783 345677
rect 97717 345672 100188 345674
rect 97717 345616 97722 345672
rect 97778 345616 100188 345672
rect 97717 345614 100188 345616
rect 97717 345611 97783 345614
rect -960 345402 480 345492
rect 3693 345402 3759 345405
rect -960 345400 3759 345402
rect -960 345344 3698 345400
rect 3754 345344 3759 345400
rect -960 345342 3759 345344
rect -960 345252 480 345342
rect 3693 345339 3759 345342
rect 172053 344994 172119 344997
rect 169924 344992 172119 344994
rect 169924 344936 172058 344992
rect 172114 344936 172119 344992
rect 169924 344934 172119 344936
rect 172053 344931 172119 344934
rect 99373 342954 99439 342957
rect 99373 342952 100188 342954
rect 99373 342896 99378 342952
rect 99434 342896 100188 342952
rect 99373 342894 100188 342896
rect 99373 342891 99439 342894
rect 172145 342274 172211 342277
rect 169924 342272 172211 342274
rect 169924 342216 172150 342272
rect 172206 342216 172211 342272
rect 169924 342214 172211 342216
rect 172145 342211 172211 342214
rect 97625 340234 97691 340237
rect 97625 340232 100188 340234
rect 97625 340176 97630 340232
rect 97686 340176 100188 340232
rect 97625 340174 100188 340176
rect 97625 340171 97691 340174
rect 172237 339554 172303 339557
rect 169924 339552 172303 339554
rect 169924 339496 172242 339552
rect 172298 339496 172303 339552
rect 169924 339494 172303 339496
rect 172237 339491 172303 339494
rect 583520 338452 584960 338692
rect 99097 337514 99163 337517
rect 99097 337512 100188 337514
rect 99097 337456 99102 337512
rect 99158 337456 100188 337512
rect 99097 337454 100188 337456
rect 99097 337451 99163 337454
rect 172421 336834 172487 336837
rect 169924 336832 172487 336834
rect 169924 336776 172426 336832
rect 172482 336776 172487 336832
rect 169924 336774 172487 336776
rect 172421 336771 172487 336774
rect 97533 334794 97599 334797
rect 97533 334792 100188 334794
rect 97533 334736 97538 334792
rect 97594 334736 100188 334792
rect 97533 334734 100188 334736
rect 97533 334731 97599 334734
rect 172421 334114 172487 334117
rect 169924 334112 172487 334114
rect 169924 334056 172426 334112
rect 172482 334056 172487 334112
rect 169924 334054 172487 334056
rect 172421 334051 172487 334054
rect -960 332196 480 332436
rect 97441 332074 97507 332077
rect 97441 332072 100188 332074
rect 97441 332016 97446 332072
rect 97502 332016 100188 332072
rect 97441 332014 100188 332016
rect 97441 332011 97507 332014
rect 172421 331394 172487 331397
rect 169924 331392 172487 331394
rect 169924 331336 172426 331392
rect 172482 331336 172487 331392
rect 169924 331334 172487 331336
rect 172421 331331 172487 331334
rect 99005 329354 99071 329357
rect 99005 329352 100188 329354
rect 99005 329296 99010 329352
rect 99066 329296 100188 329352
rect 99005 329294 100188 329296
rect 99005 329291 99071 329294
rect 172329 328674 172395 328677
rect 169924 328672 172395 328674
rect 169924 328616 172334 328672
rect 172390 328616 172395 328672
rect 169924 328614 172395 328616
rect 172329 328611 172395 328614
rect 97349 326634 97415 326637
rect 97349 326632 100188 326634
rect 97349 326576 97354 326632
rect 97410 326576 100188 326632
rect 97349 326574 100188 326576
rect 97349 326571 97415 326574
rect 172421 325954 172487 325957
rect 169924 325952 172487 325954
rect 169924 325896 172426 325952
rect 172482 325896 172487 325952
rect 169924 325894 172487 325896
rect 172421 325891 172487 325894
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 98913 323914 98979 323917
rect 98913 323912 100188 323914
rect 98913 323856 98918 323912
rect 98974 323856 100188 323912
rect 98913 323854 100188 323856
rect 98913 323851 98979 323854
rect 171317 323234 171383 323237
rect 169924 323232 171383 323234
rect 169924 323176 171322 323232
rect 171378 323176 171383 323232
rect 169924 323174 171383 323176
rect 171317 323171 171383 323174
rect 99465 321194 99531 321197
rect 99465 321192 100188 321194
rect 99465 321136 99470 321192
rect 99526 321136 100188 321192
rect 99465 321134 100188 321136
rect 99465 321131 99531 321134
rect 171501 320514 171567 320517
rect 169924 320512 171567 320514
rect 169924 320456 171506 320512
rect 171562 320456 171567 320512
rect 169924 320454 171567 320456
rect 171501 320451 171567 320454
rect -960 319290 480 319380
rect 2957 319290 3023 319293
rect -960 319288 3023 319290
rect -960 319232 2962 319288
rect 3018 319232 3023 319288
rect -960 319230 3023 319232
rect -960 319140 480 319230
rect 2957 319227 3023 319230
rect 98821 318474 98887 318477
rect 98821 318472 100188 318474
rect 98821 318416 98826 318472
rect 98882 318416 100188 318472
rect 98821 318414 100188 318416
rect 98821 318411 98887 318414
rect 171501 317794 171567 317797
rect 169924 317792 171567 317794
rect 169924 317736 171506 317792
rect 171562 317736 171567 317792
rect 169924 317734 171567 317736
rect 171501 317731 171567 317734
rect 98729 315754 98795 315757
rect 98729 315752 100188 315754
rect 98729 315696 98734 315752
rect 98790 315696 100188 315752
rect 98729 315694 100188 315696
rect 98729 315691 98795 315694
rect 172421 315074 172487 315077
rect 169924 315072 172487 315074
rect 169924 315016 172426 315072
rect 172482 315016 172487 315072
rect 169924 315014 172487 315016
rect 172421 315011 172487 315014
rect 99557 313034 99623 313037
rect 99557 313032 100188 313034
rect 99557 312976 99562 313032
rect 99618 312976 100188 313032
rect 99557 312974 100188 312976
rect 99557 312971 99623 312974
rect 172421 312354 172487 312357
rect 169924 312352 172487 312354
rect 169924 312296 172426 312352
rect 172482 312296 172487 312352
rect 169924 312294 172487 312296
rect 172421 312291 172487 312294
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect 232078 311204 232084 311268
rect 232148 311266 232154 311268
rect 232221 311266 232287 311269
rect 232148 311264 232287 311266
rect 232148 311208 232226 311264
rect 232282 311208 232287 311264
rect 232148 311206 232287 311208
rect 232148 311204 232154 311206
rect 232221 311203 232287 311206
rect 172053 310858 172119 310861
rect 172053 310856 233986 310858
rect 172053 310800 172058 310856
rect 172114 310800 233986 310856
rect 172053 310798 233986 310800
rect 172053 310795 172119 310798
rect 225781 310586 225847 310589
rect 233693 310586 233759 310589
rect 225781 310584 233759 310586
rect 225781 310528 225786 310584
rect 225842 310528 233698 310584
rect 233754 310528 233759 310584
rect 225781 310526 233759 310528
rect 233926 310586 233986 310798
rect 234061 310586 234127 310589
rect 233926 310584 234127 310586
rect 233926 310528 234066 310584
rect 234122 310528 234127 310584
rect 233926 310526 234127 310528
rect 225781 310523 225847 310526
rect 233693 310523 233759 310526
rect 234061 310523 234127 310526
rect 232078 310388 232084 310452
rect 232148 310450 232154 310452
rect 232405 310450 232471 310453
rect 232148 310448 232471 310450
rect 232148 310392 232410 310448
rect 232466 310392 232471 310448
rect 232148 310390 232471 310392
rect 232148 310388 232154 310390
rect 232405 310387 232471 310390
rect 98637 310314 98703 310317
rect 98637 310312 100188 310314
rect 98637 310256 98642 310312
rect 98698 310256 100188 310312
rect 98637 310254 100188 310256
rect 98637 310251 98703 310254
rect 231894 310252 231900 310316
rect 231964 310314 231970 310316
rect 232865 310314 232931 310317
rect 231964 310312 232931 310314
rect 231964 310256 232870 310312
rect 232926 310256 232931 310312
rect 231964 310254 232931 310256
rect 231964 310252 231970 310254
rect 232865 310251 232931 310254
rect 241237 310042 241303 310045
rect 224910 310040 241303 310042
rect 224910 309984 241242 310040
rect 241298 309984 241303 310040
rect 224910 309982 241303 309984
rect 172237 309634 172303 309637
rect 169924 309632 172303 309634
rect 169924 309576 172242 309632
rect 172298 309576 172303 309632
rect 169924 309574 172303 309576
rect 172237 309571 172303 309574
rect 170949 309498 171015 309501
rect 224910 309498 224970 309982
rect 241237 309979 241303 309982
rect 231209 309906 231275 309909
rect 240317 309906 240383 309909
rect 231209 309904 240383 309906
rect 231209 309848 231214 309904
rect 231270 309848 240322 309904
rect 240378 309848 240383 309904
rect 231209 309846 240383 309848
rect 231209 309843 231275 309846
rect 240317 309843 240383 309846
rect 232446 309708 232452 309772
rect 232516 309770 232522 309772
rect 247309 309770 247375 309773
rect 232516 309768 247375 309770
rect 232516 309712 247314 309768
rect 247370 309712 247375 309768
rect 232516 309710 247375 309712
rect 232516 309708 232522 309710
rect 247309 309707 247375 309710
rect 228541 309634 228607 309637
rect 248137 309634 248203 309637
rect 228541 309632 248203 309634
rect 228541 309576 228546 309632
rect 228602 309576 248142 309632
rect 248198 309576 248203 309632
rect 228541 309574 248203 309576
rect 228541 309571 228607 309574
rect 248137 309571 248203 309574
rect 170949 309496 224970 309498
rect 170949 309440 170954 309496
rect 171010 309440 224970 309496
rect 170949 309438 224970 309440
rect 170949 309435 171015 309438
rect 170581 309362 170647 309365
rect 244641 309362 244707 309365
rect 170581 309360 244707 309362
rect 170581 309304 170586 309360
rect 170642 309304 244646 309360
rect 244702 309304 244707 309360
rect 170581 309302 244707 309304
rect 170581 309299 170647 309302
rect 244641 309299 244707 309302
rect 170765 309226 170831 309229
rect 251725 309226 251791 309229
rect 170765 309224 251791 309226
rect 170765 309168 170770 309224
rect 170826 309168 251730 309224
rect 251786 309168 251791 309224
rect 170765 309166 251791 309168
rect 170765 309163 170831 309166
rect 251725 309163 251791 309166
rect 231301 309090 231367 309093
rect 235717 309090 235783 309093
rect 231301 309088 235783 309090
rect 231301 309032 231306 309088
rect 231362 309032 235722 309088
rect 235778 309032 235783 309088
rect 231301 309030 235783 309032
rect 231301 309027 231367 309030
rect 235717 309027 235783 309030
rect 346945 309090 347011 309093
rect 366449 309090 366515 309093
rect 346945 309088 366515 309090
rect 346945 309032 346950 309088
rect 347006 309032 366454 309088
rect 366510 309032 366515 309088
rect 346945 309030 366515 309032
rect 346945 309027 347011 309030
rect 366449 309027 366515 309030
rect 173433 308954 173499 308957
rect 234521 308954 234587 308957
rect 173433 308952 234587 308954
rect 173433 308896 173438 308952
rect 173494 308896 234526 308952
rect 234582 308896 234587 308952
rect 173433 308894 234587 308896
rect 173433 308891 173499 308894
rect 234521 308891 234587 308894
rect 347497 308954 347563 308957
rect 366265 308954 366331 308957
rect 347497 308952 366331 308954
rect 347497 308896 347502 308952
rect 347558 308896 366270 308952
rect 366326 308896 366331 308952
rect 347497 308894 366331 308896
rect 347497 308891 347563 308894
rect 366265 308891 366331 308894
rect 231485 308818 231551 308821
rect 248321 308818 248387 308821
rect 231485 308816 248387 308818
rect 231485 308760 231490 308816
rect 231546 308760 248326 308816
rect 248382 308760 248387 308816
rect 231485 308758 248387 308760
rect 231485 308755 231551 308758
rect 248321 308755 248387 308758
rect 348417 308818 348483 308821
rect 368565 308818 368631 308821
rect 348417 308816 368631 308818
rect 348417 308760 348422 308816
rect 348478 308760 368570 308816
rect 368626 308760 368631 308816
rect 348417 308758 368631 308760
rect 348417 308755 348483 308758
rect 368565 308755 368631 308758
rect 228633 308682 228699 308685
rect 252645 308682 252711 308685
rect 228633 308680 252711 308682
rect 228633 308624 228638 308680
rect 228694 308624 252650 308680
rect 252706 308624 252711 308680
rect 228633 308622 252711 308624
rect 228633 308619 228699 308622
rect 252645 308619 252711 308622
rect 349245 308682 349311 308685
rect 370037 308682 370103 308685
rect 349245 308680 370103 308682
rect 349245 308624 349250 308680
rect 349306 308624 370042 308680
rect 370098 308624 370103 308680
rect 349245 308622 370103 308624
rect 349245 308619 349311 308622
rect 370037 308619 370103 308622
rect 169334 308484 169340 308548
rect 169404 308546 169410 308548
rect 250989 308546 251055 308549
rect 169404 308544 251055 308546
rect 169404 308488 250994 308544
rect 251050 308488 251055 308544
rect 169404 308486 251055 308488
rect 169404 308484 169410 308486
rect 250989 308483 251055 308486
rect 311065 308546 311131 308549
rect 371325 308546 371391 308549
rect 311065 308544 371391 308546
rect 311065 308488 311070 308544
rect 311126 308488 371330 308544
rect 371386 308488 371391 308544
rect 311065 308486 371391 308488
rect 311065 308483 311131 308486
rect 371325 308483 371391 308486
rect 214833 308410 214899 308413
rect 298277 308410 298343 308413
rect 214833 308408 298343 308410
rect 214833 308352 214838 308408
rect 214894 308352 298282 308408
rect 298338 308352 298343 308408
rect 214833 308350 298343 308352
rect 214833 308347 214899 308350
rect 298277 308347 298343 308350
rect 329925 308410 329991 308413
rect 462957 308410 463023 308413
rect 329925 308408 463023 308410
rect 329925 308352 329930 308408
rect 329986 308352 462962 308408
rect 463018 308352 463023 308408
rect 329925 308350 463023 308352
rect 329925 308347 329991 308350
rect 462957 308347 463023 308350
rect 173249 308274 173315 308277
rect 250345 308274 250411 308277
rect 173249 308272 250411 308274
rect 173249 308216 173254 308272
rect 173310 308216 250350 308272
rect 250406 308216 250411 308272
rect 173249 308214 250411 308216
rect 173249 308211 173315 308214
rect 250345 308211 250411 308214
rect 346761 308274 346827 308277
rect 362125 308274 362191 308277
rect 346761 308272 362191 308274
rect 346761 308216 346766 308272
rect 346822 308216 362130 308272
rect 362186 308216 362191 308272
rect 346761 308214 362191 308216
rect 346761 308211 346827 308214
rect 362125 308211 362191 308214
rect 99833 307594 99899 307597
rect 99833 307592 100188 307594
rect 99833 307536 99838 307592
rect 99894 307536 100188 307592
rect 99833 307534 100188 307536
rect 99833 307531 99899 307534
rect 171409 306914 171475 306917
rect 169924 306912 171475 306914
rect 169924 306856 171414 306912
rect 171470 306856 171475 306912
rect 169924 306854 171475 306856
rect 171409 306851 171475 306854
rect 350993 306370 351059 306373
rect 370129 306370 370195 306373
rect 350993 306368 370195 306370
rect -960 306234 480 306324
rect 350993 306312 350998 306368
rect 351054 306312 370134 306368
rect 370190 306312 370195 306368
rect 350993 306310 370195 306312
rect 350993 306307 351059 306310
rect 370129 306307 370195 306310
rect 3325 306234 3391 306237
rect -960 306232 3391 306234
rect -960 306176 3330 306232
rect 3386 306176 3391 306232
rect -960 306174 3391 306176
rect -960 306084 480 306174
rect 3325 306171 3391 306174
rect 218830 306172 218836 306236
rect 218900 306234 218906 306236
rect 288341 306234 288407 306237
rect 218900 306232 288407 306234
rect 218900 306176 288346 306232
rect 288402 306176 288407 306232
rect 218900 306174 288407 306176
rect 218900 306172 218906 306174
rect 288341 306171 288407 306174
rect 349981 306234 350047 306237
rect 369025 306234 369091 306237
rect 349981 306232 369091 306234
rect 349981 306176 349986 306232
rect 350042 306176 369030 306232
rect 369086 306176 369091 306232
rect 349981 306174 369091 306176
rect 349981 306171 350047 306174
rect 369025 306171 369091 306174
rect 219014 306036 219020 306100
rect 219084 306098 219090 306100
rect 288893 306098 288959 306101
rect 219084 306096 288959 306098
rect 219084 306040 288898 306096
rect 288954 306040 288959 306096
rect 219084 306038 288959 306040
rect 219084 306036 219090 306038
rect 288893 306035 288959 306038
rect 319345 306098 319411 306101
rect 377397 306098 377463 306101
rect 319345 306096 377463 306098
rect 319345 306040 319350 306096
rect 319406 306040 377402 306096
rect 377458 306040 377463 306096
rect 319345 306038 377463 306040
rect 319345 306035 319411 306038
rect 377397 306035 377463 306038
rect 219198 305900 219204 305964
rect 219268 305962 219274 305964
rect 288709 305962 288775 305965
rect 219268 305960 288775 305962
rect 219268 305904 288714 305960
rect 288770 305904 288775 305960
rect 219268 305902 288775 305904
rect 219268 305900 219274 305902
rect 288709 305899 288775 305902
rect 298093 305962 298159 305965
rect 358261 305962 358327 305965
rect 298093 305960 358327 305962
rect 298093 305904 298098 305960
rect 298154 305904 358266 305960
rect 358322 305904 358327 305960
rect 298093 305902 358327 305904
rect 298093 305899 298159 305902
rect 358261 305899 358327 305902
rect 217358 305764 217364 305828
rect 217428 305826 217434 305828
rect 290089 305826 290155 305829
rect 217428 305824 290155 305826
rect 217428 305768 290094 305824
rect 290150 305768 290155 305824
rect 217428 305766 290155 305768
rect 217428 305764 217434 305766
rect 290089 305763 290155 305766
rect 315389 305826 315455 305829
rect 385033 305826 385099 305829
rect 315389 305824 385099 305826
rect 315389 305768 315394 305824
rect 315450 305768 385038 305824
rect 385094 305768 385099 305824
rect 315389 305766 385099 305768
rect 315389 305763 315455 305766
rect 385033 305763 385099 305766
rect 217174 305628 217180 305692
rect 217244 305690 217250 305692
rect 291745 305690 291811 305693
rect 217244 305688 291811 305690
rect 217244 305632 291750 305688
rect 291806 305632 291811 305688
rect 217244 305630 291811 305632
rect 217244 305628 217250 305630
rect 291745 305627 291811 305630
rect 345105 305690 345171 305693
rect 570597 305690 570663 305693
rect 345105 305688 570663 305690
rect 345105 305632 345110 305688
rect 345166 305632 570602 305688
rect 570658 305632 570663 305688
rect 345105 305630 570663 305632
rect 345105 305627 345171 305630
rect 570597 305627 570663 305630
rect 97901 304874 97967 304877
rect 97901 304872 100188 304874
rect 97901 304816 97906 304872
rect 97962 304816 100188 304872
rect 97901 304814 100188 304816
rect 97901 304811 97967 304814
rect 172329 304194 172395 304197
rect 169924 304192 172395 304194
rect 169924 304136 172334 304192
rect 172390 304136 172395 304192
rect 169924 304134 172395 304136
rect 172329 304131 172395 304134
rect 312353 303514 312419 303517
rect 369894 303514 369900 303516
rect 312353 303512 369900 303514
rect 312353 303456 312358 303512
rect 312414 303456 369900 303512
rect 312353 303454 369900 303456
rect 312353 303451 312419 303454
rect 369894 303452 369900 303454
rect 369964 303452 369970 303516
rect 216254 303316 216260 303380
rect 216324 303378 216330 303380
rect 287605 303378 287671 303381
rect 216324 303376 287671 303378
rect 216324 303320 287610 303376
rect 287666 303320 287671 303376
rect 216324 303318 287671 303320
rect 216324 303316 216330 303318
rect 287605 303315 287671 303318
rect 298829 303378 298895 303381
rect 367093 303378 367159 303381
rect 298829 303376 367159 303378
rect 298829 303320 298834 303376
rect 298890 303320 367098 303376
rect 367154 303320 367159 303376
rect 298829 303318 367159 303320
rect 298829 303315 298895 303318
rect 367093 303315 367159 303318
rect 215150 303180 215156 303244
rect 215220 303242 215226 303244
rect 287513 303242 287579 303245
rect 215220 303240 287579 303242
rect 215220 303184 287518 303240
rect 287574 303184 287579 303240
rect 215220 303182 287579 303184
rect 215220 303180 215226 303182
rect 287513 303179 287579 303182
rect 318241 303242 318307 303245
rect 396717 303242 396783 303245
rect 318241 303240 396783 303242
rect 318241 303184 318246 303240
rect 318302 303184 396722 303240
rect 396778 303184 396783 303240
rect 318241 303182 396783 303184
rect 318241 303179 318307 303182
rect 396717 303179 396783 303182
rect 170489 303106 170555 303109
rect 260097 303106 260163 303109
rect 170489 303104 260163 303106
rect 170489 303048 170494 303104
rect 170550 303048 260102 303104
rect 260158 303048 260163 303104
rect 170489 303046 260163 303048
rect 170489 303043 170555 303046
rect 260097 303043 260163 303046
rect 331673 303106 331739 303109
rect 489177 303106 489243 303109
rect 331673 303104 489243 303106
rect 331673 303048 331678 303104
rect 331734 303048 489182 303104
rect 489238 303048 489243 303104
rect 331673 303046 489243 303048
rect 331673 303043 331739 303046
rect 489177 303043 489243 303046
rect 184933 302970 184999 302973
rect 282637 302970 282703 302973
rect 184933 302968 282703 302970
rect 184933 302912 184938 302968
rect 184994 302912 282642 302968
rect 282698 302912 282703 302968
rect 184933 302910 282703 302912
rect 184933 302907 184999 302910
rect 282637 302907 282703 302910
rect 337285 302970 337351 302973
rect 520917 302970 520983 302973
rect 337285 302968 520983 302970
rect 337285 302912 337290 302968
rect 337346 302912 520922 302968
rect 520978 302912 520983 302968
rect 337285 302910 520983 302912
rect 337285 302907 337351 302910
rect 520917 302907 520983 302910
rect 182173 302834 182239 302837
rect 282085 302834 282151 302837
rect 182173 302832 282151 302834
rect 182173 302776 182178 302832
rect 182234 302776 282090 302832
rect 282146 302776 282151 302832
rect 182173 302774 282151 302776
rect 182173 302771 182239 302774
rect 282085 302771 282151 302774
rect 341701 302834 341767 302837
rect 545757 302834 545823 302837
rect 341701 302832 545823 302834
rect 341701 302776 341706 302832
rect 341762 302776 545762 302832
rect 545818 302776 545823 302832
rect 341701 302774 545823 302776
rect 341701 302771 341767 302774
rect 545757 302771 545823 302774
rect 99741 301610 99807 301613
rect 100158 301610 100218 302124
rect 99741 301608 100218 301610
rect 99741 301552 99746 301608
rect 99802 301552 100218 301608
rect 99741 301550 100218 301552
rect 99741 301547 99807 301550
rect 169518 301548 169524 301612
rect 169588 301610 169594 301612
rect 236269 301610 236335 301613
rect 169588 301608 236335 301610
rect 169588 301552 236274 301608
rect 236330 301552 236335 301608
rect 169588 301550 236335 301552
rect 169588 301548 169594 301550
rect 236269 301547 236335 301550
rect 172421 301474 172487 301477
rect 169924 301472 172487 301474
rect 169924 301416 172426 301472
rect 172482 301416 172487 301472
rect 169924 301414 172487 301416
rect 172421 301411 172487 301414
rect 169150 301140 169156 301204
rect 169220 301202 169226 301204
rect 248597 301202 248663 301205
rect 169220 301200 248663 301202
rect 169220 301144 248602 301200
rect 248658 301144 248663 301200
rect 169220 301142 248663 301144
rect 169220 301140 169226 301142
rect 248597 301139 248663 301142
rect 99281 300794 99347 300797
rect 245653 300794 245719 300797
rect 99281 300792 245719 300794
rect 99281 300736 99286 300792
rect 99342 300736 245658 300792
rect 245714 300736 245719 300792
rect 99281 300734 245719 300736
rect 99281 300731 99347 300734
rect 245653 300731 245719 300734
rect 211981 300522 212047 300525
rect 289997 300522 290063 300525
rect 211981 300520 290063 300522
rect 211981 300464 211986 300520
rect 212042 300464 290002 300520
rect 290058 300464 290063 300520
rect 211981 300462 290063 300464
rect 211981 300459 212047 300462
rect 289997 300459 290063 300462
rect 164233 300386 164299 300389
rect 279325 300386 279391 300389
rect 164233 300384 279391 300386
rect 164233 300328 164238 300384
rect 164294 300328 279330 300384
rect 279386 300328 279391 300384
rect 164233 300326 279391 300328
rect 164233 300323 164299 300326
rect 279325 300323 279391 300326
rect 160093 300250 160159 300253
rect 278589 300250 278655 300253
rect 160093 300248 278655 300250
rect 160093 300192 160098 300248
rect 160154 300192 278594 300248
rect 278650 300192 278655 300248
rect 160093 300190 278655 300192
rect 160093 300187 160159 300190
rect 278589 300187 278655 300190
rect 20713 300114 20779 300117
rect 255773 300114 255839 300117
rect 20713 300112 255839 300114
rect 20713 300056 20718 300112
rect 20774 300056 255778 300112
rect 255834 300056 255839 300112
rect 20713 300054 255839 300056
rect 20713 300051 20779 300054
rect 255773 300051 255839 300054
rect 299749 300114 299815 300117
rect 368422 300114 368428 300116
rect 299749 300112 368428 300114
rect 299749 300056 299754 300112
rect 299810 300056 368428 300112
rect 299749 300054 368428 300056
rect 299749 300051 299815 300054
rect 368422 300052 368428 300054
rect 368492 300052 368498 300116
rect 97441 299434 97507 299437
rect 237557 299434 237623 299437
rect 97441 299432 237623 299434
rect 97441 299376 97446 299432
rect 97502 299376 237562 299432
rect 237618 299376 237623 299432
rect 97441 299374 237623 299376
rect 97441 299371 97507 299374
rect 237557 299371 237623 299374
rect 97533 299298 97599 299301
rect 234337 299298 234403 299301
rect 97533 299296 234403 299298
rect 97533 299240 97538 299296
rect 97594 299240 234342 299296
rect 234398 299240 234403 299296
rect 97533 299238 234403 299240
rect 97533 299235 97599 299238
rect 234337 299235 234403 299238
rect 97257 299162 97323 299165
rect 169334 299162 169340 299164
rect 97257 299160 169340 299162
rect 97257 299104 97262 299160
rect 97318 299104 169340 299160
rect 97257 299102 169340 299104
rect 97257 299099 97323 299102
rect 169334 299100 169340 299102
rect 169404 299100 169410 299164
rect 580901 298754 580967 298757
rect 583520 298754 584960 298844
rect 580901 298752 584960 298754
rect 580901 298696 580906 298752
rect 580962 298696 584960 298752
rect 580901 298694 584960 298696
rect 580901 298691 580967 298694
rect 583520 298604 584960 298694
rect 101949 298074 102015 298077
rect 169150 298074 169156 298076
rect 101949 298072 169156 298074
rect 101949 298016 101954 298072
rect 102010 298016 169156 298072
rect 101949 298014 169156 298016
rect 101949 298011 102015 298014
rect 169150 298012 169156 298014
rect 169220 298012 169226 298076
rect 145741 297938 145807 297941
rect 169518 297938 169524 297940
rect 145741 297936 169524 297938
rect 145741 297880 145746 297936
rect 145802 297880 169524 297936
rect 145741 297878 169524 297880
rect 145741 297875 145807 297878
rect 169518 297876 169524 297878
rect 169588 297876 169594 297940
rect 216990 297740 216996 297804
rect 217060 297802 217066 297804
rect 293309 297802 293375 297805
rect 217060 297800 293375 297802
rect 217060 297744 293314 297800
rect 293370 297744 293375 297800
rect 217060 297742 293375 297744
rect 217060 297740 217066 297742
rect 293309 297739 293375 297742
rect 213361 297666 213427 297669
rect 290181 297666 290247 297669
rect 213361 297664 290247 297666
rect 213361 297608 213366 297664
rect 213422 297608 290186 297664
rect 290242 297608 290247 297664
rect 213361 297606 290247 297608
rect 213361 297603 213427 297606
rect 290181 297603 290247 297606
rect 213545 297530 213611 297533
rect 291561 297530 291627 297533
rect 213545 297528 291627 297530
rect 213545 297472 213550 297528
rect 213606 297472 291566 297528
rect 291622 297472 291627 297528
rect 213545 297470 291627 297472
rect 213545 297467 213611 297470
rect 291561 297467 291627 297470
rect 212073 297394 212139 297397
rect 290273 297394 290339 297397
rect 212073 297392 290339 297394
rect 212073 297336 212078 297392
rect 212134 297336 290278 297392
rect 290334 297336 290339 297392
rect 212073 297334 290339 297336
rect 212073 297331 212139 297334
rect 290273 297331 290339 297334
rect -960 293178 480 293268
rect 3601 293178 3667 293181
rect -960 293176 3667 293178
rect -960 293120 3606 293176
rect 3662 293120 3667 293176
rect -960 293118 3667 293120
rect -960 293028 480 293118
rect 3601 293115 3667 293118
rect 312077 286378 312143 286381
rect 367134 286378 367140 286380
rect 312077 286376 367140 286378
rect 312077 286320 312082 286376
rect 312138 286320 367140 286376
rect 312077 286318 367140 286320
rect 312077 286315 312143 286318
rect 367134 286316 367140 286318
rect 367204 286316 367210 286380
rect 583520 285276 584960 285516
rect 214414 284820 214420 284884
rect 214484 284882 214490 284884
rect 285949 284882 286015 284885
rect 214484 284880 286015 284882
rect 214484 284824 285954 284880
rect 286010 284824 286015 284880
rect 214484 284822 286015 284824
rect 214484 284820 214490 284822
rect 285949 284819 286015 284822
rect -960 279972 480 280212
rect 580809 272234 580875 272237
rect 583520 272234 584960 272324
rect 580809 272232 584960 272234
rect 580809 272176 580814 272232
rect 580870 272176 584960 272232
rect 580809 272174 584960 272176
rect 580809 272171 580875 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 2957 267202 3023 267205
rect -960 267200 3023 267202
rect -960 267144 2962 267200
rect 3018 267144 3023 267200
rect -960 267142 3023 267144
rect -960 267052 480 267142
rect 2957 267139 3023 267142
rect 579797 258906 579863 258909
rect 583520 258906 584960 258996
rect 579797 258904 584960 258906
rect 579797 258848 579802 258904
rect 579858 258848 584960 258904
rect 579797 258846 584960 258848
rect 579797 258843 579863 258846
rect 311065 258770 311131 258773
rect 364374 258770 364380 258772
rect 311065 258768 364380 258770
rect 311065 258712 311070 258768
rect 311126 258712 364380 258768
rect 311065 258710 364380 258712
rect 311065 258707 311131 258710
rect 364374 258708 364380 258710
rect 364444 258708 364450 258772
rect 583520 258756 584960 258846
rect 216438 255852 216444 255916
rect 216508 255914 216514 255916
rect 287145 255914 287211 255917
rect 216508 255912 287211 255914
rect 216508 255856 287150 255912
rect 287206 255856 287211 255912
rect 216508 255854 287211 255856
rect 216508 255852 216514 255854
rect 287145 255851 287211 255854
rect 310973 254690 311039 254693
rect 365662 254690 365668 254692
rect 310973 254688 365668 254690
rect 310973 254632 310978 254688
rect 311034 254632 365668 254688
rect 310973 254630 365668 254632
rect 310973 254627 311039 254630
rect 365662 254628 365668 254630
rect 365732 254628 365738 254692
rect 313273 254554 313339 254557
rect 369158 254554 369164 254556
rect 313273 254552 369164 254554
rect 313273 254496 313278 254552
rect 313334 254496 369164 254552
rect 313273 254494 369164 254496
rect 313273 254491 313339 254494
rect 369158 254492 369164 254494
rect 369228 254492 369234 254556
rect -960 254146 480 254236
rect 3325 254146 3391 254149
rect -960 254144 3391 254146
rect -960 254088 3330 254144
rect 3386 254088 3391 254144
rect -960 254086 3391 254088
rect -960 253996 480 254086
rect 3325 254083 3391 254086
rect 310789 253194 310855 253197
rect 365846 253194 365852 253196
rect 310789 253192 365852 253194
rect 310789 253136 310794 253192
rect 310850 253136 365852 253192
rect 310789 253134 365852 253136
rect 310789 253131 310855 253134
rect 365846 253132 365852 253134
rect 365916 253132 365922 253196
rect 310881 251970 310947 251973
rect 358854 251970 358860 251972
rect 310881 251968 358860 251970
rect 310881 251912 310886 251968
rect 310942 251912 358860 251968
rect 310881 251910 358860 251912
rect 310881 251907 310947 251910
rect 358854 251908 358860 251910
rect 358924 251908 358930 251972
rect 310697 251834 310763 251837
rect 362902 251834 362908 251836
rect 310697 251832 362908 251834
rect 310697 251776 310702 251832
rect 310758 251776 362908 251832
rect 310697 251774 362908 251776
rect 310697 251771 310763 251774
rect 362902 251772 362908 251774
rect 362972 251772 362978 251836
rect 303981 250882 304047 250885
rect 358118 250882 358124 250884
rect 303981 250880 358124 250882
rect 303981 250824 303986 250880
rect 304042 250824 358124 250880
rect 303981 250822 358124 250824
rect 303981 250819 304047 250822
rect 358118 250820 358124 250822
rect 358188 250820 358194 250884
rect 308397 250746 308463 250749
rect 363086 250746 363092 250748
rect 308397 250744 363092 250746
rect 308397 250688 308402 250744
rect 308458 250688 363092 250744
rect 308397 250686 363092 250688
rect 308397 250683 308463 250686
rect 363086 250684 363092 250686
rect 363156 250684 363162 250748
rect 308213 250610 308279 250613
rect 363270 250610 363276 250612
rect 308213 250608 363276 250610
rect 308213 250552 308218 250608
rect 308274 250552 363276 250608
rect 308213 250550 363276 250552
rect 308213 250547 308279 250550
rect 363270 250548 363276 250550
rect 363340 250548 363346 250612
rect 217542 250412 217548 250476
rect 217612 250474 217618 250476
rect 287053 250474 287119 250477
rect 217612 250472 287119 250474
rect 217612 250416 287058 250472
rect 287114 250416 287119 250472
rect 217612 250414 287119 250416
rect 217612 250412 217618 250414
rect 287053 250411 287119 250414
rect 303797 250474 303863 250477
rect 367318 250474 367324 250476
rect 303797 250472 367324 250474
rect 303797 250416 303802 250472
rect 303858 250416 367324 250472
rect 303797 250414 367324 250416
rect 303797 250411 303863 250414
rect 367318 250412 367324 250414
rect 367388 250412 367394 250476
rect 310605 248298 310671 248301
rect 360142 248298 360148 248300
rect 310605 248296 360148 248298
rect 310605 248240 310610 248296
rect 310666 248240 360148 248296
rect 310605 248238 360148 248240
rect 310605 248235 310671 248238
rect 360142 248236 360148 248238
rect 360212 248236 360218 248300
rect 305269 248162 305335 248165
rect 359038 248162 359044 248164
rect 305269 248160 359044 248162
rect 305269 248104 305274 248160
rect 305330 248104 359044 248160
rect 305269 248102 359044 248104
rect 305269 248099 305335 248102
rect 359038 248100 359044 248102
rect 359108 248100 359114 248164
rect 309225 248026 309291 248029
rect 363454 248026 363460 248028
rect 309225 248024 363460 248026
rect 309225 247968 309230 248024
rect 309286 247968 363460 248024
rect 309225 247966 363460 247968
rect 309225 247963 309291 247966
rect 363454 247964 363460 247966
rect 363524 247964 363530 248028
rect 309409 247890 309475 247893
rect 364742 247890 364748 247892
rect 309409 247888 364748 247890
rect 309409 247832 309414 247888
rect 309470 247832 364748 247888
rect 309409 247830 364748 247832
rect 309409 247827 309475 247830
rect 364742 247828 364748 247830
rect 364812 247828 364818 247892
rect 308121 247754 308187 247757
rect 364558 247754 364564 247756
rect 308121 247752 364564 247754
rect 308121 247696 308126 247752
rect 308182 247696 364564 247752
rect 308121 247694 364564 247696
rect 308121 247691 308187 247694
rect 364558 247692 364564 247694
rect 364628 247692 364634 247756
rect 336733 247618 336799 247621
rect 524413 247618 524479 247621
rect 336733 247616 524479 247618
rect 336733 247560 336738 247616
rect 336794 247560 524418 247616
rect 524474 247560 524479 247616
rect 336733 247558 524479 247560
rect 336733 247555 336799 247558
rect 524413 247555 524479 247558
rect 309133 245578 309199 245581
rect 358670 245578 358676 245580
rect 309133 245576 358676 245578
rect 309133 245520 309138 245576
rect 309194 245520 358676 245576
rect 309133 245518 358676 245520
rect 309133 245515 309199 245518
rect 358670 245516 358676 245518
rect 358740 245516 358746 245580
rect 578877 245578 578943 245581
rect 583520 245578 584960 245668
rect 578877 245576 584960 245578
rect 578877 245520 578882 245576
rect 578938 245520 584960 245576
rect 578877 245518 584960 245520
rect 578877 245515 578943 245518
rect 309317 245442 309383 245445
rect 360694 245442 360700 245444
rect 309317 245440 360700 245442
rect 309317 245384 309322 245440
rect 309378 245384 360700 245440
rect 309317 245382 360700 245384
rect 309317 245379 309383 245382
rect 360694 245380 360700 245382
rect 360764 245380 360770 245444
rect 583520 245428 584960 245518
rect 306465 245306 306531 245309
rect 359406 245306 359412 245308
rect 306465 245304 359412 245306
rect 306465 245248 306470 245304
rect 306526 245248 359412 245304
rect 306465 245246 359412 245248
rect 306465 245243 306531 245246
rect 359406 245244 359412 245246
rect 359476 245244 359482 245308
rect 305361 245170 305427 245173
rect 359222 245170 359228 245172
rect 305361 245168 359228 245170
rect 305361 245112 305366 245168
rect 305422 245112 359228 245168
rect 305361 245110 359228 245112
rect 305361 245107 305427 245110
rect 359222 245108 359228 245110
rect 359292 245108 359298 245172
rect 305177 245034 305243 245037
rect 360510 245034 360516 245036
rect 305177 245032 360516 245034
rect 305177 244976 305182 245032
rect 305238 244976 360516 245032
rect 305177 244974 360516 244976
rect 305177 244971 305243 244974
rect 360510 244972 360516 244974
rect 360580 244972 360586 245036
rect 304993 244898 305059 244901
rect 360326 244898 360332 244900
rect 304993 244896 360332 244898
rect 304993 244840 304998 244896
rect 305054 244840 360332 244896
rect 304993 244838 360332 244840
rect 304993 244835 305059 244838
rect 360326 244836 360332 244838
rect 360396 244836 360402 244900
rect 310513 244762 310579 244765
rect 358302 244762 358308 244764
rect 310513 244760 358308 244762
rect 310513 244704 310518 244760
rect 310574 244704 358308 244760
rect 310513 244702 358308 244704
rect 310513 244699 310579 244702
rect 358302 244700 358308 244702
rect 358372 244700 358378 244764
rect 363413 243810 363479 243813
rect 354630 243808 363479 243810
rect 354630 243752 363418 243808
rect 363474 243752 363479 243808
rect 354630 243750 363479 243752
rect 303613 243674 303679 243677
rect 354630 243674 354690 243750
rect 363413 243747 363479 243750
rect 359641 243674 359707 243677
rect 303613 243672 354690 243674
rect 303613 243616 303618 243672
rect 303674 243616 354690 243672
rect 303613 243614 354690 243616
rect 356654 243672 359707 243674
rect 356654 243616 359646 243672
rect 359702 243616 359707 243672
rect 356654 243614 359707 243616
rect 303613 243611 303679 243614
rect 298645 243538 298711 243541
rect 356654 243538 356714 243614
rect 359641 243611 359707 243614
rect 298645 243536 356714 243538
rect 298645 243480 298650 243536
rect 298706 243480 356714 243536
rect 298645 243478 356714 243480
rect 356881 243538 356947 243541
rect 358486 243538 358492 243540
rect 356881 243536 358492 243538
rect 356881 243480 356886 243536
rect 356942 243480 358492 243536
rect 356881 243478 358492 243480
rect 298645 243475 298711 243478
rect 356881 243475 356947 243478
rect 358486 243476 358492 243478
rect 358556 243476 358562 243540
rect -960 241090 480 241180
rect 3509 241090 3575 241093
rect -960 241088 3575 241090
rect -960 241032 3514 241088
rect 3570 241032 3575 241088
rect -960 241030 3575 241032
rect -960 240940 480 241030
rect 3509 241027 3575 241030
rect 583520 232386 584960 232476
rect 583342 232326 584960 232386
rect 583342 232250 583402 232326
rect 583520 232250 584960 232326
rect 583342 232236 584960 232250
rect 583342 232190 583586 232236
rect 362718 231916 362724 231980
rect 362788 231978 362794 231980
rect 583526 231978 583586 232190
rect 362788 231918 583586 231978
rect 362788 231916 362794 231918
rect -960 227884 480 228124
rect 583520 219058 584960 219148
rect 583342 218998 584960 219058
rect 583342 218922 583402 218998
rect 583520 218922 584960 218998
rect 583342 218908 584960 218922
rect 583342 218862 583586 218908
rect 369342 218044 369348 218108
rect 369412 218106 369418 218108
rect 583526 218106 583586 218862
rect 369412 218046 583586 218106
rect 369412 218044 369418 218046
rect -960 214978 480 215068
rect -960 214918 674 214978
rect -960 214842 480 214918
rect 614 214842 674 214918
rect -960 214828 674 214842
rect 246 214782 674 214828
rect 246 214298 306 214782
rect 246 214238 6930 214298
rect 6870 214026 6930 214238
rect 216070 214026 216076 214028
rect 6870 213966 216076 214026
rect 216070 213964 216076 213966
rect 216140 213964 216146 214028
rect 579613 205730 579679 205733
rect 583520 205730 584960 205820
rect 579613 205728 584960 205730
rect 579613 205672 579618 205728
rect 579674 205672 584960 205728
rect 579613 205670 584960 205672
rect 579613 205667 579679 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3049 201922 3115 201925
rect -960 201920 3115 201922
rect -960 201864 3054 201920
rect 3110 201864 3115 201920
rect -960 201862 3115 201864
rect -960 201772 480 201862
rect 3049 201859 3115 201862
rect 217685 196890 217751 196893
rect 219390 196890 220064 196924
rect 217685 196888 220064 196890
rect 217685 196832 217690 196888
rect 217746 196864 220064 196888
rect 217746 196832 219450 196864
rect 217685 196830 219450 196832
rect 217685 196827 217751 196830
rect 217317 195938 217383 195941
rect 219390 195938 220064 195972
rect 217317 195936 220064 195938
rect 217317 195880 217322 195936
rect 217378 195912 220064 195936
rect 217378 195880 219450 195912
rect 217317 195878 219450 195880
rect 217317 195875 217383 195878
rect 217777 193762 217843 193765
rect 219390 193762 220064 193796
rect 217777 193760 220064 193762
rect 217777 193704 217782 193760
rect 217838 193736 220064 193760
rect 217838 193704 219450 193736
rect 217777 193702 219450 193704
rect 217777 193699 217843 193702
rect 218605 193220 218671 193221
rect 218605 193218 218652 193220
rect 218560 193216 218652 193218
rect 218560 193160 218610 193216
rect 218560 193158 218652 193160
rect 218605 193156 218652 193158
rect 218716 193156 218722 193220
rect 218605 193155 218671 193156
rect 217133 192810 217199 192813
rect 219390 192810 220064 192844
rect 217133 192808 220064 192810
rect 217133 192752 217138 192808
rect 217194 192784 220064 192808
rect 217194 192752 219450 192784
rect 217133 192750 219450 192752
rect 217133 192747 217199 192750
rect 580717 192538 580783 192541
rect 583520 192538 584960 192628
rect 580717 192536 584960 192538
rect 580717 192480 580722 192536
rect 580778 192480 584960 192536
rect 580717 192478 584960 192480
rect 580717 192475 580783 192478
rect 583520 192388 584960 192478
rect 218421 191042 218487 191045
rect 219390 191042 220064 191076
rect 218421 191040 220064 191042
rect 218421 190984 218426 191040
rect 218482 191016 220064 191040
rect 218482 190984 219450 191016
rect 218421 190982 219450 190984
rect 218421 190979 218487 190982
rect 218513 189954 218579 189957
rect 219390 189954 220064 189988
rect 218513 189952 220064 189954
rect 218513 189896 218518 189952
rect 218574 189928 220064 189952
rect 218574 189896 219450 189928
rect 218513 189894 219450 189896
rect 218513 189891 218579 189894
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 216673 188186 216739 188189
rect 219390 188186 220064 188220
rect 216673 188184 220064 188186
rect 216673 188128 216678 188184
rect 216734 188160 220064 188184
rect 216734 188128 219450 188160
rect 216673 188126 219450 188128
rect 216673 188123 216739 188126
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 217593 169962 217659 169965
rect 219390 169962 220064 169996
rect 217593 169960 220064 169962
rect 217593 169904 217598 169960
rect 217654 169936 220064 169960
rect 217654 169904 219450 169936
rect 217593 169902 219450 169904
rect 217593 169899 217659 169902
rect 217409 168330 217475 168333
rect 219390 168330 220064 168364
rect 217409 168328 220064 168330
rect 217409 168272 217414 168328
rect 217470 168304 220064 168328
rect 217470 168272 219450 168304
rect 217409 168270 219450 168272
rect 217409 168267 217475 168270
rect 217225 168058 217291 168061
rect 219390 168058 220064 168092
rect 217225 168056 220064 168058
rect 217225 168000 217230 168056
rect 217286 168032 220064 168056
rect 217286 168000 219450 168032
rect 217225 167998 219450 168000
rect 217225 167995 217291 167998
rect 579613 165882 579679 165885
rect 583520 165882 584960 165972
rect 579613 165880 584960 165882
rect 579613 165824 579618 165880
rect 579674 165824 584960 165880
rect 579613 165822 584960 165824
rect 579613 165819 579679 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 214598 162890 214604 162892
rect -960 162830 214604 162890
rect -960 162740 480 162830
rect 214598 162828 214604 162830
rect 214668 162828 214674 162892
rect 258533 159900 258599 159901
rect 275829 159900 275895 159901
rect 277025 159900 277091 159901
rect 278129 159900 278195 159901
rect 279233 159900 279299 159901
rect 258488 159898 258494 159900
rect 258442 159838 258494 159898
rect 258558 159896 258599 159900
rect 275760 159898 275766 159900
rect 258594 159840 258599 159896
rect 258488 159836 258494 159838
rect 258558 159836 258599 159840
rect 275738 159838 275766 159898
rect 275760 159836 275766 159838
rect 275830 159896 275895 159900
rect 276984 159898 276990 159900
rect 275830 159840 275834 159896
rect 275890 159840 275895 159896
rect 275830 159836 275895 159840
rect 276934 159838 276990 159898
rect 277054 159896 277091 159900
rect 278072 159898 278078 159900
rect 277086 159840 277091 159896
rect 276984 159836 276990 159838
rect 277054 159836 277091 159840
rect 278038 159838 278078 159898
rect 278142 159896 278195 159900
rect 279160 159898 279166 159900
rect 278190 159840 278195 159896
rect 278072 159836 278078 159838
rect 278142 159836 278195 159840
rect 279142 159838 279166 159898
rect 279160 159836 279166 159838
rect 279230 159896 279299 159900
rect 279230 159840 279238 159896
rect 279294 159840 279299 159896
rect 279230 159836 279299 159840
rect 258533 159835 258599 159836
rect 275829 159835 275895 159836
rect 277025 159835 277091 159836
rect 278129 159835 278195 159836
rect 279233 159835 279299 159836
rect 300945 159764 301011 159765
rect 300920 159762 300926 159764
rect 300854 159702 300926 159762
rect 300990 159760 301011 159764
rect 301006 159704 301011 159760
rect 300920 159700 300926 159702
rect 300990 159700 301011 159704
rect 300945 159699 301011 159700
rect 255957 159628 256023 159629
rect 271045 159628 271111 159629
rect 274449 159628 274515 159629
rect 255904 159626 255910 159628
rect 255866 159566 255910 159626
rect 255974 159624 256023 159628
rect 271000 159626 271006 159628
rect 256018 159568 256023 159624
rect 255904 159564 255910 159566
rect 255974 159564 256023 159568
rect 270954 159566 271006 159626
rect 271070 159624 271111 159628
rect 274400 159626 274406 159628
rect 271106 159568 271111 159624
rect 271000 159564 271006 159566
rect 271070 159564 271111 159568
rect 274358 159566 274406 159626
rect 274470 159624 274515 159628
rect 274510 159568 274515 159624
rect 274400 159564 274406 159566
rect 274470 159564 274515 159568
rect 255957 159563 256023 159564
rect 271045 159563 271111 159564
rect 274449 159563 274515 159564
rect 357341 159490 357407 159493
rect 362125 159490 362191 159493
rect 357341 159488 362191 159490
rect 357341 159432 357346 159488
rect 357402 159432 362130 159488
rect 362186 159432 362191 159488
rect 357341 159430 362191 159432
rect 357341 159427 357407 159430
rect 362125 159427 362191 159430
rect 296713 159354 296779 159357
rect 369301 159354 369367 159357
rect 296713 159352 369367 159354
rect 296713 159296 296718 159352
rect 296774 159296 369306 159352
rect 369362 159296 369367 159352
rect 296713 159294 369367 159296
rect 296713 159291 296779 159294
rect 369301 159291 369367 159294
rect 254526 159156 254532 159220
rect 254596 159218 254602 159220
rect 365069 159218 365135 159221
rect 254596 159216 365135 159218
rect 254596 159160 365074 159216
rect 365130 159160 365135 159216
rect 254596 159158 365135 159160
rect 254596 159156 254602 159158
rect 365069 159155 365135 159158
rect 250846 159020 250852 159084
rect 250916 159082 250922 159084
rect 372061 159082 372127 159085
rect 250916 159080 372127 159082
rect 250916 159024 372066 159080
rect 372122 159024 372127 159080
rect 250916 159022 372127 159024
rect 250916 159020 250922 159022
rect 372061 159019 372127 159022
rect 243118 158884 243124 158948
rect 243188 158946 243194 158948
rect 366449 158946 366515 158949
rect 243188 158944 366515 158946
rect 243188 158888 366454 158944
rect 366510 158888 366515 158944
rect 243188 158886 366515 158888
rect 243188 158884 243194 158886
rect 366449 158883 366515 158886
rect 236126 158748 236132 158812
rect 236196 158810 236202 158812
rect 357341 158810 357407 158813
rect 236196 158808 357407 158810
rect 236196 158752 357346 158808
rect 357402 158752 357407 158808
rect 236196 158750 357407 158752
rect 236196 158748 236202 158750
rect 357341 158747 357407 158750
rect 358077 158810 358143 158813
rect 358670 158810 358676 158812
rect 358077 158808 358676 158810
rect 358077 158752 358082 158808
rect 358138 158752 358676 158808
rect 358077 158750 358676 158752
rect 358077 158747 358143 158750
rect 358670 158748 358676 158750
rect 358740 158748 358746 158812
rect 360694 158748 360700 158812
rect 360764 158810 360770 158812
rect 361113 158810 361179 158813
rect 360764 158808 361179 158810
rect 360764 158752 361118 158808
rect 361174 158752 361179 158808
rect 360764 158750 361179 158752
rect 360764 158748 360770 158750
rect 361113 158747 361179 158750
rect 364742 158748 364748 158812
rect 364812 158810 364818 158812
rect 365253 158810 365319 158813
rect 364812 158808 365319 158810
rect 364812 158752 365258 158808
rect 365314 158752 365319 158808
rect 364812 158750 365319 158752
rect 364812 158748 364818 158750
rect 365253 158747 365319 158750
rect 218830 158612 218836 158676
rect 218900 158674 218906 158676
rect 220813 158674 220879 158677
rect 218900 158672 220879 158674
rect 218900 158616 220818 158672
rect 220874 158616 220879 158672
rect 218900 158614 220879 158616
rect 218900 158612 218906 158614
rect 220813 158611 220879 158614
rect 238109 158676 238175 158677
rect 239581 158676 239647 158677
rect 238109 158672 238156 158676
rect 238220 158674 238226 158676
rect 238109 158616 238114 158672
rect 238109 158612 238156 158616
rect 238220 158614 238266 158674
rect 239581 158672 239628 158676
rect 239692 158674 239698 158676
rect 239581 158616 239586 158672
rect 238220 158612 238226 158614
rect 239581 158612 239628 158616
rect 239692 158614 239738 158674
rect 239692 158612 239698 158614
rect 240542 158612 240548 158676
rect 240612 158674 240618 158676
rect 240685 158674 240751 158677
rect 248321 158676 248387 158677
rect 250161 158676 250227 158677
rect 248270 158674 248276 158676
rect 240612 158672 240751 158674
rect 240612 158616 240690 158672
rect 240746 158616 240751 158672
rect 240612 158614 240751 158616
rect 248230 158614 248276 158674
rect 248340 158672 248387 158676
rect 250110 158674 250116 158676
rect 248382 158616 248387 158672
rect 240612 158612 240618 158614
rect 238109 158611 238175 158612
rect 239581 158611 239647 158612
rect 240685 158611 240751 158614
rect 248270 158612 248276 158614
rect 248340 158612 248387 158616
rect 250070 158614 250116 158674
rect 250180 158672 250227 158676
rect 250222 158616 250227 158672
rect 250110 158612 250116 158614
rect 250180 158612 250227 158616
rect 255998 158612 256004 158676
rect 256068 158674 256074 158676
rect 256601 158674 256667 158677
rect 257153 158676 257219 158677
rect 257102 158674 257108 158676
rect 256068 158672 256667 158674
rect 256068 158616 256606 158672
rect 256662 158616 256667 158672
rect 256068 158614 256667 158616
rect 257062 158614 257108 158674
rect 257172 158672 257219 158676
rect 257214 158616 257219 158672
rect 256068 158612 256074 158614
rect 248321 158611 248387 158612
rect 250161 158611 250227 158612
rect 256601 158611 256667 158614
rect 257102 158612 257108 158614
rect 257172 158612 257219 158616
rect 258206 158612 258212 158676
rect 258276 158674 258282 158676
rect 258625 158674 258691 158677
rect 259545 158676 259611 158677
rect 259494 158674 259500 158676
rect 258276 158672 258691 158674
rect 258276 158616 258630 158672
rect 258686 158616 258691 158672
rect 258276 158614 258691 158616
rect 259454 158614 259500 158674
rect 259564 158672 259611 158676
rect 259606 158616 259611 158672
rect 258276 158612 258282 158614
rect 257153 158611 257219 158612
rect 258625 158611 258691 158614
rect 259494 158612 259500 158614
rect 259564 158612 259611 158616
rect 261150 158612 261156 158676
rect 261220 158674 261226 158676
rect 261753 158674 261819 158677
rect 262857 158676 262923 158677
rect 265985 158676 266051 158677
rect 267641 158676 267707 158677
rect 268745 158676 268811 158677
rect 262806 158674 262812 158676
rect 261220 158672 261819 158674
rect 261220 158616 261758 158672
rect 261814 158616 261819 158672
rect 261220 158614 261819 158616
rect 262766 158614 262812 158674
rect 262876 158672 262923 158676
rect 265934 158674 265940 158676
rect 262918 158616 262923 158672
rect 261220 158612 261226 158614
rect 259545 158611 259611 158612
rect 261753 158611 261819 158614
rect 262806 158612 262812 158614
rect 262876 158612 262923 158616
rect 265894 158614 265940 158674
rect 266004 158672 266051 158676
rect 267590 158674 267596 158676
rect 266046 158616 266051 158672
rect 265934 158612 265940 158614
rect 266004 158612 266051 158616
rect 267550 158614 267596 158674
rect 267660 158672 267707 158676
rect 268694 158674 268700 158676
rect 267702 158616 267707 158672
rect 267590 158612 267596 158614
rect 267660 158612 267707 158616
rect 268654 158614 268700 158674
rect 268764 158672 268811 158676
rect 268806 158616 268811 158672
rect 268694 158612 268700 158614
rect 268764 158612 268811 158616
rect 269798 158612 269804 158676
rect 269868 158674 269874 158676
rect 270217 158674 270283 158677
rect 271137 158676 271203 158677
rect 272241 158676 272307 158677
rect 271086 158674 271092 158676
rect 269868 158672 270283 158674
rect 269868 158616 270222 158672
rect 270278 158616 270283 158672
rect 269868 158614 270283 158616
rect 271046 158614 271092 158674
rect 271156 158672 271203 158676
rect 272190 158674 272196 158676
rect 271198 158616 271203 158672
rect 269868 158612 269874 158614
rect 262857 158611 262923 158612
rect 265985 158611 266051 158612
rect 267641 158611 267707 158612
rect 268745 158611 268811 158612
rect 270217 158611 270283 158614
rect 271086 158612 271092 158614
rect 271156 158612 271203 158616
rect 272150 158614 272196 158674
rect 272260 158672 272307 158676
rect 272302 158616 272307 158672
rect 272190 158612 272196 158614
rect 272260 158612 272307 158616
rect 298502 158612 298508 158676
rect 298572 158674 298578 158676
rect 298921 158674 298987 158677
rect 303521 158676 303587 158677
rect 306097 158676 306163 158677
rect 308673 158676 308739 158677
rect 313457 158676 313523 158677
rect 315849 158676 315915 158677
rect 318609 158676 318675 158677
rect 303470 158674 303476 158676
rect 298572 158672 298987 158674
rect 298572 158616 298926 158672
rect 298982 158616 298987 158672
rect 298572 158614 298987 158616
rect 303430 158614 303476 158674
rect 303540 158672 303587 158676
rect 306046 158674 306052 158676
rect 303582 158616 303587 158672
rect 298572 158612 298578 158614
rect 271137 158611 271203 158612
rect 272241 158611 272307 158612
rect 298921 158611 298987 158614
rect 303470 158612 303476 158614
rect 303540 158612 303587 158616
rect 306006 158614 306052 158674
rect 306116 158672 306163 158676
rect 308622 158674 308628 158676
rect 306158 158616 306163 158672
rect 306046 158612 306052 158614
rect 306116 158612 306163 158616
rect 308582 158614 308628 158674
rect 308692 158672 308739 158676
rect 313406 158674 313412 158676
rect 308734 158616 308739 158672
rect 308622 158612 308628 158614
rect 308692 158612 308739 158616
rect 313366 158614 313412 158674
rect 313476 158672 313523 158676
rect 315798 158674 315804 158676
rect 313518 158616 313523 158672
rect 313406 158612 313412 158614
rect 313476 158612 313523 158616
rect 315758 158614 315804 158674
rect 315868 158672 315915 158676
rect 318558 158674 318564 158676
rect 315910 158616 315915 158672
rect 315798 158612 315804 158614
rect 315868 158612 315915 158616
rect 318518 158614 318564 158674
rect 318628 158672 318675 158676
rect 318670 158616 318675 158672
rect 318558 158612 318564 158614
rect 318628 158612 318675 158616
rect 320950 158612 320956 158676
rect 321020 158674 321026 158676
rect 321185 158674 321251 158677
rect 323393 158676 323459 158677
rect 325969 158676 326035 158677
rect 323342 158674 323348 158676
rect 321020 158672 321251 158674
rect 321020 158616 321190 158672
rect 321246 158616 321251 158672
rect 321020 158614 321251 158616
rect 323302 158614 323348 158674
rect 323412 158672 323459 158676
rect 325918 158674 325924 158676
rect 323454 158616 323459 158672
rect 321020 158612 321026 158614
rect 303521 158611 303587 158612
rect 306097 158611 306163 158612
rect 308673 158611 308739 158612
rect 313457 158611 313523 158612
rect 315849 158611 315915 158612
rect 318609 158611 318675 158612
rect 321185 158611 321251 158614
rect 323342 158612 323348 158614
rect 323412 158612 323459 158616
rect 325878 158614 325924 158674
rect 325988 158672 326035 158676
rect 326030 158616 326035 158672
rect 325918 158612 325924 158614
rect 325988 158612 326035 158616
rect 323393 158611 323459 158612
rect 325969 158611 326035 158612
rect 219014 158476 219020 158540
rect 219084 158538 219090 158540
rect 224953 158538 225019 158541
rect 252369 158540 252435 158541
rect 260649 158540 260715 158541
rect 276105 158540 276171 158541
rect 252318 158538 252324 158540
rect 219084 158536 225019 158538
rect 219084 158480 224958 158536
rect 225014 158480 225019 158536
rect 219084 158478 225019 158480
rect 252278 158478 252324 158538
rect 252388 158536 252435 158540
rect 260598 158538 260604 158540
rect 252430 158480 252435 158536
rect 219084 158476 219090 158478
rect 224953 158475 225019 158478
rect 252318 158476 252324 158478
rect 252388 158476 252435 158480
rect 260558 158478 260604 158538
rect 260668 158536 260715 158540
rect 276054 158538 276060 158540
rect 260710 158480 260715 158536
rect 260598 158476 260604 158478
rect 260668 158476 260715 158480
rect 276014 158478 276060 158538
rect 276124 158536 276171 158540
rect 276166 158480 276171 158536
rect 276054 158476 276060 158478
rect 276124 158476 276171 158480
rect 281022 158476 281028 158540
rect 281092 158538 281098 158540
rect 281349 158538 281415 158541
rect 281092 158536 281415 158538
rect 281092 158480 281354 158536
rect 281410 158480 281415 158536
rect 281092 158478 281415 158480
rect 281092 158476 281098 158478
rect 252369 158475 252435 158476
rect 260649 158475 260715 158476
rect 276105 158475 276171 158476
rect 281349 158475 281415 158478
rect 285990 158476 285996 158540
rect 286060 158538 286066 158540
rect 286225 158538 286291 158541
rect 286060 158536 286291 158538
rect 286060 158480 286230 158536
rect 286286 158480 286291 158536
rect 286060 158478 286291 158480
rect 286060 158476 286066 158478
rect 286225 158475 286291 158478
rect 353937 158538 354003 158541
rect 358261 158538 358327 158541
rect 353937 158536 358327 158538
rect 353937 158480 353942 158536
rect 353998 158480 358266 158536
rect 358322 158480 358327 158536
rect 353937 158478 358327 158480
rect 353937 158475 354003 158478
rect 358261 158475 358327 158478
rect 219198 158340 219204 158404
rect 219268 158402 219274 158404
rect 227713 158402 227779 158405
rect 273345 158404 273411 158405
rect 291009 158404 291075 158405
rect 273294 158402 273300 158404
rect 219268 158400 227779 158402
rect 219268 158344 227718 158400
rect 227774 158344 227779 158400
rect 219268 158342 227779 158344
rect 273254 158342 273300 158402
rect 273364 158400 273411 158404
rect 290958 158402 290964 158404
rect 273406 158344 273411 158400
rect 219268 158340 219274 158342
rect 227713 158339 227779 158342
rect 273294 158340 273300 158342
rect 273364 158340 273411 158344
rect 290918 158342 290964 158402
rect 291028 158400 291075 158404
rect 291070 158344 291075 158400
rect 290958 158340 290964 158342
rect 291028 158340 291075 158344
rect 295926 158340 295932 158404
rect 295996 158402 296002 158404
rect 296253 158402 296319 158405
rect 295996 158400 296319 158402
rect 295996 158344 296258 158400
rect 296314 158344 296319 158400
rect 295996 158342 296319 158344
rect 295996 158340 296002 158342
rect 273345 158339 273411 158340
rect 291009 158339 291075 158340
rect 296253 158339 296319 158342
rect 354121 158402 354187 158405
rect 363781 158402 363847 158405
rect 354121 158400 363847 158402
rect 354121 158344 354126 158400
rect 354182 158344 363786 158400
rect 363842 158344 363847 158400
rect 354121 158342 363847 158344
rect 354121 158339 354187 158342
rect 363781 158339 363847 158342
rect 216254 158204 216260 158268
rect 216324 158266 216330 158268
rect 219433 158266 219499 158269
rect 216324 158264 219499 158266
rect 216324 158208 219438 158264
rect 219494 158208 219499 158264
rect 216324 158206 219499 158208
rect 216324 158204 216330 158206
rect 219433 158203 219499 158206
rect 244222 158204 244228 158268
rect 244292 158266 244298 158268
rect 245377 158266 245443 158269
rect 244292 158264 245443 158266
rect 244292 158208 245382 158264
rect 245438 158208 245443 158264
rect 244292 158206 245443 158208
rect 244292 158204 244298 158206
rect 245377 158203 245443 158206
rect 311014 158204 311020 158268
rect 311084 158266 311090 158268
rect 311249 158266 311315 158269
rect 311084 158264 311315 158266
rect 311084 158208 311254 158264
rect 311310 158208 311315 158264
rect 311084 158206 311315 158208
rect 311084 158204 311090 158206
rect 311249 158203 311315 158206
rect 348417 158266 348483 158269
rect 362401 158266 362467 158269
rect 348417 158264 362467 158266
rect 348417 158208 348422 158264
rect 348478 158208 362406 158264
rect 362462 158208 362467 158264
rect 348417 158206 362467 158208
rect 348417 158203 348483 158206
rect 362401 158203 362467 158206
rect 217358 158068 217364 158132
rect 217428 158130 217434 158132
rect 231853 158130 231919 158133
rect 217428 158128 231919 158130
rect 217428 158072 231858 158128
rect 231914 158072 231919 158128
rect 217428 158070 231919 158072
rect 217428 158068 217434 158070
rect 231853 158067 231919 158070
rect 246614 158068 246620 158132
rect 246684 158130 246690 158132
rect 246849 158130 246915 158133
rect 246684 158128 246915 158130
rect 246684 158072 246854 158128
rect 246910 158072 246915 158128
rect 246684 158070 246915 158072
rect 246684 158068 246690 158070
rect 246849 158067 246915 158070
rect 351177 158130 351243 158133
rect 365161 158130 365227 158133
rect 351177 158128 365227 158130
rect 351177 158072 351182 158128
rect 351238 158072 365166 158128
rect 365222 158072 365227 158128
rect 351177 158070 365227 158072
rect 351177 158067 351243 158070
rect 365161 158067 365227 158070
rect 217174 157932 217180 157996
rect 217244 157994 217250 157996
rect 238753 157994 238819 157997
rect 248689 157996 248755 157997
rect 248638 157994 248644 157996
rect 217244 157992 238819 157994
rect 217244 157936 238758 157992
rect 238814 157936 238819 157992
rect 217244 157934 238819 157936
rect 248598 157934 248644 157994
rect 248708 157992 248755 157996
rect 248750 157936 248755 157992
rect 217244 157932 217250 157934
rect 238753 157931 238819 157934
rect 248638 157932 248644 157934
rect 248708 157932 248755 157936
rect 251398 157932 251404 157996
rect 251468 157994 251474 157996
rect 252093 157994 252159 157997
rect 251468 157992 252159 157994
rect 251468 157936 252098 157992
rect 252154 157936 252159 157992
rect 251468 157934 252159 157936
rect 251468 157932 251474 157934
rect 248689 157931 248755 157932
rect 252093 157931 252159 157934
rect 253422 157932 253428 157996
rect 253492 157994 253498 157996
rect 253565 157994 253631 157997
rect 253492 157992 253631 157994
rect 253492 157936 253570 157992
rect 253626 157936 253631 157992
rect 253492 157934 253631 157936
rect 253492 157932 253498 157934
rect 253565 157931 253631 157934
rect 261702 157932 261708 157996
rect 261772 157994 261778 157996
rect 261937 157994 262003 157997
rect 261772 157992 262003 157994
rect 261772 157936 261942 157992
rect 261998 157936 262003 157992
rect 261772 157934 262003 157936
rect 261772 157932 261778 157934
rect 261937 157931 262003 157934
rect 266486 157932 266492 157996
rect 266556 157994 266562 157996
rect 266721 157994 266787 157997
rect 266556 157992 266787 157994
rect 266556 157936 266726 157992
rect 266782 157936 266787 157992
rect 266556 157934 266787 157936
rect 266556 157932 266562 157934
rect 266721 157931 266787 157934
rect 268326 157932 268332 157996
rect 268396 157994 268402 157996
rect 268929 157994 268995 157997
rect 268396 157992 268995 157994
rect 268396 157936 268934 157992
rect 268990 157936 268995 157992
rect 268396 157934 268995 157936
rect 268396 157932 268402 157934
rect 268929 157931 268995 157934
rect 345657 157994 345723 157997
rect 359641 157994 359707 157997
rect 345657 157992 359707 157994
rect 345657 157936 345662 157992
rect 345718 157936 359646 157992
rect 359702 157936 359707 157992
rect 345657 157934 359707 157936
rect 345657 157931 345723 157934
rect 359641 157931 359707 157934
rect 214649 157858 214715 157861
rect 223573 157858 223639 157861
rect 214649 157856 223639 157858
rect 214649 157800 214654 157856
rect 214710 157800 223578 157856
rect 223634 157800 223639 157856
rect 214649 157798 223639 157800
rect 214649 157795 214715 157798
rect 223573 157795 223639 157798
rect 237230 157796 237236 157860
rect 237300 157858 237306 157860
rect 366265 157858 366331 157861
rect 237300 157856 366331 157858
rect 237300 157800 366270 157856
rect 366326 157800 366331 157856
rect 237300 157798 366331 157800
rect 237300 157796 237306 157798
rect 366265 157795 366331 157798
rect 263910 157660 263916 157724
rect 263980 157722 263986 157724
rect 264421 157722 264487 157725
rect 263980 157720 264487 157722
rect 263980 157664 264426 157720
rect 264482 157664 264487 157720
rect 263980 157662 264487 157664
rect 263980 157660 263986 157662
rect 264421 157659 264487 157662
rect 265382 157660 265388 157724
rect 265452 157722 265458 157724
rect 265985 157722 266051 157725
rect 265452 157720 266051 157722
rect 265452 157664 265990 157720
rect 266046 157664 266051 157720
rect 265452 157662 266051 157664
rect 265452 157660 265458 157662
rect 265985 157659 266051 157662
rect 273662 157660 273668 157724
rect 273732 157722 273738 157724
rect 274449 157722 274515 157725
rect 273732 157720 274515 157722
rect 273732 157664 274454 157720
rect 274510 157664 274515 157720
rect 273732 157662 274515 157664
rect 273732 157660 273738 157662
rect 274449 157659 274515 157662
rect 278446 157660 278452 157724
rect 278516 157722 278522 157724
rect 278681 157722 278747 157725
rect 278516 157720 278747 157722
rect 278516 157664 278686 157720
rect 278742 157664 278747 157720
rect 278516 157662 278747 157664
rect 278516 157660 278522 157662
rect 278681 157659 278747 157662
rect 283598 157660 283604 157724
rect 283668 157722 283674 157724
rect 284109 157722 284175 157725
rect 283668 157720 284175 157722
rect 283668 157664 284114 157720
rect 284170 157664 284175 157720
rect 283668 157662 284175 157664
rect 283668 157660 283674 157662
rect 284109 157659 284175 157662
rect 288249 157588 288315 157589
rect 293585 157588 293651 157589
rect 288198 157586 288204 157588
rect 288158 157526 288204 157586
rect 288268 157584 288315 157588
rect 293534 157586 293540 157588
rect 288310 157528 288315 157584
rect 288198 157524 288204 157526
rect 288268 157524 288315 157528
rect 293494 157526 293540 157586
rect 293604 157584 293651 157588
rect 293646 157528 293651 157584
rect 293534 157524 293540 157526
rect 293604 157524 293651 157528
rect 288249 157523 288315 157524
rect 293585 157523 293651 157524
rect 253657 157452 253723 157453
rect 241830 157388 241836 157452
rect 241900 157388 241906 157452
rect 245510 157388 245516 157452
rect 245580 157388 245586 157452
rect 253606 157450 253612 157452
rect 253566 157390 253612 157450
rect 253676 157448 253723 157452
rect 253718 157392 253723 157448
rect 253606 157388 253612 157390
rect 253676 157388 253723 157392
rect 263542 157388 263548 157452
rect 263612 157450 263618 157452
rect 263961 157450 264027 157453
rect 263612 157448 264027 157450
rect 263612 157392 263966 157448
rect 264022 157392 264027 157448
rect 263612 157390 264027 157392
rect 263612 157388 263618 157390
rect 241838 156906 241898 157388
rect 245518 157314 245578 157388
rect 253657 157387 253723 157388
rect 263961 157387 264027 157390
rect 253197 157314 253263 157317
rect 373165 157314 373231 157317
rect 245518 157254 248430 157314
rect 248370 157178 248430 157254
rect 253197 157312 373231 157314
rect 253197 157256 253202 157312
rect 253258 157256 373170 157312
rect 373226 157256 373231 157312
rect 253197 157254 373231 157256
rect 253197 157251 253263 157254
rect 373165 157251 373231 157254
rect 368565 157178 368631 157181
rect 248370 157176 368631 157178
rect 248370 157120 368570 157176
rect 368626 157120 368631 157176
rect 248370 157118 368631 157120
rect 368565 157115 368631 157118
rect 247718 156980 247724 157044
rect 247788 157042 247794 157044
rect 369025 157042 369091 157045
rect 247788 157040 369091 157042
rect 247788 156984 369030 157040
rect 369086 156984 369091 157040
rect 247788 156982 369091 156984
rect 247788 156980 247794 156982
rect 369025 156979 369091 156982
rect 253197 156906 253263 156909
rect 370313 156906 370379 156909
rect 241838 156904 253263 156906
rect 241838 156848 253202 156904
rect 253258 156848 253263 156904
rect 241838 156846 253263 156848
rect 253197 156843 253263 156846
rect 258030 156904 370379 156906
rect 258030 156848 370318 156904
rect 370374 156848 370379 156904
rect 258030 156846 370379 156848
rect 252369 156770 252435 156773
rect 258030 156770 258090 156846
rect 370313 156843 370379 156846
rect 252369 156768 258090 156770
rect 252369 156712 252374 156768
rect 252430 156712 258090 156768
rect 252369 156710 258090 156712
rect 252369 156707 252435 156710
rect 246849 155954 246915 155957
rect 370037 155954 370103 155957
rect 246849 155952 370103 155954
rect 246849 155896 246854 155952
rect 246910 155896 370042 155952
rect 370098 155896 370103 155952
rect 246849 155894 370103 155896
rect 246849 155891 246915 155894
rect 370037 155891 370103 155894
rect 248689 155818 248755 155821
rect 370129 155818 370195 155821
rect 248689 155816 370195 155818
rect 248689 155760 248694 155816
rect 248750 155760 370134 155816
rect 370190 155760 370195 155816
rect 248689 155758 370195 155760
rect 248689 155755 248755 155758
rect 370129 155755 370195 155758
rect 293953 155546 294019 155549
rect 362309 155546 362375 155549
rect 293953 155544 362375 155546
rect 293953 155488 293958 155544
rect 294014 155488 362314 155544
rect 362370 155488 362375 155544
rect 293953 155486 362375 155488
rect 293953 155483 294019 155486
rect 362309 155483 362375 155486
rect 216990 155348 216996 155412
rect 217060 155410 217066 155412
rect 251265 155410 251331 155413
rect 217060 155408 251331 155410
rect 217060 155352 251270 155408
rect 251326 155352 251331 155408
rect 217060 155350 251331 155352
rect 217060 155348 217066 155350
rect 251265 155347 251331 155350
rect 292573 155410 292639 155413
rect 368422 155410 368428 155412
rect 292573 155408 368428 155410
rect 292573 155352 292578 155408
rect 292634 155352 368428 155408
rect 292573 155350 368428 155352
rect 292573 155347 292639 155350
rect 368422 155348 368428 155350
rect 368492 155348 368498 155412
rect 210785 155274 210851 155277
rect 269113 155274 269179 155277
rect 210785 155272 269179 155274
rect 210785 155216 210790 155272
rect 210846 155216 269118 155272
rect 269174 155216 269179 155272
rect 210785 155214 269179 155216
rect 210785 155211 210851 155214
rect 269113 155211 269179 155214
rect 291193 155274 291259 155277
rect 367921 155274 367987 155277
rect 291193 155272 367987 155274
rect 291193 155216 291198 155272
rect 291254 155216 367926 155272
rect 367982 155216 367987 155272
rect 291193 155214 367987 155216
rect 291193 155211 291259 155214
rect 367921 155211 367987 155214
rect 580625 152690 580691 152693
rect 583520 152690 584960 152780
rect 580625 152688 584960 152690
rect 580625 152632 580630 152688
rect 580686 152632 584960 152688
rect 580625 152630 584960 152632
rect 580625 152627 580691 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3509 149834 3575 149837
rect -960 149832 3575 149834
rect -960 149776 3514 149832
rect 3570 149776 3575 149832
rect -960 149774 3575 149776
rect -960 149684 480 149774
rect 3509 149771 3575 149774
rect 580533 139362 580599 139365
rect 583520 139362 584960 139452
rect 580533 139360 584960 139362
rect 580533 139304 580538 139360
rect 580594 139304 584960 139360
rect 580533 139302 584960 139304
rect 580533 139299 580599 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 583520 126034 584960 126124
rect 583342 125974 584960 126034
rect 583342 125898 583402 125974
rect 583520 125898 584960 125974
rect 583342 125884 584960 125898
rect 583342 125838 583586 125884
rect 368974 125564 368980 125628
rect 369044 125626 369050 125628
rect 583526 125626 583586 125838
rect 369044 125566 583586 125626
rect 369044 125564 369050 125566
rect -960 123572 480 123812
rect 580441 112842 580507 112845
rect 583520 112842 584960 112932
rect 580441 112840 584960 112842
rect 580441 112784 580446 112840
rect 580502 112784 584960 112840
rect 580441 112782 584960 112784
rect 580441 112779 580507 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 367870 99452 367876 99516
rect 367940 99514 367946 99516
rect 583520 99514 584960 99604
rect 367940 99454 584960 99514
rect 367940 99452 367946 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 583520 86186 584960 86276
rect 583342 86126 584960 86186
rect 583342 86050 583402 86126
rect 583520 86050 584960 86126
rect 583342 86036 584960 86050
rect 583342 85990 583586 86036
rect 367686 85580 367692 85644
rect 367756 85642 367762 85644
rect 583526 85642 583586 85990
rect 367756 85582 583586 85642
rect 367756 85580 367762 85582
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 583520 72994 584960 73084
rect 583342 72934 584960 72994
rect 583342 72858 583402 72934
rect 583520 72858 584960 72934
rect 583342 72844 584960 72858
rect 583342 72798 583586 72844
rect 362534 71844 362540 71908
rect 362604 71906 362610 71908
rect 583526 71906 583586 72798
rect 362604 71846 583586 71906
rect 362604 71844 362610 71846
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 583520 46338 584960 46428
rect 583342 46278 584960 46338
rect 583342 46202 583402 46278
rect 583520 46202 584960 46278
rect 583342 46188 584960 46202
rect 583342 46142 583586 46188
rect -960 45522 480 45612
rect 364926 45596 364932 45660
rect 364996 45658 365002 45660
rect 583526 45658 583586 46142
rect 364996 45598 583586 45658
rect 364996 45596 365002 45598
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 579613 33146 579679 33149
rect 583520 33146 584960 33236
rect 579613 33144 584960 33146
rect 579613 33088 579618 33144
rect 579674 33088 584960 33144
rect 579613 33086 584960 33088
rect 579613 33083 579679 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 580349 19818 580415 19821
rect 583520 19818 584960 19908
rect 580349 19816 584960 19818
rect 580349 19760 580354 19816
rect 580410 19760 584960 19816
rect 580349 19758 584960 19760
rect 580349 19755 580415 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 350441 6898 350507 6901
rect 363454 6898 363460 6900
rect 350441 6896 363460 6898
rect 350441 6840 350446 6896
rect 350502 6840 363460 6896
rect 350441 6838 363460 6840
rect 350441 6835 350507 6838
rect 363454 6836 363460 6838
rect 363524 6836 363530 6900
rect 351637 6762 351703 6765
rect 365805 6762 365871 6765
rect 351637 6760 365871 6762
rect 351637 6704 351642 6760
rect 351698 6704 365810 6760
rect 365866 6704 365871 6760
rect 351637 6702 365871 6704
rect 351637 6699 351703 6702
rect 365805 6699 365871 6702
rect 348049 6626 348115 6629
rect 363270 6626 363276 6628
rect 348049 6624 363276 6626
rect -960 6490 480 6580
rect 348049 6568 348054 6624
rect 348110 6568 363276 6624
rect 348049 6566 363276 6568
rect 348049 6563 348115 6566
rect 363270 6564 363276 6566
rect 363340 6564 363346 6628
rect 580257 6626 580323 6629
rect 583520 6626 584960 6716
rect 580257 6624 584960 6626
rect 580257 6568 580262 6624
rect 580318 6568 584960 6624
rect 580257 6566 584960 6568
rect 580257 6563 580323 6566
rect 344553 6490 344619 6493
rect 363086 6490 363092 6492
rect -960 6430 674 6490
rect -960 6354 480 6430
rect 614 6354 674 6430
rect 344553 6488 363092 6490
rect 344553 6432 344558 6488
rect 344614 6432 363092 6488
rect 344553 6430 363092 6432
rect 344553 6427 344619 6430
rect 363086 6428 363092 6430
rect 363156 6428 363162 6492
rect 583520 6476 584960 6566
rect -960 6340 674 6354
rect 246 6294 674 6340
rect 323301 6354 323367 6357
rect 358118 6354 358124 6356
rect 323301 6352 358124 6354
rect 323301 6296 323306 6352
rect 323362 6296 358124 6352
rect 323301 6294 358124 6296
rect 246 5810 306 6294
rect 323301 6291 323367 6294
rect 358118 6292 358124 6294
rect 358188 6292 358194 6356
rect 320909 6218 320975 6221
rect 367318 6218 367324 6220
rect 320909 6216 367324 6218
rect 320909 6160 320914 6216
rect 320970 6160 367324 6216
rect 320909 6158 367324 6160
rect 320909 6155 320975 6158
rect 367318 6156 367324 6158
rect 367388 6156 367394 6220
rect 246 5750 6930 5810
rect 6870 5674 6930 5750
rect 215886 5674 215892 5676
rect 6870 5614 215892 5674
rect 215886 5612 215892 5614
rect 215956 5612 215962 5676
rect 343357 4042 343423 4045
rect 356421 4042 356487 4045
rect 343357 4040 356487 4042
rect 343357 3984 343362 4040
rect 343418 3984 356426 4040
rect 356482 3984 356487 4040
rect 343357 3982 356487 3984
rect 343357 3979 343423 3982
rect 356421 3979 356487 3982
rect 356605 4042 356671 4045
rect 360326 4042 360332 4044
rect 356605 4040 360332 4042
rect 356605 3984 356610 4040
rect 356666 3984 360332 4040
rect 356605 3982 360332 3984
rect 356605 3979 356671 3982
rect 360326 3980 360332 3982
rect 360396 3980 360402 4044
rect 335077 3906 335143 3909
rect 359406 3906 359412 3908
rect 335077 3904 359412 3906
rect 335077 3848 335082 3904
rect 335138 3848 359412 3904
rect 335077 3846 359412 3848
rect 335077 3843 335143 3846
rect 359406 3844 359412 3846
rect 359476 3844 359482 3908
rect 331581 3770 331647 3773
rect 356605 3770 356671 3773
rect 359038 3770 359044 3772
rect 331581 3768 356671 3770
rect 331581 3712 331586 3768
rect 331642 3712 356610 3768
rect 356666 3712 356671 3768
rect 331581 3710 356671 3712
rect 331581 3707 331647 3710
rect 356605 3707 356671 3710
rect 356838 3710 359044 3770
rect 327993 3634 328059 3637
rect 356697 3634 356763 3637
rect 327993 3632 356763 3634
rect 327993 3576 327998 3632
rect 328054 3576 356702 3632
rect 356758 3576 356763 3632
rect 327993 3574 356763 3576
rect 327993 3571 328059 3574
rect 356697 3571 356763 3574
rect 214465 3498 214531 3501
rect 215150 3498 215156 3500
rect 214465 3496 215156 3498
rect 214465 3440 214470 3496
rect 214526 3440 215156 3496
rect 214465 3438 215156 3440
rect 214465 3435 214531 3438
rect 215150 3436 215156 3438
rect 215220 3436 215226 3500
rect 215661 3498 215727 3501
rect 216438 3498 216444 3500
rect 215661 3496 216444 3498
rect 215661 3440 215666 3496
rect 215722 3440 216444 3496
rect 215661 3438 216444 3440
rect 215661 3435 215727 3438
rect 216438 3436 216444 3438
rect 216508 3436 216514 3500
rect 216857 3498 216923 3501
rect 217542 3498 217548 3500
rect 216857 3496 217548 3498
rect 216857 3440 216862 3496
rect 216918 3440 217548 3496
rect 216857 3438 217548 3440
rect 216857 3435 216923 3438
rect 217542 3436 217548 3438
rect 217612 3436 217618 3500
rect 218646 3436 218652 3500
rect 218716 3498 218722 3500
rect 219249 3498 219315 3501
rect 218716 3496 219315 3498
rect 218716 3440 219254 3496
rect 219310 3440 219315 3496
rect 218716 3438 219315 3440
rect 218716 3436 218722 3438
rect 219249 3435 219315 3438
rect 325601 3498 325667 3501
rect 356838 3498 356898 3710
rect 359038 3708 359044 3710
rect 359108 3708 359114 3772
rect 357525 3634 357591 3637
rect 358486 3634 358492 3636
rect 357525 3632 358492 3634
rect 357525 3576 357530 3632
rect 357586 3576 358492 3632
rect 357525 3574 358492 3576
rect 357525 3571 357591 3574
rect 358486 3572 358492 3574
rect 358556 3572 358562 3636
rect 365662 3572 365668 3636
rect 365732 3634 365738 3636
rect 365805 3634 365871 3637
rect 365732 3632 365871 3634
rect 365732 3576 365810 3632
rect 365866 3576 365871 3632
rect 365732 3574 365871 3576
rect 365732 3572 365738 3574
rect 365805 3571 365871 3574
rect 325601 3496 356898 3498
rect 325601 3440 325606 3496
rect 325662 3440 356898 3496
rect 325601 3438 356898 3440
rect 325601 3435 325667 3438
rect 358302 3436 358308 3500
rect 358372 3498 358378 3500
rect 358721 3498 358787 3501
rect 358372 3496 358787 3498
rect 358372 3440 358726 3496
rect 358782 3440 358787 3496
rect 358372 3438 358787 3440
rect 358372 3436 358378 3438
rect 358721 3435 358787 3438
rect 358854 3436 358860 3500
rect 358924 3498 358930 3500
rect 359917 3498 359983 3501
rect 358924 3496 359983 3498
rect 358924 3440 359922 3496
rect 359978 3440 359983 3496
rect 358924 3438 359983 3440
rect 358924 3436 358930 3438
rect 359917 3435 359983 3438
rect 360142 3436 360148 3500
rect 360212 3498 360218 3500
rect 361113 3498 361179 3501
rect 360212 3496 361179 3498
rect 360212 3440 361118 3496
rect 361174 3440 361179 3496
rect 360212 3438 361179 3440
rect 360212 3436 360218 3438
rect 361113 3435 361179 3438
rect 362902 3436 362908 3500
rect 362972 3498 362978 3500
rect 363505 3498 363571 3501
rect 362972 3496 363571 3498
rect 362972 3440 363510 3496
rect 363566 3440 363571 3496
rect 362972 3438 363571 3440
rect 362972 3436 362978 3438
rect 363505 3435 363571 3438
rect 364374 3436 364380 3500
rect 364444 3498 364450 3500
rect 364609 3498 364675 3501
rect 364444 3496 364675 3498
rect 364444 3440 364614 3496
rect 364670 3440 364675 3496
rect 364444 3438 364675 3440
rect 364444 3436 364450 3438
rect 364609 3435 364675 3438
rect 365846 3436 365852 3500
rect 365916 3498 365922 3500
rect 367001 3498 367067 3501
rect 365916 3496 367067 3498
rect 365916 3440 367006 3496
rect 367062 3440 367067 3496
rect 365916 3438 367067 3440
rect 365916 3436 365922 3438
rect 367001 3435 367067 3438
rect 367134 3436 367140 3500
rect 367204 3498 367210 3500
rect 368197 3498 368263 3501
rect 367204 3496 368263 3498
rect 367204 3440 368202 3496
rect 368258 3440 368263 3496
rect 367204 3438 368263 3440
rect 367204 3436 367210 3438
rect 368197 3435 368263 3438
rect 369894 3436 369900 3500
rect 369964 3498 369970 3500
rect 370589 3498 370655 3501
rect 369964 3496 370655 3498
rect 369964 3440 370594 3496
rect 370650 3440 370655 3496
rect 369964 3438 370655 3440
rect 369964 3436 369970 3438
rect 370589 3435 370655 3438
rect 205081 3362 205147 3365
rect 214414 3362 214420 3364
rect 205081 3360 214420 3362
rect 205081 3304 205086 3360
rect 205142 3304 214420 3360
rect 205081 3302 214420 3304
rect 205081 3299 205147 3302
rect 214414 3300 214420 3302
rect 214484 3300 214490 3364
rect 215201 3362 215267 3365
rect 222745 3362 222811 3365
rect 215201 3360 222811 3362
rect 215201 3304 215206 3360
rect 215262 3304 222750 3360
rect 222806 3304 222811 3360
rect 215201 3302 222811 3304
rect 215201 3299 215267 3302
rect 222745 3299 222811 3302
rect 324405 3362 324471 3365
rect 359222 3362 359228 3364
rect 324405 3360 359228 3362
rect 324405 3304 324410 3360
rect 324466 3304 359228 3360
rect 324405 3302 359228 3304
rect 324405 3299 324471 3302
rect 359222 3300 359228 3302
rect 359292 3300 359298 3364
rect 369158 3300 369164 3364
rect 369228 3362 369234 3364
rect 379973 3362 380039 3365
rect 369228 3360 380039 3362
rect 369228 3304 379978 3360
rect 380034 3304 380039 3360
rect 369228 3302 380039 3304
rect 369228 3300 369234 3302
rect 379973 3299 380039 3302
rect 346945 3226 347011 3229
rect 356697 3226 356763 3229
rect 360510 3226 360516 3228
rect 346945 3224 354690 3226
rect 346945 3168 346950 3224
rect 347006 3168 354690 3224
rect 346945 3166 354690 3168
rect 346945 3163 347011 3166
rect 354630 3090 354690 3166
rect 356697 3224 360516 3226
rect 356697 3168 356702 3224
rect 356758 3168 360516 3224
rect 356697 3166 360516 3168
rect 356697 3163 356763 3166
rect 360510 3164 360516 3166
rect 360580 3164 360586 3228
rect 364558 3090 364564 3092
rect 354630 3030 364564 3090
rect 364558 3028 364564 3030
rect 364628 3028 364634 3092
rect 356421 2954 356487 2957
rect 363137 2954 363203 2957
rect 356421 2952 363203 2954
rect 356421 2896 356426 2952
rect 356482 2896 363142 2952
rect 363198 2896 363203 2952
rect 356421 2894 363203 2896
rect 356421 2891 356487 2894
rect 363137 2891 363203 2894
<< via3 >>
rect 238340 477260 238404 477324
rect 241836 477124 241900 477188
rect 253428 477124 253492 477188
rect 256188 476988 256252 477052
rect 320956 476988 321020 477052
rect 239628 476852 239692 476916
rect 240548 476852 240612 476916
rect 236132 476716 236196 476780
rect 258028 476716 258092 476780
rect 308628 476716 308692 476780
rect 313412 476716 313476 476780
rect 265940 476580 266004 476644
rect 270908 476580 270972 476644
rect 261156 476444 261220 476508
rect 273668 476444 273732 476508
rect 318564 476444 318628 476508
rect 323348 476444 323412 476508
rect 325924 476444 325988 476508
rect 244228 476308 244292 476372
rect 247724 476308 247788 476372
rect 250116 476308 250180 476372
rect 251404 476308 251468 476372
rect 259500 476308 259564 476372
rect 263548 476308 263612 476372
rect 266492 476308 266556 476372
rect 268332 476308 268396 476372
rect 273300 476308 273364 476372
rect 276060 476308 276124 476372
rect 278084 476308 278148 476372
rect 311020 476308 311084 476372
rect 237236 476232 237300 476236
rect 237236 476176 237250 476232
rect 237250 476176 237300 476232
rect 237236 476172 237300 476176
rect 243124 476172 243188 476236
rect 245516 476232 245580 476236
rect 245516 476176 245530 476232
rect 245530 476176 245580 476232
rect 245516 476172 245580 476176
rect 246620 476172 246684 476236
rect 248276 476232 248340 476236
rect 248276 476176 248326 476232
rect 248326 476176 248340 476232
rect 248276 476172 248340 476176
rect 248644 476172 248708 476236
rect 250852 476172 250916 476236
rect 252324 476172 252388 476236
rect 253612 476172 253676 476236
rect 254532 476172 254596 476236
rect 255820 476172 255884 476236
rect 257108 476172 257172 476236
rect 258580 476172 258644 476236
rect 260604 476172 260668 476236
rect 261708 476172 261772 476236
rect 262812 476172 262876 476236
rect 263916 476172 263980 476236
rect 265388 476172 265452 476236
rect 267596 476232 267660 476236
rect 267596 476176 267610 476232
rect 267610 476176 267660 476232
rect 267596 476172 267660 476176
rect 268700 476172 268764 476236
rect 269804 476172 269868 476236
rect 271276 476172 271340 476236
rect 272196 476172 272260 476236
rect 274404 476232 274468 476236
rect 274404 476176 274418 476232
rect 274418 476176 274468 476232
rect 274404 476172 274468 476176
rect 275876 476232 275940 476236
rect 275876 476176 275926 476232
rect 275926 476176 275940 476232
rect 275876 476172 275940 476176
rect 276980 476172 277044 476236
rect 278452 476172 278516 476236
rect 279188 476172 279252 476236
rect 281028 476172 281092 476236
rect 283604 476172 283668 476236
rect 285996 476172 286060 476236
rect 288204 476172 288268 476236
rect 290964 476172 291028 476236
rect 293540 476172 293604 476236
rect 295932 476172 295996 476236
rect 298508 476172 298572 476236
rect 300900 476172 300964 476236
rect 303476 476232 303540 476236
rect 303476 476176 303526 476232
rect 303526 476176 303540 476232
rect 303476 476172 303540 476176
rect 306052 476172 306116 476236
rect 315804 476172 315868 476236
rect 369348 445844 369412 445908
rect 367876 445708 367940 445772
rect 216076 444892 216140 444956
rect 214604 444756 214668 444820
rect 364932 444620 364996 444684
rect 368980 444484 369044 444548
rect 367692 444348 367756 444412
rect 362540 443260 362604 443324
rect 215892 441764 215956 441828
rect 362724 441628 362788 441692
rect 232084 374036 232148 374100
rect 231900 373220 231964 373284
rect 232084 311204 232148 311268
rect 232084 310388 232148 310452
rect 231900 310252 231964 310316
rect 232452 309708 232516 309772
rect 169340 308484 169404 308548
rect 218836 306172 218900 306236
rect 219020 306036 219084 306100
rect 219204 305900 219268 305964
rect 217364 305764 217428 305828
rect 217180 305628 217244 305692
rect 369900 303452 369964 303516
rect 216260 303316 216324 303380
rect 215156 303180 215220 303244
rect 169524 301548 169588 301612
rect 169156 301140 169220 301204
rect 368428 300052 368492 300116
rect 169340 299100 169404 299164
rect 169156 298012 169220 298076
rect 169524 297876 169588 297940
rect 216996 297740 217060 297804
rect 367140 286316 367204 286380
rect 214420 284820 214484 284884
rect 364380 258708 364444 258772
rect 216444 255852 216508 255916
rect 365668 254628 365732 254692
rect 369164 254492 369228 254556
rect 365852 253132 365916 253196
rect 358860 251908 358924 251972
rect 362908 251772 362972 251836
rect 358124 250820 358188 250884
rect 363092 250684 363156 250748
rect 363276 250548 363340 250612
rect 217548 250412 217612 250476
rect 367324 250412 367388 250476
rect 360148 248236 360212 248300
rect 359044 248100 359108 248164
rect 363460 247964 363524 248028
rect 364748 247828 364812 247892
rect 364564 247692 364628 247756
rect 358676 245516 358740 245580
rect 360700 245380 360764 245444
rect 359412 245244 359476 245308
rect 359228 245108 359292 245172
rect 360516 244972 360580 245036
rect 360332 244836 360396 244900
rect 358308 244700 358372 244764
rect 358492 243476 358556 243540
rect 362724 231916 362788 231980
rect 369348 218044 369412 218108
rect 216076 213964 216140 214028
rect 218652 193216 218716 193220
rect 218652 193160 218666 193216
rect 218666 193160 218716 193216
rect 218652 193156 218716 193160
rect 214604 162828 214668 162892
rect 258494 159896 258558 159900
rect 258494 159840 258538 159896
rect 258538 159840 258558 159896
rect 258494 159836 258558 159840
rect 275766 159836 275830 159900
rect 276990 159896 277054 159900
rect 276990 159840 277030 159896
rect 277030 159840 277054 159896
rect 276990 159836 277054 159840
rect 278078 159896 278142 159900
rect 278078 159840 278134 159896
rect 278134 159840 278142 159896
rect 278078 159836 278142 159840
rect 279166 159836 279230 159900
rect 300926 159760 300990 159764
rect 300926 159704 300950 159760
rect 300950 159704 300990 159760
rect 300926 159700 300990 159704
rect 255910 159624 255974 159628
rect 255910 159568 255962 159624
rect 255962 159568 255974 159624
rect 255910 159564 255974 159568
rect 271006 159624 271070 159628
rect 271006 159568 271050 159624
rect 271050 159568 271070 159624
rect 271006 159564 271070 159568
rect 274406 159624 274470 159628
rect 274406 159568 274454 159624
rect 274454 159568 274470 159624
rect 274406 159564 274470 159568
rect 254532 159156 254596 159220
rect 250852 159020 250916 159084
rect 243124 158884 243188 158948
rect 236132 158748 236196 158812
rect 358676 158748 358740 158812
rect 360700 158748 360764 158812
rect 364748 158748 364812 158812
rect 218836 158612 218900 158676
rect 238156 158672 238220 158676
rect 238156 158616 238170 158672
rect 238170 158616 238220 158672
rect 238156 158612 238220 158616
rect 239628 158672 239692 158676
rect 239628 158616 239642 158672
rect 239642 158616 239692 158672
rect 239628 158612 239692 158616
rect 240548 158612 240612 158676
rect 248276 158672 248340 158676
rect 248276 158616 248326 158672
rect 248326 158616 248340 158672
rect 248276 158612 248340 158616
rect 250116 158672 250180 158676
rect 250116 158616 250166 158672
rect 250166 158616 250180 158672
rect 250116 158612 250180 158616
rect 256004 158612 256068 158676
rect 257108 158672 257172 158676
rect 257108 158616 257158 158672
rect 257158 158616 257172 158672
rect 257108 158612 257172 158616
rect 258212 158612 258276 158676
rect 259500 158672 259564 158676
rect 259500 158616 259550 158672
rect 259550 158616 259564 158672
rect 259500 158612 259564 158616
rect 261156 158612 261220 158676
rect 262812 158672 262876 158676
rect 262812 158616 262862 158672
rect 262862 158616 262876 158672
rect 262812 158612 262876 158616
rect 265940 158672 266004 158676
rect 265940 158616 265990 158672
rect 265990 158616 266004 158672
rect 265940 158612 266004 158616
rect 267596 158672 267660 158676
rect 267596 158616 267646 158672
rect 267646 158616 267660 158672
rect 267596 158612 267660 158616
rect 268700 158672 268764 158676
rect 268700 158616 268750 158672
rect 268750 158616 268764 158672
rect 268700 158612 268764 158616
rect 269804 158612 269868 158676
rect 271092 158672 271156 158676
rect 271092 158616 271142 158672
rect 271142 158616 271156 158672
rect 271092 158612 271156 158616
rect 272196 158672 272260 158676
rect 272196 158616 272246 158672
rect 272246 158616 272260 158672
rect 272196 158612 272260 158616
rect 298508 158612 298572 158676
rect 303476 158672 303540 158676
rect 303476 158616 303526 158672
rect 303526 158616 303540 158672
rect 303476 158612 303540 158616
rect 306052 158672 306116 158676
rect 306052 158616 306102 158672
rect 306102 158616 306116 158672
rect 306052 158612 306116 158616
rect 308628 158672 308692 158676
rect 308628 158616 308678 158672
rect 308678 158616 308692 158672
rect 308628 158612 308692 158616
rect 313412 158672 313476 158676
rect 313412 158616 313462 158672
rect 313462 158616 313476 158672
rect 313412 158612 313476 158616
rect 315804 158672 315868 158676
rect 315804 158616 315854 158672
rect 315854 158616 315868 158672
rect 315804 158612 315868 158616
rect 318564 158672 318628 158676
rect 318564 158616 318614 158672
rect 318614 158616 318628 158672
rect 318564 158612 318628 158616
rect 320956 158612 321020 158676
rect 323348 158672 323412 158676
rect 323348 158616 323398 158672
rect 323398 158616 323412 158672
rect 323348 158612 323412 158616
rect 325924 158672 325988 158676
rect 325924 158616 325974 158672
rect 325974 158616 325988 158672
rect 325924 158612 325988 158616
rect 219020 158476 219084 158540
rect 252324 158536 252388 158540
rect 252324 158480 252374 158536
rect 252374 158480 252388 158536
rect 252324 158476 252388 158480
rect 260604 158536 260668 158540
rect 260604 158480 260654 158536
rect 260654 158480 260668 158536
rect 260604 158476 260668 158480
rect 276060 158536 276124 158540
rect 276060 158480 276110 158536
rect 276110 158480 276124 158536
rect 276060 158476 276124 158480
rect 281028 158476 281092 158540
rect 285996 158476 286060 158540
rect 219204 158340 219268 158404
rect 273300 158400 273364 158404
rect 273300 158344 273350 158400
rect 273350 158344 273364 158400
rect 273300 158340 273364 158344
rect 290964 158400 291028 158404
rect 290964 158344 291014 158400
rect 291014 158344 291028 158400
rect 290964 158340 291028 158344
rect 295932 158340 295996 158404
rect 216260 158204 216324 158268
rect 244228 158204 244292 158268
rect 311020 158204 311084 158268
rect 217364 158068 217428 158132
rect 246620 158068 246684 158132
rect 217180 157932 217244 157996
rect 248644 157992 248708 157996
rect 248644 157936 248694 157992
rect 248694 157936 248708 157992
rect 248644 157932 248708 157936
rect 251404 157932 251468 157996
rect 253428 157932 253492 157996
rect 261708 157932 261772 157996
rect 266492 157932 266556 157996
rect 268332 157932 268396 157996
rect 237236 157796 237300 157860
rect 263916 157660 263980 157724
rect 265388 157660 265452 157724
rect 273668 157660 273732 157724
rect 278452 157660 278516 157724
rect 283604 157660 283668 157724
rect 288204 157584 288268 157588
rect 288204 157528 288254 157584
rect 288254 157528 288268 157584
rect 288204 157524 288268 157528
rect 293540 157584 293604 157588
rect 293540 157528 293590 157584
rect 293590 157528 293604 157584
rect 293540 157524 293604 157528
rect 241836 157388 241900 157452
rect 245516 157388 245580 157452
rect 253612 157448 253676 157452
rect 253612 157392 253662 157448
rect 253662 157392 253676 157448
rect 253612 157388 253676 157392
rect 263548 157388 263612 157452
rect 247724 156980 247788 157044
rect 216996 155348 217060 155412
rect 368428 155348 368492 155412
rect 368980 125564 369044 125628
rect 367876 99452 367940 99516
rect 367692 85580 367756 85644
rect 362540 71844 362604 71908
rect 364932 45596 364996 45660
rect 363460 6836 363524 6900
rect 363276 6564 363340 6628
rect 363092 6428 363156 6492
rect 358124 6292 358188 6356
rect 367324 6156 367388 6220
rect 215892 5612 215956 5676
rect 360332 3980 360396 4044
rect 359412 3844 359476 3908
rect 215156 3436 215220 3500
rect 216444 3436 216508 3500
rect 217548 3436 217612 3500
rect 218652 3436 218716 3500
rect 359044 3708 359108 3772
rect 358492 3572 358556 3636
rect 365668 3572 365732 3636
rect 358308 3436 358372 3500
rect 358860 3436 358924 3500
rect 360148 3436 360212 3500
rect 362908 3436 362972 3500
rect 364380 3436 364444 3500
rect 365852 3436 365916 3500
rect 367140 3436 367204 3500
rect 369900 3436 369964 3500
rect 214420 3300 214484 3364
rect 359228 3300 359292 3364
rect 369164 3300 369228 3364
rect 360516 3164 360580 3228
rect 364564 3028 364628 3092
<< metal4 >>
rect -9036 711868 -8416 711900
rect -9036 711632 -9004 711868
rect -8768 711632 -8684 711868
rect -8448 711632 -8416 711868
rect -9036 711548 -8416 711632
rect -9036 711312 -9004 711548
rect -8768 711312 -8684 711548
rect -8448 711312 -8416 711548
rect -9036 682954 -8416 711312
rect -9036 682718 -9004 682954
rect -8768 682718 -8684 682954
rect -8448 682718 -8416 682954
rect -9036 682634 -8416 682718
rect -9036 682398 -9004 682634
rect -8768 682398 -8684 682634
rect -8448 682398 -8416 682634
rect -9036 646954 -8416 682398
rect -9036 646718 -9004 646954
rect -8768 646718 -8684 646954
rect -8448 646718 -8416 646954
rect -9036 646634 -8416 646718
rect -9036 646398 -9004 646634
rect -8768 646398 -8684 646634
rect -8448 646398 -8416 646634
rect -9036 610954 -8416 646398
rect -9036 610718 -9004 610954
rect -8768 610718 -8684 610954
rect -8448 610718 -8416 610954
rect -9036 610634 -8416 610718
rect -9036 610398 -9004 610634
rect -8768 610398 -8684 610634
rect -8448 610398 -8416 610634
rect -9036 574954 -8416 610398
rect -9036 574718 -9004 574954
rect -8768 574718 -8684 574954
rect -8448 574718 -8416 574954
rect -9036 574634 -8416 574718
rect -9036 574398 -9004 574634
rect -8768 574398 -8684 574634
rect -8448 574398 -8416 574634
rect -9036 538954 -8416 574398
rect -9036 538718 -9004 538954
rect -8768 538718 -8684 538954
rect -8448 538718 -8416 538954
rect -9036 538634 -8416 538718
rect -9036 538398 -9004 538634
rect -8768 538398 -8684 538634
rect -8448 538398 -8416 538634
rect -9036 502954 -8416 538398
rect -9036 502718 -9004 502954
rect -8768 502718 -8684 502954
rect -8448 502718 -8416 502954
rect -9036 502634 -8416 502718
rect -9036 502398 -9004 502634
rect -8768 502398 -8684 502634
rect -8448 502398 -8416 502634
rect -9036 466954 -8416 502398
rect -9036 466718 -9004 466954
rect -8768 466718 -8684 466954
rect -8448 466718 -8416 466954
rect -9036 466634 -8416 466718
rect -9036 466398 -9004 466634
rect -8768 466398 -8684 466634
rect -8448 466398 -8416 466634
rect -9036 430954 -8416 466398
rect -9036 430718 -9004 430954
rect -8768 430718 -8684 430954
rect -8448 430718 -8416 430954
rect -9036 430634 -8416 430718
rect -9036 430398 -9004 430634
rect -8768 430398 -8684 430634
rect -8448 430398 -8416 430634
rect -9036 394954 -8416 430398
rect -9036 394718 -9004 394954
rect -8768 394718 -8684 394954
rect -8448 394718 -8416 394954
rect -9036 394634 -8416 394718
rect -9036 394398 -9004 394634
rect -8768 394398 -8684 394634
rect -8448 394398 -8416 394634
rect -9036 358954 -8416 394398
rect -9036 358718 -9004 358954
rect -8768 358718 -8684 358954
rect -8448 358718 -8416 358954
rect -9036 358634 -8416 358718
rect -9036 358398 -9004 358634
rect -8768 358398 -8684 358634
rect -8448 358398 -8416 358634
rect -9036 322954 -8416 358398
rect -9036 322718 -9004 322954
rect -8768 322718 -8684 322954
rect -8448 322718 -8416 322954
rect -9036 322634 -8416 322718
rect -9036 322398 -9004 322634
rect -8768 322398 -8684 322634
rect -8448 322398 -8416 322634
rect -9036 286954 -8416 322398
rect -9036 286718 -9004 286954
rect -8768 286718 -8684 286954
rect -8448 286718 -8416 286954
rect -9036 286634 -8416 286718
rect -9036 286398 -9004 286634
rect -8768 286398 -8684 286634
rect -8448 286398 -8416 286634
rect -9036 250954 -8416 286398
rect -9036 250718 -9004 250954
rect -8768 250718 -8684 250954
rect -8448 250718 -8416 250954
rect -9036 250634 -8416 250718
rect -9036 250398 -9004 250634
rect -8768 250398 -8684 250634
rect -8448 250398 -8416 250634
rect -9036 214954 -8416 250398
rect -9036 214718 -9004 214954
rect -8768 214718 -8684 214954
rect -8448 214718 -8416 214954
rect -9036 214634 -8416 214718
rect -9036 214398 -9004 214634
rect -8768 214398 -8684 214634
rect -8448 214398 -8416 214634
rect -9036 178954 -8416 214398
rect -9036 178718 -9004 178954
rect -8768 178718 -8684 178954
rect -8448 178718 -8416 178954
rect -9036 178634 -8416 178718
rect -9036 178398 -9004 178634
rect -8768 178398 -8684 178634
rect -8448 178398 -8416 178634
rect -9036 142954 -8416 178398
rect -9036 142718 -9004 142954
rect -8768 142718 -8684 142954
rect -8448 142718 -8416 142954
rect -9036 142634 -8416 142718
rect -9036 142398 -9004 142634
rect -8768 142398 -8684 142634
rect -8448 142398 -8416 142634
rect -9036 106954 -8416 142398
rect -9036 106718 -9004 106954
rect -8768 106718 -8684 106954
rect -8448 106718 -8416 106954
rect -9036 106634 -8416 106718
rect -9036 106398 -9004 106634
rect -8768 106398 -8684 106634
rect -8448 106398 -8416 106634
rect -9036 70954 -8416 106398
rect -9036 70718 -9004 70954
rect -8768 70718 -8684 70954
rect -8448 70718 -8416 70954
rect -9036 70634 -8416 70718
rect -9036 70398 -9004 70634
rect -8768 70398 -8684 70634
rect -8448 70398 -8416 70634
rect -9036 34954 -8416 70398
rect -9036 34718 -9004 34954
rect -8768 34718 -8684 34954
rect -8448 34718 -8416 34954
rect -9036 34634 -8416 34718
rect -9036 34398 -9004 34634
rect -8768 34398 -8684 34634
rect -8448 34398 -8416 34634
rect -9036 -7376 -8416 34398
rect -8076 710908 -7456 710940
rect -8076 710672 -8044 710908
rect -7808 710672 -7724 710908
rect -7488 710672 -7456 710908
rect -8076 710588 -7456 710672
rect -8076 710352 -8044 710588
rect -7808 710352 -7724 710588
rect -7488 710352 -7456 710588
rect -8076 678454 -7456 710352
rect -8076 678218 -8044 678454
rect -7808 678218 -7724 678454
rect -7488 678218 -7456 678454
rect -8076 678134 -7456 678218
rect -8076 677898 -8044 678134
rect -7808 677898 -7724 678134
rect -7488 677898 -7456 678134
rect -8076 642454 -7456 677898
rect -8076 642218 -8044 642454
rect -7808 642218 -7724 642454
rect -7488 642218 -7456 642454
rect -8076 642134 -7456 642218
rect -8076 641898 -8044 642134
rect -7808 641898 -7724 642134
rect -7488 641898 -7456 642134
rect -8076 606454 -7456 641898
rect -8076 606218 -8044 606454
rect -7808 606218 -7724 606454
rect -7488 606218 -7456 606454
rect -8076 606134 -7456 606218
rect -8076 605898 -8044 606134
rect -7808 605898 -7724 606134
rect -7488 605898 -7456 606134
rect -8076 570454 -7456 605898
rect -8076 570218 -8044 570454
rect -7808 570218 -7724 570454
rect -7488 570218 -7456 570454
rect -8076 570134 -7456 570218
rect -8076 569898 -8044 570134
rect -7808 569898 -7724 570134
rect -7488 569898 -7456 570134
rect -8076 534454 -7456 569898
rect -8076 534218 -8044 534454
rect -7808 534218 -7724 534454
rect -7488 534218 -7456 534454
rect -8076 534134 -7456 534218
rect -8076 533898 -8044 534134
rect -7808 533898 -7724 534134
rect -7488 533898 -7456 534134
rect -8076 498454 -7456 533898
rect -8076 498218 -8044 498454
rect -7808 498218 -7724 498454
rect -7488 498218 -7456 498454
rect -8076 498134 -7456 498218
rect -8076 497898 -8044 498134
rect -7808 497898 -7724 498134
rect -7488 497898 -7456 498134
rect -8076 462454 -7456 497898
rect -8076 462218 -8044 462454
rect -7808 462218 -7724 462454
rect -7488 462218 -7456 462454
rect -8076 462134 -7456 462218
rect -8076 461898 -8044 462134
rect -7808 461898 -7724 462134
rect -7488 461898 -7456 462134
rect -8076 426454 -7456 461898
rect -8076 426218 -8044 426454
rect -7808 426218 -7724 426454
rect -7488 426218 -7456 426454
rect -8076 426134 -7456 426218
rect -8076 425898 -8044 426134
rect -7808 425898 -7724 426134
rect -7488 425898 -7456 426134
rect -8076 390454 -7456 425898
rect -8076 390218 -8044 390454
rect -7808 390218 -7724 390454
rect -7488 390218 -7456 390454
rect -8076 390134 -7456 390218
rect -8076 389898 -8044 390134
rect -7808 389898 -7724 390134
rect -7488 389898 -7456 390134
rect -8076 354454 -7456 389898
rect -8076 354218 -8044 354454
rect -7808 354218 -7724 354454
rect -7488 354218 -7456 354454
rect -8076 354134 -7456 354218
rect -8076 353898 -8044 354134
rect -7808 353898 -7724 354134
rect -7488 353898 -7456 354134
rect -8076 318454 -7456 353898
rect -8076 318218 -8044 318454
rect -7808 318218 -7724 318454
rect -7488 318218 -7456 318454
rect -8076 318134 -7456 318218
rect -8076 317898 -8044 318134
rect -7808 317898 -7724 318134
rect -7488 317898 -7456 318134
rect -8076 282454 -7456 317898
rect -8076 282218 -8044 282454
rect -7808 282218 -7724 282454
rect -7488 282218 -7456 282454
rect -8076 282134 -7456 282218
rect -8076 281898 -8044 282134
rect -7808 281898 -7724 282134
rect -7488 281898 -7456 282134
rect -8076 246454 -7456 281898
rect -8076 246218 -8044 246454
rect -7808 246218 -7724 246454
rect -7488 246218 -7456 246454
rect -8076 246134 -7456 246218
rect -8076 245898 -8044 246134
rect -7808 245898 -7724 246134
rect -7488 245898 -7456 246134
rect -8076 210454 -7456 245898
rect -8076 210218 -8044 210454
rect -7808 210218 -7724 210454
rect -7488 210218 -7456 210454
rect -8076 210134 -7456 210218
rect -8076 209898 -8044 210134
rect -7808 209898 -7724 210134
rect -7488 209898 -7456 210134
rect -8076 174454 -7456 209898
rect -8076 174218 -8044 174454
rect -7808 174218 -7724 174454
rect -7488 174218 -7456 174454
rect -8076 174134 -7456 174218
rect -8076 173898 -8044 174134
rect -7808 173898 -7724 174134
rect -7488 173898 -7456 174134
rect -8076 138454 -7456 173898
rect -8076 138218 -8044 138454
rect -7808 138218 -7724 138454
rect -7488 138218 -7456 138454
rect -8076 138134 -7456 138218
rect -8076 137898 -8044 138134
rect -7808 137898 -7724 138134
rect -7488 137898 -7456 138134
rect -8076 102454 -7456 137898
rect -8076 102218 -8044 102454
rect -7808 102218 -7724 102454
rect -7488 102218 -7456 102454
rect -8076 102134 -7456 102218
rect -8076 101898 -8044 102134
rect -7808 101898 -7724 102134
rect -7488 101898 -7456 102134
rect -8076 66454 -7456 101898
rect -8076 66218 -8044 66454
rect -7808 66218 -7724 66454
rect -7488 66218 -7456 66454
rect -8076 66134 -7456 66218
rect -8076 65898 -8044 66134
rect -7808 65898 -7724 66134
rect -7488 65898 -7456 66134
rect -8076 30454 -7456 65898
rect -8076 30218 -8044 30454
rect -7808 30218 -7724 30454
rect -7488 30218 -7456 30454
rect -8076 30134 -7456 30218
rect -8076 29898 -8044 30134
rect -7808 29898 -7724 30134
rect -7488 29898 -7456 30134
rect -8076 -6416 -7456 29898
rect -7116 709948 -6496 709980
rect -7116 709712 -7084 709948
rect -6848 709712 -6764 709948
rect -6528 709712 -6496 709948
rect -7116 709628 -6496 709712
rect -7116 709392 -7084 709628
rect -6848 709392 -6764 709628
rect -6528 709392 -6496 709628
rect -7116 673954 -6496 709392
rect -7116 673718 -7084 673954
rect -6848 673718 -6764 673954
rect -6528 673718 -6496 673954
rect -7116 673634 -6496 673718
rect -7116 673398 -7084 673634
rect -6848 673398 -6764 673634
rect -6528 673398 -6496 673634
rect -7116 637954 -6496 673398
rect -7116 637718 -7084 637954
rect -6848 637718 -6764 637954
rect -6528 637718 -6496 637954
rect -7116 637634 -6496 637718
rect -7116 637398 -7084 637634
rect -6848 637398 -6764 637634
rect -6528 637398 -6496 637634
rect -7116 601954 -6496 637398
rect -7116 601718 -7084 601954
rect -6848 601718 -6764 601954
rect -6528 601718 -6496 601954
rect -7116 601634 -6496 601718
rect -7116 601398 -7084 601634
rect -6848 601398 -6764 601634
rect -6528 601398 -6496 601634
rect -7116 565954 -6496 601398
rect -7116 565718 -7084 565954
rect -6848 565718 -6764 565954
rect -6528 565718 -6496 565954
rect -7116 565634 -6496 565718
rect -7116 565398 -7084 565634
rect -6848 565398 -6764 565634
rect -6528 565398 -6496 565634
rect -7116 529954 -6496 565398
rect -7116 529718 -7084 529954
rect -6848 529718 -6764 529954
rect -6528 529718 -6496 529954
rect -7116 529634 -6496 529718
rect -7116 529398 -7084 529634
rect -6848 529398 -6764 529634
rect -6528 529398 -6496 529634
rect -7116 493954 -6496 529398
rect -7116 493718 -7084 493954
rect -6848 493718 -6764 493954
rect -6528 493718 -6496 493954
rect -7116 493634 -6496 493718
rect -7116 493398 -7084 493634
rect -6848 493398 -6764 493634
rect -6528 493398 -6496 493634
rect -7116 457954 -6496 493398
rect -7116 457718 -7084 457954
rect -6848 457718 -6764 457954
rect -6528 457718 -6496 457954
rect -7116 457634 -6496 457718
rect -7116 457398 -7084 457634
rect -6848 457398 -6764 457634
rect -6528 457398 -6496 457634
rect -7116 421954 -6496 457398
rect -7116 421718 -7084 421954
rect -6848 421718 -6764 421954
rect -6528 421718 -6496 421954
rect -7116 421634 -6496 421718
rect -7116 421398 -7084 421634
rect -6848 421398 -6764 421634
rect -6528 421398 -6496 421634
rect -7116 385954 -6496 421398
rect -7116 385718 -7084 385954
rect -6848 385718 -6764 385954
rect -6528 385718 -6496 385954
rect -7116 385634 -6496 385718
rect -7116 385398 -7084 385634
rect -6848 385398 -6764 385634
rect -6528 385398 -6496 385634
rect -7116 349954 -6496 385398
rect -7116 349718 -7084 349954
rect -6848 349718 -6764 349954
rect -6528 349718 -6496 349954
rect -7116 349634 -6496 349718
rect -7116 349398 -7084 349634
rect -6848 349398 -6764 349634
rect -6528 349398 -6496 349634
rect -7116 313954 -6496 349398
rect -7116 313718 -7084 313954
rect -6848 313718 -6764 313954
rect -6528 313718 -6496 313954
rect -7116 313634 -6496 313718
rect -7116 313398 -7084 313634
rect -6848 313398 -6764 313634
rect -6528 313398 -6496 313634
rect -7116 277954 -6496 313398
rect -7116 277718 -7084 277954
rect -6848 277718 -6764 277954
rect -6528 277718 -6496 277954
rect -7116 277634 -6496 277718
rect -7116 277398 -7084 277634
rect -6848 277398 -6764 277634
rect -6528 277398 -6496 277634
rect -7116 241954 -6496 277398
rect -7116 241718 -7084 241954
rect -6848 241718 -6764 241954
rect -6528 241718 -6496 241954
rect -7116 241634 -6496 241718
rect -7116 241398 -7084 241634
rect -6848 241398 -6764 241634
rect -6528 241398 -6496 241634
rect -7116 205954 -6496 241398
rect -7116 205718 -7084 205954
rect -6848 205718 -6764 205954
rect -6528 205718 -6496 205954
rect -7116 205634 -6496 205718
rect -7116 205398 -7084 205634
rect -6848 205398 -6764 205634
rect -6528 205398 -6496 205634
rect -7116 169954 -6496 205398
rect -7116 169718 -7084 169954
rect -6848 169718 -6764 169954
rect -6528 169718 -6496 169954
rect -7116 169634 -6496 169718
rect -7116 169398 -7084 169634
rect -6848 169398 -6764 169634
rect -6528 169398 -6496 169634
rect -7116 133954 -6496 169398
rect -7116 133718 -7084 133954
rect -6848 133718 -6764 133954
rect -6528 133718 -6496 133954
rect -7116 133634 -6496 133718
rect -7116 133398 -7084 133634
rect -6848 133398 -6764 133634
rect -6528 133398 -6496 133634
rect -7116 97954 -6496 133398
rect -7116 97718 -7084 97954
rect -6848 97718 -6764 97954
rect -6528 97718 -6496 97954
rect -7116 97634 -6496 97718
rect -7116 97398 -7084 97634
rect -6848 97398 -6764 97634
rect -6528 97398 -6496 97634
rect -7116 61954 -6496 97398
rect -7116 61718 -7084 61954
rect -6848 61718 -6764 61954
rect -6528 61718 -6496 61954
rect -7116 61634 -6496 61718
rect -7116 61398 -7084 61634
rect -6848 61398 -6764 61634
rect -6528 61398 -6496 61634
rect -7116 25954 -6496 61398
rect -7116 25718 -7084 25954
rect -6848 25718 -6764 25954
rect -6528 25718 -6496 25954
rect -7116 25634 -6496 25718
rect -7116 25398 -7084 25634
rect -6848 25398 -6764 25634
rect -6528 25398 -6496 25634
rect -7116 -5456 -6496 25398
rect -6156 708988 -5536 709020
rect -6156 708752 -6124 708988
rect -5888 708752 -5804 708988
rect -5568 708752 -5536 708988
rect -6156 708668 -5536 708752
rect -6156 708432 -6124 708668
rect -5888 708432 -5804 708668
rect -5568 708432 -5536 708668
rect -6156 669454 -5536 708432
rect -6156 669218 -6124 669454
rect -5888 669218 -5804 669454
rect -5568 669218 -5536 669454
rect -6156 669134 -5536 669218
rect -6156 668898 -6124 669134
rect -5888 668898 -5804 669134
rect -5568 668898 -5536 669134
rect -6156 633454 -5536 668898
rect -6156 633218 -6124 633454
rect -5888 633218 -5804 633454
rect -5568 633218 -5536 633454
rect -6156 633134 -5536 633218
rect -6156 632898 -6124 633134
rect -5888 632898 -5804 633134
rect -5568 632898 -5536 633134
rect -6156 597454 -5536 632898
rect -6156 597218 -6124 597454
rect -5888 597218 -5804 597454
rect -5568 597218 -5536 597454
rect -6156 597134 -5536 597218
rect -6156 596898 -6124 597134
rect -5888 596898 -5804 597134
rect -5568 596898 -5536 597134
rect -6156 561454 -5536 596898
rect -6156 561218 -6124 561454
rect -5888 561218 -5804 561454
rect -5568 561218 -5536 561454
rect -6156 561134 -5536 561218
rect -6156 560898 -6124 561134
rect -5888 560898 -5804 561134
rect -5568 560898 -5536 561134
rect -6156 525454 -5536 560898
rect -6156 525218 -6124 525454
rect -5888 525218 -5804 525454
rect -5568 525218 -5536 525454
rect -6156 525134 -5536 525218
rect -6156 524898 -6124 525134
rect -5888 524898 -5804 525134
rect -5568 524898 -5536 525134
rect -6156 489454 -5536 524898
rect -6156 489218 -6124 489454
rect -5888 489218 -5804 489454
rect -5568 489218 -5536 489454
rect -6156 489134 -5536 489218
rect -6156 488898 -6124 489134
rect -5888 488898 -5804 489134
rect -5568 488898 -5536 489134
rect -6156 453454 -5536 488898
rect -6156 453218 -6124 453454
rect -5888 453218 -5804 453454
rect -5568 453218 -5536 453454
rect -6156 453134 -5536 453218
rect -6156 452898 -6124 453134
rect -5888 452898 -5804 453134
rect -5568 452898 -5536 453134
rect -6156 417454 -5536 452898
rect -6156 417218 -6124 417454
rect -5888 417218 -5804 417454
rect -5568 417218 -5536 417454
rect -6156 417134 -5536 417218
rect -6156 416898 -6124 417134
rect -5888 416898 -5804 417134
rect -5568 416898 -5536 417134
rect -6156 381454 -5536 416898
rect -6156 381218 -6124 381454
rect -5888 381218 -5804 381454
rect -5568 381218 -5536 381454
rect -6156 381134 -5536 381218
rect -6156 380898 -6124 381134
rect -5888 380898 -5804 381134
rect -5568 380898 -5536 381134
rect -6156 345454 -5536 380898
rect -6156 345218 -6124 345454
rect -5888 345218 -5804 345454
rect -5568 345218 -5536 345454
rect -6156 345134 -5536 345218
rect -6156 344898 -6124 345134
rect -5888 344898 -5804 345134
rect -5568 344898 -5536 345134
rect -6156 309454 -5536 344898
rect -6156 309218 -6124 309454
rect -5888 309218 -5804 309454
rect -5568 309218 -5536 309454
rect -6156 309134 -5536 309218
rect -6156 308898 -6124 309134
rect -5888 308898 -5804 309134
rect -5568 308898 -5536 309134
rect -6156 273454 -5536 308898
rect -6156 273218 -6124 273454
rect -5888 273218 -5804 273454
rect -5568 273218 -5536 273454
rect -6156 273134 -5536 273218
rect -6156 272898 -6124 273134
rect -5888 272898 -5804 273134
rect -5568 272898 -5536 273134
rect -6156 237454 -5536 272898
rect -6156 237218 -6124 237454
rect -5888 237218 -5804 237454
rect -5568 237218 -5536 237454
rect -6156 237134 -5536 237218
rect -6156 236898 -6124 237134
rect -5888 236898 -5804 237134
rect -5568 236898 -5536 237134
rect -6156 201454 -5536 236898
rect -6156 201218 -6124 201454
rect -5888 201218 -5804 201454
rect -5568 201218 -5536 201454
rect -6156 201134 -5536 201218
rect -6156 200898 -6124 201134
rect -5888 200898 -5804 201134
rect -5568 200898 -5536 201134
rect -6156 165454 -5536 200898
rect -6156 165218 -6124 165454
rect -5888 165218 -5804 165454
rect -5568 165218 -5536 165454
rect -6156 165134 -5536 165218
rect -6156 164898 -6124 165134
rect -5888 164898 -5804 165134
rect -5568 164898 -5536 165134
rect -6156 129454 -5536 164898
rect -6156 129218 -6124 129454
rect -5888 129218 -5804 129454
rect -5568 129218 -5536 129454
rect -6156 129134 -5536 129218
rect -6156 128898 -6124 129134
rect -5888 128898 -5804 129134
rect -5568 128898 -5536 129134
rect -6156 93454 -5536 128898
rect -6156 93218 -6124 93454
rect -5888 93218 -5804 93454
rect -5568 93218 -5536 93454
rect -6156 93134 -5536 93218
rect -6156 92898 -6124 93134
rect -5888 92898 -5804 93134
rect -5568 92898 -5536 93134
rect -6156 57454 -5536 92898
rect -6156 57218 -6124 57454
rect -5888 57218 -5804 57454
rect -5568 57218 -5536 57454
rect -6156 57134 -5536 57218
rect -6156 56898 -6124 57134
rect -5888 56898 -5804 57134
rect -5568 56898 -5536 57134
rect -6156 21454 -5536 56898
rect -6156 21218 -6124 21454
rect -5888 21218 -5804 21454
rect -5568 21218 -5536 21454
rect -6156 21134 -5536 21218
rect -6156 20898 -6124 21134
rect -5888 20898 -5804 21134
rect -5568 20898 -5536 21134
rect -6156 -4496 -5536 20898
rect -5196 708028 -4576 708060
rect -5196 707792 -5164 708028
rect -4928 707792 -4844 708028
rect -4608 707792 -4576 708028
rect -5196 707708 -4576 707792
rect -5196 707472 -5164 707708
rect -4928 707472 -4844 707708
rect -4608 707472 -4576 707708
rect -5196 700954 -4576 707472
rect -5196 700718 -5164 700954
rect -4928 700718 -4844 700954
rect -4608 700718 -4576 700954
rect -5196 700634 -4576 700718
rect -5196 700398 -5164 700634
rect -4928 700398 -4844 700634
rect -4608 700398 -4576 700634
rect -5196 664954 -4576 700398
rect -5196 664718 -5164 664954
rect -4928 664718 -4844 664954
rect -4608 664718 -4576 664954
rect -5196 664634 -4576 664718
rect -5196 664398 -5164 664634
rect -4928 664398 -4844 664634
rect -4608 664398 -4576 664634
rect -5196 628954 -4576 664398
rect -5196 628718 -5164 628954
rect -4928 628718 -4844 628954
rect -4608 628718 -4576 628954
rect -5196 628634 -4576 628718
rect -5196 628398 -5164 628634
rect -4928 628398 -4844 628634
rect -4608 628398 -4576 628634
rect -5196 592954 -4576 628398
rect -5196 592718 -5164 592954
rect -4928 592718 -4844 592954
rect -4608 592718 -4576 592954
rect -5196 592634 -4576 592718
rect -5196 592398 -5164 592634
rect -4928 592398 -4844 592634
rect -4608 592398 -4576 592634
rect -5196 556954 -4576 592398
rect -5196 556718 -5164 556954
rect -4928 556718 -4844 556954
rect -4608 556718 -4576 556954
rect -5196 556634 -4576 556718
rect -5196 556398 -5164 556634
rect -4928 556398 -4844 556634
rect -4608 556398 -4576 556634
rect -5196 520954 -4576 556398
rect -5196 520718 -5164 520954
rect -4928 520718 -4844 520954
rect -4608 520718 -4576 520954
rect -5196 520634 -4576 520718
rect -5196 520398 -5164 520634
rect -4928 520398 -4844 520634
rect -4608 520398 -4576 520634
rect -5196 484954 -4576 520398
rect -5196 484718 -5164 484954
rect -4928 484718 -4844 484954
rect -4608 484718 -4576 484954
rect -5196 484634 -4576 484718
rect -5196 484398 -5164 484634
rect -4928 484398 -4844 484634
rect -4608 484398 -4576 484634
rect -5196 448954 -4576 484398
rect -5196 448718 -5164 448954
rect -4928 448718 -4844 448954
rect -4608 448718 -4576 448954
rect -5196 448634 -4576 448718
rect -5196 448398 -5164 448634
rect -4928 448398 -4844 448634
rect -4608 448398 -4576 448634
rect -5196 412954 -4576 448398
rect -5196 412718 -5164 412954
rect -4928 412718 -4844 412954
rect -4608 412718 -4576 412954
rect -5196 412634 -4576 412718
rect -5196 412398 -5164 412634
rect -4928 412398 -4844 412634
rect -4608 412398 -4576 412634
rect -5196 376954 -4576 412398
rect -5196 376718 -5164 376954
rect -4928 376718 -4844 376954
rect -4608 376718 -4576 376954
rect -5196 376634 -4576 376718
rect -5196 376398 -5164 376634
rect -4928 376398 -4844 376634
rect -4608 376398 -4576 376634
rect -5196 340954 -4576 376398
rect -5196 340718 -5164 340954
rect -4928 340718 -4844 340954
rect -4608 340718 -4576 340954
rect -5196 340634 -4576 340718
rect -5196 340398 -5164 340634
rect -4928 340398 -4844 340634
rect -4608 340398 -4576 340634
rect -5196 304954 -4576 340398
rect -5196 304718 -5164 304954
rect -4928 304718 -4844 304954
rect -4608 304718 -4576 304954
rect -5196 304634 -4576 304718
rect -5196 304398 -5164 304634
rect -4928 304398 -4844 304634
rect -4608 304398 -4576 304634
rect -5196 268954 -4576 304398
rect -5196 268718 -5164 268954
rect -4928 268718 -4844 268954
rect -4608 268718 -4576 268954
rect -5196 268634 -4576 268718
rect -5196 268398 -5164 268634
rect -4928 268398 -4844 268634
rect -4608 268398 -4576 268634
rect -5196 232954 -4576 268398
rect -5196 232718 -5164 232954
rect -4928 232718 -4844 232954
rect -4608 232718 -4576 232954
rect -5196 232634 -4576 232718
rect -5196 232398 -5164 232634
rect -4928 232398 -4844 232634
rect -4608 232398 -4576 232634
rect -5196 196954 -4576 232398
rect -5196 196718 -5164 196954
rect -4928 196718 -4844 196954
rect -4608 196718 -4576 196954
rect -5196 196634 -4576 196718
rect -5196 196398 -5164 196634
rect -4928 196398 -4844 196634
rect -4608 196398 -4576 196634
rect -5196 160954 -4576 196398
rect -5196 160718 -5164 160954
rect -4928 160718 -4844 160954
rect -4608 160718 -4576 160954
rect -5196 160634 -4576 160718
rect -5196 160398 -5164 160634
rect -4928 160398 -4844 160634
rect -4608 160398 -4576 160634
rect -5196 124954 -4576 160398
rect -5196 124718 -5164 124954
rect -4928 124718 -4844 124954
rect -4608 124718 -4576 124954
rect -5196 124634 -4576 124718
rect -5196 124398 -5164 124634
rect -4928 124398 -4844 124634
rect -4608 124398 -4576 124634
rect -5196 88954 -4576 124398
rect -5196 88718 -5164 88954
rect -4928 88718 -4844 88954
rect -4608 88718 -4576 88954
rect -5196 88634 -4576 88718
rect -5196 88398 -5164 88634
rect -4928 88398 -4844 88634
rect -4608 88398 -4576 88634
rect -5196 52954 -4576 88398
rect -5196 52718 -5164 52954
rect -4928 52718 -4844 52954
rect -4608 52718 -4576 52954
rect -5196 52634 -4576 52718
rect -5196 52398 -5164 52634
rect -4928 52398 -4844 52634
rect -4608 52398 -4576 52634
rect -5196 16954 -4576 52398
rect -5196 16718 -5164 16954
rect -4928 16718 -4844 16954
rect -4608 16718 -4576 16954
rect -5196 16634 -4576 16718
rect -5196 16398 -5164 16634
rect -4928 16398 -4844 16634
rect -4608 16398 -4576 16634
rect -5196 -3536 -4576 16398
rect -4236 707068 -3616 707100
rect -4236 706832 -4204 707068
rect -3968 706832 -3884 707068
rect -3648 706832 -3616 707068
rect -4236 706748 -3616 706832
rect -4236 706512 -4204 706748
rect -3968 706512 -3884 706748
rect -3648 706512 -3616 706748
rect -4236 696454 -3616 706512
rect -4236 696218 -4204 696454
rect -3968 696218 -3884 696454
rect -3648 696218 -3616 696454
rect -4236 696134 -3616 696218
rect -4236 695898 -4204 696134
rect -3968 695898 -3884 696134
rect -3648 695898 -3616 696134
rect -4236 660454 -3616 695898
rect -4236 660218 -4204 660454
rect -3968 660218 -3884 660454
rect -3648 660218 -3616 660454
rect -4236 660134 -3616 660218
rect -4236 659898 -4204 660134
rect -3968 659898 -3884 660134
rect -3648 659898 -3616 660134
rect -4236 624454 -3616 659898
rect -4236 624218 -4204 624454
rect -3968 624218 -3884 624454
rect -3648 624218 -3616 624454
rect -4236 624134 -3616 624218
rect -4236 623898 -4204 624134
rect -3968 623898 -3884 624134
rect -3648 623898 -3616 624134
rect -4236 588454 -3616 623898
rect -4236 588218 -4204 588454
rect -3968 588218 -3884 588454
rect -3648 588218 -3616 588454
rect -4236 588134 -3616 588218
rect -4236 587898 -4204 588134
rect -3968 587898 -3884 588134
rect -3648 587898 -3616 588134
rect -4236 552454 -3616 587898
rect -4236 552218 -4204 552454
rect -3968 552218 -3884 552454
rect -3648 552218 -3616 552454
rect -4236 552134 -3616 552218
rect -4236 551898 -4204 552134
rect -3968 551898 -3884 552134
rect -3648 551898 -3616 552134
rect -4236 516454 -3616 551898
rect -4236 516218 -4204 516454
rect -3968 516218 -3884 516454
rect -3648 516218 -3616 516454
rect -4236 516134 -3616 516218
rect -4236 515898 -4204 516134
rect -3968 515898 -3884 516134
rect -3648 515898 -3616 516134
rect -4236 480454 -3616 515898
rect -4236 480218 -4204 480454
rect -3968 480218 -3884 480454
rect -3648 480218 -3616 480454
rect -4236 480134 -3616 480218
rect -4236 479898 -4204 480134
rect -3968 479898 -3884 480134
rect -3648 479898 -3616 480134
rect -4236 444454 -3616 479898
rect -4236 444218 -4204 444454
rect -3968 444218 -3884 444454
rect -3648 444218 -3616 444454
rect -4236 444134 -3616 444218
rect -4236 443898 -4204 444134
rect -3968 443898 -3884 444134
rect -3648 443898 -3616 444134
rect -4236 408454 -3616 443898
rect -4236 408218 -4204 408454
rect -3968 408218 -3884 408454
rect -3648 408218 -3616 408454
rect -4236 408134 -3616 408218
rect -4236 407898 -4204 408134
rect -3968 407898 -3884 408134
rect -3648 407898 -3616 408134
rect -4236 372454 -3616 407898
rect -4236 372218 -4204 372454
rect -3968 372218 -3884 372454
rect -3648 372218 -3616 372454
rect -4236 372134 -3616 372218
rect -4236 371898 -4204 372134
rect -3968 371898 -3884 372134
rect -3648 371898 -3616 372134
rect -4236 336454 -3616 371898
rect -4236 336218 -4204 336454
rect -3968 336218 -3884 336454
rect -3648 336218 -3616 336454
rect -4236 336134 -3616 336218
rect -4236 335898 -4204 336134
rect -3968 335898 -3884 336134
rect -3648 335898 -3616 336134
rect -4236 300454 -3616 335898
rect -4236 300218 -4204 300454
rect -3968 300218 -3884 300454
rect -3648 300218 -3616 300454
rect -4236 300134 -3616 300218
rect -4236 299898 -4204 300134
rect -3968 299898 -3884 300134
rect -3648 299898 -3616 300134
rect -4236 264454 -3616 299898
rect -4236 264218 -4204 264454
rect -3968 264218 -3884 264454
rect -3648 264218 -3616 264454
rect -4236 264134 -3616 264218
rect -4236 263898 -4204 264134
rect -3968 263898 -3884 264134
rect -3648 263898 -3616 264134
rect -4236 228454 -3616 263898
rect -4236 228218 -4204 228454
rect -3968 228218 -3884 228454
rect -3648 228218 -3616 228454
rect -4236 228134 -3616 228218
rect -4236 227898 -4204 228134
rect -3968 227898 -3884 228134
rect -3648 227898 -3616 228134
rect -4236 192454 -3616 227898
rect -4236 192218 -4204 192454
rect -3968 192218 -3884 192454
rect -3648 192218 -3616 192454
rect -4236 192134 -3616 192218
rect -4236 191898 -4204 192134
rect -3968 191898 -3884 192134
rect -3648 191898 -3616 192134
rect -4236 156454 -3616 191898
rect -4236 156218 -4204 156454
rect -3968 156218 -3884 156454
rect -3648 156218 -3616 156454
rect -4236 156134 -3616 156218
rect -4236 155898 -4204 156134
rect -3968 155898 -3884 156134
rect -3648 155898 -3616 156134
rect -4236 120454 -3616 155898
rect -4236 120218 -4204 120454
rect -3968 120218 -3884 120454
rect -3648 120218 -3616 120454
rect -4236 120134 -3616 120218
rect -4236 119898 -4204 120134
rect -3968 119898 -3884 120134
rect -3648 119898 -3616 120134
rect -4236 84454 -3616 119898
rect -4236 84218 -4204 84454
rect -3968 84218 -3884 84454
rect -3648 84218 -3616 84454
rect -4236 84134 -3616 84218
rect -4236 83898 -4204 84134
rect -3968 83898 -3884 84134
rect -3648 83898 -3616 84134
rect -4236 48454 -3616 83898
rect -4236 48218 -4204 48454
rect -3968 48218 -3884 48454
rect -3648 48218 -3616 48454
rect -4236 48134 -3616 48218
rect -4236 47898 -4204 48134
rect -3968 47898 -3884 48134
rect -3648 47898 -3616 48134
rect -4236 12454 -3616 47898
rect -4236 12218 -4204 12454
rect -3968 12218 -3884 12454
rect -3648 12218 -3616 12454
rect -4236 12134 -3616 12218
rect -4236 11898 -4204 12134
rect -3968 11898 -3884 12134
rect -3648 11898 -3616 12134
rect -4236 -2576 -3616 11898
rect -3276 706108 -2656 706140
rect -3276 705872 -3244 706108
rect -3008 705872 -2924 706108
rect -2688 705872 -2656 706108
rect -3276 705788 -2656 705872
rect -3276 705552 -3244 705788
rect -3008 705552 -2924 705788
rect -2688 705552 -2656 705788
rect -3276 691954 -2656 705552
rect -3276 691718 -3244 691954
rect -3008 691718 -2924 691954
rect -2688 691718 -2656 691954
rect -3276 691634 -2656 691718
rect -3276 691398 -3244 691634
rect -3008 691398 -2924 691634
rect -2688 691398 -2656 691634
rect -3276 655954 -2656 691398
rect -3276 655718 -3244 655954
rect -3008 655718 -2924 655954
rect -2688 655718 -2656 655954
rect -3276 655634 -2656 655718
rect -3276 655398 -3244 655634
rect -3008 655398 -2924 655634
rect -2688 655398 -2656 655634
rect -3276 619954 -2656 655398
rect -3276 619718 -3244 619954
rect -3008 619718 -2924 619954
rect -2688 619718 -2656 619954
rect -3276 619634 -2656 619718
rect -3276 619398 -3244 619634
rect -3008 619398 -2924 619634
rect -2688 619398 -2656 619634
rect -3276 583954 -2656 619398
rect -3276 583718 -3244 583954
rect -3008 583718 -2924 583954
rect -2688 583718 -2656 583954
rect -3276 583634 -2656 583718
rect -3276 583398 -3244 583634
rect -3008 583398 -2924 583634
rect -2688 583398 -2656 583634
rect -3276 547954 -2656 583398
rect -3276 547718 -3244 547954
rect -3008 547718 -2924 547954
rect -2688 547718 -2656 547954
rect -3276 547634 -2656 547718
rect -3276 547398 -3244 547634
rect -3008 547398 -2924 547634
rect -2688 547398 -2656 547634
rect -3276 511954 -2656 547398
rect -3276 511718 -3244 511954
rect -3008 511718 -2924 511954
rect -2688 511718 -2656 511954
rect -3276 511634 -2656 511718
rect -3276 511398 -3244 511634
rect -3008 511398 -2924 511634
rect -2688 511398 -2656 511634
rect -3276 475954 -2656 511398
rect -3276 475718 -3244 475954
rect -3008 475718 -2924 475954
rect -2688 475718 -2656 475954
rect -3276 475634 -2656 475718
rect -3276 475398 -3244 475634
rect -3008 475398 -2924 475634
rect -2688 475398 -2656 475634
rect -3276 439954 -2656 475398
rect -3276 439718 -3244 439954
rect -3008 439718 -2924 439954
rect -2688 439718 -2656 439954
rect -3276 439634 -2656 439718
rect -3276 439398 -3244 439634
rect -3008 439398 -2924 439634
rect -2688 439398 -2656 439634
rect -3276 403954 -2656 439398
rect -3276 403718 -3244 403954
rect -3008 403718 -2924 403954
rect -2688 403718 -2656 403954
rect -3276 403634 -2656 403718
rect -3276 403398 -3244 403634
rect -3008 403398 -2924 403634
rect -2688 403398 -2656 403634
rect -3276 367954 -2656 403398
rect -3276 367718 -3244 367954
rect -3008 367718 -2924 367954
rect -2688 367718 -2656 367954
rect -3276 367634 -2656 367718
rect -3276 367398 -3244 367634
rect -3008 367398 -2924 367634
rect -2688 367398 -2656 367634
rect -3276 331954 -2656 367398
rect -3276 331718 -3244 331954
rect -3008 331718 -2924 331954
rect -2688 331718 -2656 331954
rect -3276 331634 -2656 331718
rect -3276 331398 -3244 331634
rect -3008 331398 -2924 331634
rect -2688 331398 -2656 331634
rect -3276 295954 -2656 331398
rect -3276 295718 -3244 295954
rect -3008 295718 -2924 295954
rect -2688 295718 -2656 295954
rect -3276 295634 -2656 295718
rect -3276 295398 -3244 295634
rect -3008 295398 -2924 295634
rect -2688 295398 -2656 295634
rect -3276 259954 -2656 295398
rect -3276 259718 -3244 259954
rect -3008 259718 -2924 259954
rect -2688 259718 -2656 259954
rect -3276 259634 -2656 259718
rect -3276 259398 -3244 259634
rect -3008 259398 -2924 259634
rect -2688 259398 -2656 259634
rect -3276 223954 -2656 259398
rect -3276 223718 -3244 223954
rect -3008 223718 -2924 223954
rect -2688 223718 -2656 223954
rect -3276 223634 -2656 223718
rect -3276 223398 -3244 223634
rect -3008 223398 -2924 223634
rect -2688 223398 -2656 223634
rect -3276 187954 -2656 223398
rect -3276 187718 -3244 187954
rect -3008 187718 -2924 187954
rect -2688 187718 -2656 187954
rect -3276 187634 -2656 187718
rect -3276 187398 -3244 187634
rect -3008 187398 -2924 187634
rect -2688 187398 -2656 187634
rect -3276 151954 -2656 187398
rect -3276 151718 -3244 151954
rect -3008 151718 -2924 151954
rect -2688 151718 -2656 151954
rect -3276 151634 -2656 151718
rect -3276 151398 -3244 151634
rect -3008 151398 -2924 151634
rect -2688 151398 -2656 151634
rect -3276 115954 -2656 151398
rect -3276 115718 -3244 115954
rect -3008 115718 -2924 115954
rect -2688 115718 -2656 115954
rect -3276 115634 -2656 115718
rect -3276 115398 -3244 115634
rect -3008 115398 -2924 115634
rect -2688 115398 -2656 115634
rect -3276 79954 -2656 115398
rect -3276 79718 -3244 79954
rect -3008 79718 -2924 79954
rect -2688 79718 -2656 79954
rect -3276 79634 -2656 79718
rect -3276 79398 -3244 79634
rect -3008 79398 -2924 79634
rect -2688 79398 -2656 79634
rect -3276 43954 -2656 79398
rect -3276 43718 -3244 43954
rect -3008 43718 -2924 43954
rect -2688 43718 -2656 43954
rect -3276 43634 -2656 43718
rect -3276 43398 -3244 43634
rect -3008 43398 -2924 43634
rect -2688 43398 -2656 43634
rect -3276 7954 -2656 43398
rect -3276 7718 -3244 7954
rect -3008 7718 -2924 7954
rect -2688 7718 -2656 7954
rect -3276 7634 -2656 7718
rect -3276 7398 -3244 7634
rect -3008 7398 -2924 7634
rect -2688 7398 -2656 7634
rect -3276 -1616 -2656 7398
rect -2316 705148 -1696 705180
rect -2316 704912 -2284 705148
rect -2048 704912 -1964 705148
rect -1728 704912 -1696 705148
rect -2316 704828 -1696 704912
rect -2316 704592 -2284 704828
rect -2048 704592 -1964 704828
rect -1728 704592 -1696 704828
rect -2316 687454 -1696 704592
rect -2316 687218 -2284 687454
rect -2048 687218 -1964 687454
rect -1728 687218 -1696 687454
rect -2316 687134 -1696 687218
rect -2316 686898 -2284 687134
rect -2048 686898 -1964 687134
rect -1728 686898 -1696 687134
rect -2316 651454 -1696 686898
rect -2316 651218 -2284 651454
rect -2048 651218 -1964 651454
rect -1728 651218 -1696 651454
rect -2316 651134 -1696 651218
rect -2316 650898 -2284 651134
rect -2048 650898 -1964 651134
rect -1728 650898 -1696 651134
rect -2316 615454 -1696 650898
rect -2316 615218 -2284 615454
rect -2048 615218 -1964 615454
rect -1728 615218 -1696 615454
rect -2316 615134 -1696 615218
rect -2316 614898 -2284 615134
rect -2048 614898 -1964 615134
rect -1728 614898 -1696 615134
rect -2316 579454 -1696 614898
rect -2316 579218 -2284 579454
rect -2048 579218 -1964 579454
rect -1728 579218 -1696 579454
rect -2316 579134 -1696 579218
rect -2316 578898 -2284 579134
rect -2048 578898 -1964 579134
rect -1728 578898 -1696 579134
rect -2316 543454 -1696 578898
rect -2316 543218 -2284 543454
rect -2048 543218 -1964 543454
rect -1728 543218 -1696 543454
rect -2316 543134 -1696 543218
rect -2316 542898 -2284 543134
rect -2048 542898 -1964 543134
rect -1728 542898 -1696 543134
rect -2316 507454 -1696 542898
rect -2316 507218 -2284 507454
rect -2048 507218 -1964 507454
rect -1728 507218 -1696 507454
rect -2316 507134 -1696 507218
rect -2316 506898 -2284 507134
rect -2048 506898 -1964 507134
rect -1728 506898 -1696 507134
rect -2316 471454 -1696 506898
rect -2316 471218 -2284 471454
rect -2048 471218 -1964 471454
rect -1728 471218 -1696 471454
rect -2316 471134 -1696 471218
rect -2316 470898 -2284 471134
rect -2048 470898 -1964 471134
rect -1728 470898 -1696 471134
rect -2316 435454 -1696 470898
rect -2316 435218 -2284 435454
rect -2048 435218 -1964 435454
rect -1728 435218 -1696 435454
rect -2316 435134 -1696 435218
rect -2316 434898 -2284 435134
rect -2048 434898 -1964 435134
rect -1728 434898 -1696 435134
rect -2316 399454 -1696 434898
rect -2316 399218 -2284 399454
rect -2048 399218 -1964 399454
rect -1728 399218 -1696 399454
rect -2316 399134 -1696 399218
rect -2316 398898 -2284 399134
rect -2048 398898 -1964 399134
rect -1728 398898 -1696 399134
rect -2316 363454 -1696 398898
rect -2316 363218 -2284 363454
rect -2048 363218 -1964 363454
rect -1728 363218 -1696 363454
rect -2316 363134 -1696 363218
rect -2316 362898 -2284 363134
rect -2048 362898 -1964 363134
rect -1728 362898 -1696 363134
rect -2316 327454 -1696 362898
rect -2316 327218 -2284 327454
rect -2048 327218 -1964 327454
rect -1728 327218 -1696 327454
rect -2316 327134 -1696 327218
rect -2316 326898 -2284 327134
rect -2048 326898 -1964 327134
rect -1728 326898 -1696 327134
rect -2316 291454 -1696 326898
rect -2316 291218 -2284 291454
rect -2048 291218 -1964 291454
rect -1728 291218 -1696 291454
rect -2316 291134 -1696 291218
rect -2316 290898 -2284 291134
rect -2048 290898 -1964 291134
rect -1728 290898 -1696 291134
rect -2316 255454 -1696 290898
rect -2316 255218 -2284 255454
rect -2048 255218 -1964 255454
rect -1728 255218 -1696 255454
rect -2316 255134 -1696 255218
rect -2316 254898 -2284 255134
rect -2048 254898 -1964 255134
rect -1728 254898 -1696 255134
rect -2316 219454 -1696 254898
rect -2316 219218 -2284 219454
rect -2048 219218 -1964 219454
rect -1728 219218 -1696 219454
rect -2316 219134 -1696 219218
rect -2316 218898 -2284 219134
rect -2048 218898 -1964 219134
rect -1728 218898 -1696 219134
rect -2316 183454 -1696 218898
rect -2316 183218 -2284 183454
rect -2048 183218 -1964 183454
rect -1728 183218 -1696 183454
rect -2316 183134 -1696 183218
rect -2316 182898 -2284 183134
rect -2048 182898 -1964 183134
rect -1728 182898 -1696 183134
rect -2316 147454 -1696 182898
rect -2316 147218 -2284 147454
rect -2048 147218 -1964 147454
rect -1728 147218 -1696 147454
rect -2316 147134 -1696 147218
rect -2316 146898 -2284 147134
rect -2048 146898 -1964 147134
rect -1728 146898 -1696 147134
rect -2316 111454 -1696 146898
rect -2316 111218 -2284 111454
rect -2048 111218 -1964 111454
rect -1728 111218 -1696 111454
rect -2316 111134 -1696 111218
rect -2316 110898 -2284 111134
rect -2048 110898 -1964 111134
rect -1728 110898 -1696 111134
rect -2316 75454 -1696 110898
rect -2316 75218 -2284 75454
rect -2048 75218 -1964 75454
rect -1728 75218 -1696 75454
rect -2316 75134 -1696 75218
rect -2316 74898 -2284 75134
rect -2048 74898 -1964 75134
rect -1728 74898 -1696 75134
rect -2316 39454 -1696 74898
rect -2316 39218 -2284 39454
rect -2048 39218 -1964 39454
rect -1728 39218 -1696 39454
rect -2316 39134 -1696 39218
rect -2316 38898 -2284 39134
rect -2048 38898 -1964 39134
rect -1728 38898 -1696 39134
rect -2316 3454 -1696 38898
rect -2316 3218 -2284 3454
rect -2048 3218 -1964 3454
rect -1728 3218 -1696 3454
rect -2316 3134 -1696 3218
rect -2316 2898 -2284 3134
rect -2048 2898 -1964 3134
rect -1728 2898 -1696 3134
rect -2316 -656 -1696 2898
rect -2316 -892 -2284 -656
rect -2048 -892 -1964 -656
rect -1728 -892 -1696 -656
rect -2316 -976 -1696 -892
rect -2316 -1212 -2284 -976
rect -2048 -1212 -1964 -976
rect -1728 -1212 -1696 -976
rect -2316 -1244 -1696 -1212
rect 1794 705148 2414 711900
rect 1794 704912 1826 705148
rect 2062 704912 2146 705148
rect 2382 704912 2414 705148
rect 1794 704828 2414 704912
rect 1794 704592 1826 704828
rect 2062 704592 2146 704828
rect 2382 704592 2414 704828
rect 1794 687454 2414 704592
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -656 2414 2898
rect 1794 -892 1826 -656
rect 2062 -892 2146 -656
rect 2382 -892 2414 -656
rect 1794 -976 2414 -892
rect 1794 -1212 1826 -976
rect 2062 -1212 2146 -976
rect 2382 -1212 2414 -976
rect -3276 -1852 -3244 -1616
rect -3008 -1852 -2924 -1616
rect -2688 -1852 -2656 -1616
rect -3276 -1936 -2656 -1852
rect -3276 -2172 -3244 -1936
rect -3008 -2172 -2924 -1936
rect -2688 -2172 -2656 -1936
rect -3276 -2204 -2656 -2172
rect -4236 -2812 -4204 -2576
rect -3968 -2812 -3884 -2576
rect -3648 -2812 -3616 -2576
rect -4236 -2896 -3616 -2812
rect -4236 -3132 -4204 -2896
rect -3968 -3132 -3884 -2896
rect -3648 -3132 -3616 -2896
rect -4236 -3164 -3616 -3132
rect -5196 -3772 -5164 -3536
rect -4928 -3772 -4844 -3536
rect -4608 -3772 -4576 -3536
rect -5196 -3856 -4576 -3772
rect -5196 -4092 -5164 -3856
rect -4928 -4092 -4844 -3856
rect -4608 -4092 -4576 -3856
rect -5196 -4124 -4576 -4092
rect -6156 -4732 -6124 -4496
rect -5888 -4732 -5804 -4496
rect -5568 -4732 -5536 -4496
rect -6156 -4816 -5536 -4732
rect -6156 -5052 -6124 -4816
rect -5888 -5052 -5804 -4816
rect -5568 -5052 -5536 -4816
rect -6156 -5084 -5536 -5052
rect -7116 -5692 -7084 -5456
rect -6848 -5692 -6764 -5456
rect -6528 -5692 -6496 -5456
rect -7116 -5776 -6496 -5692
rect -7116 -6012 -7084 -5776
rect -6848 -6012 -6764 -5776
rect -6528 -6012 -6496 -5776
rect -7116 -6044 -6496 -6012
rect -8076 -6652 -8044 -6416
rect -7808 -6652 -7724 -6416
rect -7488 -6652 -7456 -6416
rect -8076 -6736 -7456 -6652
rect -8076 -6972 -8044 -6736
rect -7808 -6972 -7724 -6736
rect -7488 -6972 -7456 -6736
rect -8076 -7004 -7456 -6972
rect -9036 -7612 -9004 -7376
rect -8768 -7612 -8684 -7376
rect -8448 -7612 -8416 -7376
rect -9036 -7696 -8416 -7612
rect -9036 -7932 -9004 -7696
rect -8768 -7932 -8684 -7696
rect -8448 -7932 -8416 -7696
rect -9036 -7964 -8416 -7932
rect 1794 -7964 2414 -1212
rect 6294 706108 6914 711900
rect 6294 705872 6326 706108
rect 6562 705872 6646 706108
rect 6882 705872 6914 706108
rect 6294 705788 6914 705872
rect 6294 705552 6326 705788
rect 6562 705552 6646 705788
rect 6882 705552 6914 705788
rect 6294 691954 6914 705552
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1616 6914 7398
rect 6294 -1852 6326 -1616
rect 6562 -1852 6646 -1616
rect 6882 -1852 6914 -1616
rect 6294 -1936 6914 -1852
rect 6294 -2172 6326 -1936
rect 6562 -2172 6646 -1936
rect 6882 -2172 6914 -1936
rect 6294 -7964 6914 -2172
rect 10794 707068 11414 711900
rect 10794 706832 10826 707068
rect 11062 706832 11146 707068
rect 11382 706832 11414 707068
rect 10794 706748 11414 706832
rect 10794 706512 10826 706748
rect 11062 706512 11146 706748
rect 11382 706512 11414 706748
rect 10794 696454 11414 706512
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2576 11414 11898
rect 10794 -2812 10826 -2576
rect 11062 -2812 11146 -2576
rect 11382 -2812 11414 -2576
rect 10794 -2896 11414 -2812
rect 10794 -3132 10826 -2896
rect 11062 -3132 11146 -2896
rect 11382 -3132 11414 -2896
rect 10794 -7964 11414 -3132
rect 15294 708028 15914 711900
rect 15294 707792 15326 708028
rect 15562 707792 15646 708028
rect 15882 707792 15914 708028
rect 15294 707708 15914 707792
rect 15294 707472 15326 707708
rect 15562 707472 15646 707708
rect 15882 707472 15914 707708
rect 15294 700954 15914 707472
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3536 15914 16398
rect 15294 -3772 15326 -3536
rect 15562 -3772 15646 -3536
rect 15882 -3772 15914 -3536
rect 15294 -3856 15914 -3772
rect 15294 -4092 15326 -3856
rect 15562 -4092 15646 -3856
rect 15882 -4092 15914 -3856
rect 15294 -7964 15914 -4092
rect 19794 708988 20414 711900
rect 19794 708752 19826 708988
rect 20062 708752 20146 708988
rect 20382 708752 20414 708988
rect 19794 708668 20414 708752
rect 19794 708432 19826 708668
rect 20062 708432 20146 708668
rect 20382 708432 20414 708668
rect 19794 669454 20414 708432
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4496 20414 20898
rect 19794 -4732 19826 -4496
rect 20062 -4732 20146 -4496
rect 20382 -4732 20414 -4496
rect 19794 -4816 20414 -4732
rect 19794 -5052 19826 -4816
rect 20062 -5052 20146 -4816
rect 20382 -5052 20414 -4816
rect 19794 -7964 20414 -5052
rect 24294 709948 24914 711900
rect 24294 709712 24326 709948
rect 24562 709712 24646 709948
rect 24882 709712 24914 709948
rect 24294 709628 24914 709712
rect 24294 709392 24326 709628
rect 24562 709392 24646 709628
rect 24882 709392 24914 709628
rect 24294 673954 24914 709392
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5456 24914 25398
rect 24294 -5692 24326 -5456
rect 24562 -5692 24646 -5456
rect 24882 -5692 24914 -5456
rect 24294 -5776 24914 -5692
rect 24294 -6012 24326 -5776
rect 24562 -6012 24646 -5776
rect 24882 -6012 24914 -5776
rect 24294 -7964 24914 -6012
rect 28794 710908 29414 711900
rect 28794 710672 28826 710908
rect 29062 710672 29146 710908
rect 29382 710672 29414 710908
rect 28794 710588 29414 710672
rect 28794 710352 28826 710588
rect 29062 710352 29146 710588
rect 29382 710352 29414 710588
rect 28794 678454 29414 710352
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6416 29414 29898
rect 28794 -6652 28826 -6416
rect 29062 -6652 29146 -6416
rect 29382 -6652 29414 -6416
rect 28794 -6736 29414 -6652
rect 28794 -6972 28826 -6736
rect 29062 -6972 29146 -6736
rect 29382 -6972 29414 -6736
rect 28794 -7964 29414 -6972
rect 33294 711868 33914 711900
rect 33294 711632 33326 711868
rect 33562 711632 33646 711868
rect 33882 711632 33914 711868
rect 33294 711548 33914 711632
rect 33294 711312 33326 711548
rect 33562 711312 33646 711548
rect 33882 711312 33914 711548
rect 33294 682954 33914 711312
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7376 33914 34398
rect 33294 -7612 33326 -7376
rect 33562 -7612 33646 -7376
rect 33882 -7612 33914 -7376
rect 33294 -7696 33914 -7612
rect 33294 -7932 33326 -7696
rect 33562 -7932 33646 -7696
rect 33882 -7932 33914 -7696
rect 33294 -7964 33914 -7932
rect 37794 705148 38414 711900
rect 37794 704912 37826 705148
rect 38062 704912 38146 705148
rect 38382 704912 38414 705148
rect 37794 704828 38414 704912
rect 37794 704592 37826 704828
rect 38062 704592 38146 704828
rect 38382 704592 38414 704828
rect 37794 687454 38414 704592
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -656 38414 2898
rect 37794 -892 37826 -656
rect 38062 -892 38146 -656
rect 38382 -892 38414 -656
rect 37794 -976 38414 -892
rect 37794 -1212 37826 -976
rect 38062 -1212 38146 -976
rect 38382 -1212 38414 -976
rect 37794 -7964 38414 -1212
rect 42294 706108 42914 711900
rect 42294 705872 42326 706108
rect 42562 705872 42646 706108
rect 42882 705872 42914 706108
rect 42294 705788 42914 705872
rect 42294 705552 42326 705788
rect 42562 705552 42646 705788
rect 42882 705552 42914 705788
rect 42294 691954 42914 705552
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1616 42914 7398
rect 42294 -1852 42326 -1616
rect 42562 -1852 42646 -1616
rect 42882 -1852 42914 -1616
rect 42294 -1936 42914 -1852
rect 42294 -2172 42326 -1936
rect 42562 -2172 42646 -1936
rect 42882 -2172 42914 -1936
rect 42294 -7964 42914 -2172
rect 46794 707068 47414 711900
rect 46794 706832 46826 707068
rect 47062 706832 47146 707068
rect 47382 706832 47414 707068
rect 46794 706748 47414 706832
rect 46794 706512 46826 706748
rect 47062 706512 47146 706748
rect 47382 706512 47414 706748
rect 46794 696454 47414 706512
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2576 47414 11898
rect 46794 -2812 46826 -2576
rect 47062 -2812 47146 -2576
rect 47382 -2812 47414 -2576
rect 46794 -2896 47414 -2812
rect 46794 -3132 46826 -2896
rect 47062 -3132 47146 -2896
rect 47382 -3132 47414 -2896
rect 46794 -7964 47414 -3132
rect 51294 708028 51914 711900
rect 51294 707792 51326 708028
rect 51562 707792 51646 708028
rect 51882 707792 51914 708028
rect 51294 707708 51914 707792
rect 51294 707472 51326 707708
rect 51562 707472 51646 707708
rect 51882 707472 51914 707708
rect 51294 700954 51914 707472
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3536 51914 16398
rect 51294 -3772 51326 -3536
rect 51562 -3772 51646 -3536
rect 51882 -3772 51914 -3536
rect 51294 -3856 51914 -3772
rect 51294 -4092 51326 -3856
rect 51562 -4092 51646 -3856
rect 51882 -4092 51914 -3856
rect 51294 -7964 51914 -4092
rect 55794 708988 56414 711900
rect 55794 708752 55826 708988
rect 56062 708752 56146 708988
rect 56382 708752 56414 708988
rect 55794 708668 56414 708752
rect 55794 708432 55826 708668
rect 56062 708432 56146 708668
rect 56382 708432 56414 708668
rect 55794 669454 56414 708432
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4496 56414 20898
rect 55794 -4732 55826 -4496
rect 56062 -4732 56146 -4496
rect 56382 -4732 56414 -4496
rect 55794 -4816 56414 -4732
rect 55794 -5052 55826 -4816
rect 56062 -5052 56146 -4816
rect 56382 -5052 56414 -4816
rect 55794 -7964 56414 -5052
rect 60294 709948 60914 711900
rect 60294 709712 60326 709948
rect 60562 709712 60646 709948
rect 60882 709712 60914 709948
rect 60294 709628 60914 709712
rect 60294 709392 60326 709628
rect 60562 709392 60646 709628
rect 60882 709392 60914 709628
rect 60294 673954 60914 709392
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 60294 205954 60914 241398
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5456 60914 25398
rect 60294 -5692 60326 -5456
rect 60562 -5692 60646 -5456
rect 60882 -5692 60914 -5456
rect 60294 -5776 60914 -5692
rect 60294 -6012 60326 -5776
rect 60562 -6012 60646 -5776
rect 60882 -6012 60914 -5776
rect 60294 -7964 60914 -6012
rect 64794 710908 65414 711900
rect 64794 710672 64826 710908
rect 65062 710672 65146 710908
rect 65382 710672 65414 710908
rect 64794 710588 65414 710672
rect 64794 710352 64826 710588
rect 65062 710352 65146 710588
rect 65382 710352 65414 710588
rect 64794 678454 65414 710352
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6416 65414 29898
rect 64794 -6652 64826 -6416
rect 65062 -6652 65146 -6416
rect 65382 -6652 65414 -6416
rect 64794 -6736 65414 -6652
rect 64794 -6972 64826 -6736
rect 65062 -6972 65146 -6736
rect 65382 -6972 65414 -6736
rect 64794 -7964 65414 -6972
rect 69294 711868 69914 711900
rect 69294 711632 69326 711868
rect 69562 711632 69646 711868
rect 69882 711632 69914 711868
rect 69294 711548 69914 711632
rect 69294 711312 69326 711548
rect 69562 711312 69646 711548
rect 69882 711312 69914 711548
rect 69294 682954 69914 711312
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 214954 69914 250398
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7376 69914 34398
rect 69294 -7612 69326 -7376
rect 69562 -7612 69646 -7376
rect 69882 -7612 69914 -7376
rect 69294 -7696 69914 -7612
rect 69294 -7932 69326 -7696
rect 69562 -7932 69646 -7696
rect 69882 -7932 69914 -7696
rect 69294 -7964 69914 -7932
rect 73794 705148 74414 711900
rect 73794 704912 73826 705148
rect 74062 704912 74146 705148
rect 74382 704912 74414 705148
rect 73794 704828 74414 704912
rect 73794 704592 73826 704828
rect 74062 704592 74146 704828
rect 74382 704592 74414 704828
rect 73794 687454 74414 704592
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -656 74414 2898
rect 73794 -892 73826 -656
rect 74062 -892 74146 -656
rect 74382 -892 74414 -656
rect 73794 -976 74414 -892
rect 73794 -1212 73826 -976
rect 74062 -1212 74146 -976
rect 74382 -1212 74414 -976
rect 73794 -7964 74414 -1212
rect 78294 706108 78914 711900
rect 78294 705872 78326 706108
rect 78562 705872 78646 706108
rect 78882 705872 78914 706108
rect 78294 705788 78914 705872
rect 78294 705552 78326 705788
rect 78562 705552 78646 705788
rect 78882 705552 78914 705788
rect 78294 691954 78914 705552
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 223954 78914 259398
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1616 78914 7398
rect 78294 -1852 78326 -1616
rect 78562 -1852 78646 -1616
rect 78882 -1852 78914 -1616
rect 78294 -1936 78914 -1852
rect 78294 -2172 78326 -1936
rect 78562 -2172 78646 -1936
rect 78882 -2172 78914 -1936
rect 78294 -7964 78914 -2172
rect 82794 707068 83414 711900
rect 82794 706832 82826 707068
rect 83062 706832 83146 707068
rect 83382 706832 83414 707068
rect 82794 706748 83414 706832
rect 82794 706512 82826 706748
rect 83062 706512 83146 706748
rect 83382 706512 83414 706748
rect 82794 696454 83414 706512
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 228454 83414 263898
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2576 83414 11898
rect 82794 -2812 82826 -2576
rect 83062 -2812 83146 -2576
rect 83382 -2812 83414 -2576
rect 82794 -2896 83414 -2812
rect 82794 -3132 82826 -2896
rect 83062 -3132 83146 -2896
rect 83382 -3132 83414 -2896
rect 82794 -7964 83414 -3132
rect 87294 708028 87914 711900
rect 87294 707792 87326 708028
rect 87562 707792 87646 708028
rect 87882 707792 87914 708028
rect 87294 707708 87914 707792
rect 87294 707472 87326 707708
rect 87562 707472 87646 707708
rect 87882 707472 87914 707708
rect 87294 700954 87914 707472
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 232954 87914 268398
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3536 87914 16398
rect 87294 -3772 87326 -3536
rect 87562 -3772 87646 -3536
rect 87882 -3772 87914 -3536
rect 87294 -3856 87914 -3772
rect 87294 -4092 87326 -3856
rect 87562 -4092 87646 -3856
rect 87882 -4092 87914 -3856
rect 87294 -7964 87914 -4092
rect 91794 708988 92414 711900
rect 91794 708752 91826 708988
rect 92062 708752 92146 708988
rect 92382 708752 92414 708988
rect 91794 708668 92414 708752
rect 91794 708432 91826 708668
rect 92062 708432 92146 708668
rect 92382 708432 92414 708668
rect 91794 669454 92414 708432
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4496 92414 20898
rect 91794 -4732 91826 -4496
rect 92062 -4732 92146 -4496
rect 92382 -4732 92414 -4496
rect 91794 -4816 92414 -4732
rect 91794 -5052 91826 -4816
rect 92062 -5052 92146 -4816
rect 92382 -5052 92414 -4816
rect 91794 -7964 92414 -5052
rect 96294 709948 96914 711900
rect 96294 709712 96326 709948
rect 96562 709712 96646 709948
rect 96882 709712 96914 709948
rect 96294 709628 96914 709712
rect 96294 709392 96326 709628
rect 96562 709392 96646 709628
rect 96882 709392 96914 709628
rect 96294 673954 96914 709392
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 100794 710908 101414 711900
rect 100794 710672 100826 710908
rect 101062 710672 101146 710908
rect 101382 710672 101414 710908
rect 100794 710588 101414 710672
rect 100794 710352 100826 710588
rect 101062 710352 101146 710588
rect 101382 710352 101414 710588
rect 100794 678454 101414 710352
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 374164 101414 389898
rect 105294 711868 105914 711900
rect 105294 711632 105326 711868
rect 105562 711632 105646 711868
rect 105882 711632 105914 711868
rect 105294 711548 105914 711632
rect 105294 711312 105326 711548
rect 105562 711312 105646 711548
rect 105882 711312 105914 711548
rect 105294 682954 105914 711312
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 374164 105914 394398
rect 109794 705148 110414 711900
rect 109794 704912 109826 705148
rect 110062 704912 110146 705148
rect 110382 704912 110414 705148
rect 109794 704828 110414 704912
rect 109794 704592 109826 704828
rect 110062 704592 110146 704828
rect 110382 704592 110414 704828
rect 109794 687454 110414 704592
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 374164 110414 398898
rect 114294 706108 114914 711900
rect 114294 705872 114326 706108
rect 114562 705872 114646 706108
rect 114882 705872 114914 706108
rect 114294 705788 114914 705872
rect 114294 705552 114326 705788
rect 114562 705552 114646 705788
rect 114882 705552 114914 705788
rect 114294 691954 114914 705552
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 374164 114914 403398
rect 118794 707068 119414 711900
rect 118794 706832 118826 707068
rect 119062 706832 119146 707068
rect 119382 706832 119414 707068
rect 118794 706748 119414 706832
rect 118794 706512 118826 706748
rect 119062 706512 119146 706748
rect 119382 706512 119414 706748
rect 118794 696454 119414 706512
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 374164 119414 407898
rect 123294 708028 123914 711900
rect 123294 707792 123326 708028
rect 123562 707792 123646 708028
rect 123882 707792 123914 708028
rect 123294 707708 123914 707792
rect 123294 707472 123326 707708
rect 123562 707472 123646 707708
rect 123882 707472 123914 707708
rect 123294 700954 123914 707472
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 374164 123914 376398
rect 127794 708988 128414 711900
rect 127794 708752 127826 708988
rect 128062 708752 128146 708988
rect 128382 708752 128414 708988
rect 127794 708668 128414 708752
rect 127794 708432 127826 708668
rect 128062 708432 128146 708668
rect 128382 708432 128414 708668
rect 127794 669454 128414 708432
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 374164 128414 380898
rect 132294 709948 132914 711900
rect 132294 709712 132326 709948
rect 132562 709712 132646 709948
rect 132882 709712 132914 709948
rect 132294 709628 132914 709712
rect 132294 709392 132326 709628
rect 132562 709392 132646 709628
rect 132882 709392 132914 709628
rect 132294 673954 132914 709392
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 374164 132914 385398
rect 136794 710908 137414 711900
rect 136794 710672 136826 710908
rect 137062 710672 137146 710908
rect 137382 710672 137414 710908
rect 136794 710588 137414 710672
rect 136794 710352 136826 710588
rect 137062 710352 137146 710588
rect 137382 710352 137414 710588
rect 136794 678454 137414 710352
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 374164 137414 389898
rect 141294 711868 141914 711900
rect 141294 711632 141326 711868
rect 141562 711632 141646 711868
rect 141882 711632 141914 711868
rect 141294 711548 141914 711632
rect 141294 711312 141326 711548
rect 141562 711312 141646 711548
rect 141882 711312 141914 711548
rect 141294 682954 141914 711312
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 374164 141914 394398
rect 145794 705148 146414 711900
rect 145794 704912 145826 705148
rect 146062 704912 146146 705148
rect 146382 704912 146414 705148
rect 145794 704828 146414 704912
rect 145794 704592 145826 704828
rect 146062 704592 146146 704828
rect 146382 704592 146414 704828
rect 145794 687454 146414 704592
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 374164 146414 398898
rect 150294 706108 150914 711900
rect 150294 705872 150326 706108
rect 150562 705872 150646 706108
rect 150882 705872 150914 706108
rect 150294 705788 150914 705872
rect 150294 705552 150326 705788
rect 150562 705552 150646 705788
rect 150882 705552 150914 705788
rect 150294 691954 150914 705552
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 374164 150914 403398
rect 154794 707068 155414 711900
rect 154794 706832 154826 707068
rect 155062 706832 155146 707068
rect 155382 706832 155414 707068
rect 154794 706748 155414 706832
rect 154794 706512 154826 706748
rect 155062 706512 155146 706748
rect 155382 706512 155414 706748
rect 154794 696454 155414 706512
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 374164 155414 407898
rect 159294 708028 159914 711900
rect 159294 707792 159326 708028
rect 159562 707792 159646 708028
rect 159882 707792 159914 708028
rect 159294 707708 159914 707792
rect 159294 707472 159326 707708
rect 159562 707472 159646 707708
rect 159882 707472 159914 707708
rect 159294 700954 159914 707472
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 374164 159914 376398
rect 163794 708988 164414 711900
rect 163794 708752 163826 708988
rect 164062 708752 164146 708988
rect 164382 708752 164414 708988
rect 163794 708668 164414 708752
rect 163794 708432 163826 708668
rect 164062 708432 164146 708668
rect 164382 708432 164414 708668
rect 163794 669454 164414 708432
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 374164 164414 380898
rect 168294 709948 168914 711900
rect 168294 709712 168326 709948
rect 168562 709712 168646 709948
rect 168882 709712 168914 709948
rect 168294 709628 168914 709712
rect 168294 709392 168326 709628
rect 168562 709392 168646 709628
rect 168882 709392 168914 709628
rect 168294 673954 168914 709392
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 374164 168914 385398
rect 172794 710908 173414 711900
rect 172794 710672 172826 710908
rect 173062 710672 173146 710908
rect 173382 710672 173414 710908
rect 172794 710588 173414 710672
rect 172794 710352 172826 710588
rect 173062 710352 173146 710588
rect 173382 710352 173414 710588
rect 172794 678454 173414 710352
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 119568 367954 119888 367986
rect 119568 367718 119610 367954
rect 119846 367718 119888 367954
rect 119568 367634 119888 367718
rect 119568 367398 119610 367634
rect 119846 367398 119888 367634
rect 119568 367366 119888 367398
rect 150288 367954 150608 367986
rect 150288 367718 150330 367954
rect 150566 367718 150608 367954
rect 150288 367634 150608 367718
rect 150288 367398 150330 367634
rect 150566 367398 150608 367634
rect 150288 367366 150608 367398
rect 104208 363454 104528 363486
rect 104208 363218 104250 363454
rect 104486 363218 104528 363454
rect 104208 363134 104528 363218
rect 104208 362898 104250 363134
rect 104486 362898 104528 363134
rect 104208 362866 104528 362898
rect 134928 363454 135248 363486
rect 134928 363218 134970 363454
rect 135206 363218 135248 363454
rect 134928 363134 135248 363218
rect 134928 362898 134970 363134
rect 135206 362898 135248 363134
rect 134928 362866 135248 362898
rect 165648 363454 165968 363486
rect 165648 363218 165690 363454
rect 165926 363218 165968 363454
rect 165648 363134 165968 363218
rect 165648 362898 165690 363134
rect 165926 362898 165968 363134
rect 165648 362866 165968 362898
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 119568 331954 119888 331986
rect 119568 331718 119610 331954
rect 119846 331718 119888 331954
rect 119568 331634 119888 331718
rect 119568 331398 119610 331634
rect 119846 331398 119888 331634
rect 119568 331366 119888 331398
rect 150288 331954 150608 331986
rect 150288 331718 150330 331954
rect 150566 331718 150608 331954
rect 150288 331634 150608 331718
rect 150288 331398 150330 331634
rect 150566 331398 150608 331634
rect 150288 331366 150608 331398
rect 104208 327454 104528 327486
rect 104208 327218 104250 327454
rect 104486 327218 104528 327454
rect 104208 327134 104528 327218
rect 104208 326898 104250 327134
rect 104486 326898 104528 327134
rect 104208 326866 104528 326898
rect 134928 327454 135248 327486
rect 134928 327218 134970 327454
rect 135206 327218 135248 327454
rect 134928 327134 135248 327218
rect 134928 326898 134970 327134
rect 135206 326898 135248 327134
rect 134928 326866 135248 326898
rect 165648 327454 165968 327486
rect 165648 327218 165690 327454
rect 165926 327218 165968 327454
rect 165648 327134 165968 327218
rect 165648 326898 165690 327134
rect 165926 326898 165968 327134
rect 165648 326866 165968 326898
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 169339 308548 169405 308549
rect 169339 308484 169340 308548
rect 169404 308484 169405 308548
rect 169339 308483 169405 308484
rect 169155 301204 169221 301205
rect 169155 301140 169156 301204
rect 169220 301140 169221 301204
rect 169155 301139 169221 301140
rect 169158 298077 169218 301139
rect 169342 299165 169402 308483
rect 169523 301612 169589 301613
rect 169523 301548 169524 301612
rect 169588 301548 169589 301612
rect 169523 301547 169589 301548
rect 169339 299164 169405 299165
rect 169339 299100 169340 299164
rect 169404 299100 169405 299164
rect 169339 299099 169405 299100
rect 169155 298076 169221 298077
rect 169155 298012 169156 298076
rect 169220 298012 169221 298076
rect 169155 298011 169221 298012
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 241954 96914 277398
rect 96294 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 96914 241954
rect 96294 241634 96914 241718
rect 96294 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 96914 241634
rect 96294 205954 96914 241398
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5456 96914 25398
rect 96294 -5692 96326 -5456
rect 96562 -5692 96646 -5456
rect 96882 -5692 96914 -5456
rect 96294 -5776 96914 -5692
rect 96294 -6012 96326 -5776
rect 96562 -6012 96646 -5776
rect 96882 -6012 96914 -5776
rect 96294 -7964 96914 -6012
rect 100794 282454 101414 298000
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 246454 101414 281898
rect 100794 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 101414 246454
rect 100794 246134 101414 246218
rect 100794 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 101414 246134
rect 100794 210454 101414 245898
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 100794 174454 101414 209898
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 138454 101414 173898
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6416 101414 29898
rect 100794 -6652 100826 -6416
rect 101062 -6652 101146 -6416
rect 101382 -6652 101414 -6416
rect 100794 -6736 101414 -6652
rect 100794 -6972 100826 -6736
rect 101062 -6972 101146 -6736
rect 101382 -6972 101414 -6736
rect 100794 -7964 101414 -6972
rect 105294 286954 105914 298000
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 214954 105914 250398
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 105294 142954 105914 178398
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7376 105914 34398
rect 105294 -7612 105326 -7376
rect 105562 -7612 105646 -7376
rect 105882 -7612 105914 -7376
rect 105294 -7696 105914 -7612
rect 105294 -7932 105326 -7696
rect 105562 -7932 105646 -7696
rect 105882 -7932 105914 -7696
rect 105294 -7964 105914 -7932
rect 109794 291454 110414 298000
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -656 110414 2898
rect 109794 -892 109826 -656
rect 110062 -892 110146 -656
rect 110382 -892 110414 -656
rect 109794 -976 110414 -892
rect 109794 -1212 109826 -976
rect 110062 -1212 110146 -976
rect 110382 -1212 110414 -976
rect 109794 -7964 110414 -1212
rect 114294 295954 114914 298000
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 259954 114914 295398
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 223954 114914 259398
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 151954 114914 187398
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114294 115954 114914 151398
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1616 114914 7398
rect 114294 -1852 114326 -1616
rect 114562 -1852 114646 -1616
rect 114882 -1852 114914 -1616
rect 114294 -1936 114914 -1852
rect 114294 -2172 114326 -1936
rect 114562 -2172 114646 -1936
rect 114882 -2172 114914 -1936
rect 114294 -7964 114914 -2172
rect 118794 264454 119414 298000
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118794 228454 119414 263898
rect 118794 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 119414 228454
rect 118794 228134 119414 228218
rect 118794 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 119414 228134
rect 118794 192454 119414 227898
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 120454 119414 155898
rect 118794 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 119414 120454
rect 118794 120134 119414 120218
rect 118794 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 119414 120134
rect 118794 84454 119414 119898
rect 118794 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 119414 84454
rect 118794 84134 119414 84218
rect 118794 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 119414 84134
rect 118794 48454 119414 83898
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2576 119414 11898
rect 118794 -2812 118826 -2576
rect 119062 -2812 119146 -2576
rect 119382 -2812 119414 -2576
rect 118794 -2896 119414 -2812
rect 118794 -3132 118826 -2896
rect 119062 -3132 119146 -2896
rect 119382 -3132 119414 -2896
rect 118794 -7964 119414 -3132
rect 123294 268954 123914 298000
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 232954 123914 268398
rect 123294 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 123914 232954
rect 123294 232634 123914 232718
rect 123294 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 123914 232634
rect 123294 196954 123914 232398
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 123294 124954 123914 160398
rect 123294 124718 123326 124954
rect 123562 124718 123646 124954
rect 123882 124718 123914 124954
rect 123294 124634 123914 124718
rect 123294 124398 123326 124634
rect 123562 124398 123646 124634
rect 123882 124398 123914 124634
rect 123294 88954 123914 124398
rect 123294 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 123914 88954
rect 123294 88634 123914 88718
rect 123294 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 123914 88634
rect 123294 52954 123914 88398
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3536 123914 16398
rect 123294 -3772 123326 -3536
rect 123562 -3772 123646 -3536
rect 123882 -3772 123914 -3536
rect 123294 -3856 123914 -3772
rect 123294 -4092 123326 -3856
rect 123562 -4092 123646 -3856
rect 123882 -4092 123914 -3856
rect 123294 -7964 123914 -4092
rect 127794 273454 128414 298000
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4496 128414 20898
rect 127794 -4732 127826 -4496
rect 128062 -4732 128146 -4496
rect 128382 -4732 128414 -4496
rect 127794 -4816 128414 -4732
rect 127794 -5052 127826 -4816
rect 128062 -5052 128146 -4816
rect 128382 -5052 128414 -4816
rect 127794 -7964 128414 -5052
rect 132294 277954 132914 298000
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 241954 132914 277398
rect 132294 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 132914 241954
rect 132294 241634 132914 241718
rect 132294 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 132914 241634
rect 132294 205954 132914 241398
rect 132294 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 132914 205954
rect 132294 205634 132914 205718
rect 132294 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 132914 205634
rect 132294 169954 132914 205398
rect 132294 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 132914 169954
rect 132294 169634 132914 169718
rect 132294 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 132914 169634
rect 132294 133954 132914 169398
rect 132294 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 132914 133954
rect 132294 133634 132914 133718
rect 132294 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 132914 133634
rect 132294 97954 132914 133398
rect 132294 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 132914 97954
rect 132294 97634 132914 97718
rect 132294 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 132914 97634
rect 132294 61954 132914 97398
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5456 132914 25398
rect 132294 -5692 132326 -5456
rect 132562 -5692 132646 -5456
rect 132882 -5692 132914 -5456
rect 132294 -5776 132914 -5692
rect 132294 -6012 132326 -5776
rect 132562 -6012 132646 -5776
rect 132882 -6012 132914 -5776
rect 132294 -7964 132914 -6012
rect 136794 282454 137414 298000
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 246454 137414 281898
rect 136794 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 137414 246454
rect 136794 246134 137414 246218
rect 136794 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 137414 246134
rect 136794 210454 137414 245898
rect 136794 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 137414 210454
rect 136794 210134 137414 210218
rect 136794 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 137414 210134
rect 136794 174454 137414 209898
rect 136794 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 137414 174454
rect 136794 174134 137414 174218
rect 136794 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 137414 174134
rect 136794 138454 137414 173898
rect 136794 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 137414 138454
rect 136794 138134 137414 138218
rect 136794 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 137414 138134
rect 136794 102454 137414 137898
rect 136794 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 137414 102454
rect 136794 102134 137414 102218
rect 136794 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 137414 102134
rect 136794 66454 137414 101898
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6416 137414 29898
rect 136794 -6652 136826 -6416
rect 137062 -6652 137146 -6416
rect 137382 -6652 137414 -6416
rect 136794 -6736 137414 -6652
rect 136794 -6972 136826 -6736
rect 137062 -6972 137146 -6736
rect 137382 -6972 137414 -6736
rect 136794 -7964 137414 -6972
rect 141294 286954 141914 298000
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 214954 141914 250398
rect 141294 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 141914 214954
rect 141294 214634 141914 214718
rect 141294 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 141914 214634
rect 141294 178954 141914 214398
rect 141294 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 141914 178954
rect 141294 178634 141914 178718
rect 141294 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 141914 178634
rect 141294 142954 141914 178398
rect 141294 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 141914 142954
rect 141294 142634 141914 142718
rect 141294 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 141914 142634
rect 141294 106954 141914 142398
rect 141294 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 141914 106954
rect 141294 106634 141914 106718
rect 141294 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 141914 106634
rect 141294 70954 141914 106398
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7376 141914 34398
rect 141294 -7612 141326 -7376
rect 141562 -7612 141646 -7376
rect 141882 -7612 141914 -7376
rect 141294 -7696 141914 -7612
rect 141294 -7932 141326 -7696
rect 141562 -7932 141646 -7696
rect 141882 -7932 141914 -7696
rect 141294 -7964 141914 -7932
rect 145794 291454 146414 298000
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -656 146414 2898
rect 145794 -892 145826 -656
rect 146062 -892 146146 -656
rect 146382 -892 146414 -656
rect 145794 -976 146414 -892
rect 145794 -1212 145826 -976
rect 146062 -1212 146146 -976
rect 146382 -1212 146414 -976
rect 145794 -7964 146414 -1212
rect 150294 295954 150914 298000
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 223954 150914 259398
rect 150294 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 150914 223954
rect 150294 223634 150914 223718
rect 150294 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 150914 223634
rect 150294 187954 150914 223398
rect 150294 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 150914 187954
rect 150294 187634 150914 187718
rect 150294 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 150914 187634
rect 150294 151954 150914 187398
rect 150294 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 150914 151954
rect 150294 151634 150914 151718
rect 150294 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 150914 151634
rect 150294 115954 150914 151398
rect 150294 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 150914 115954
rect 150294 115634 150914 115718
rect 150294 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 150914 115634
rect 150294 79954 150914 115398
rect 150294 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 150914 79954
rect 150294 79634 150914 79718
rect 150294 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 150914 79634
rect 150294 43954 150914 79398
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1616 150914 7398
rect 150294 -1852 150326 -1616
rect 150562 -1852 150646 -1616
rect 150882 -1852 150914 -1616
rect 150294 -1936 150914 -1852
rect 150294 -2172 150326 -1936
rect 150562 -2172 150646 -1936
rect 150882 -2172 150914 -1936
rect 150294 -7964 150914 -2172
rect 154794 264454 155414 298000
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 228454 155414 263898
rect 154794 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 155414 228454
rect 154794 228134 155414 228218
rect 154794 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 155414 228134
rect 154794 192454 155414 227898
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 154794 156454 155414 191898
rect 154794 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 155414 156454
rect 154794 156134 155414 156218
rect 154794 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 155414 156134
rect 154794 120454 155414 155898
rect 154794 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 155414 120454
rect 154794 120134 155414 120218
rect 154794 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 155414 120134
rect 154794 84454 155414 119898
rect 154794 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 155414 84454
rect 154794 84134 155414 84218
rect 154794 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 155414 84134
rect 154794 48454 155414 83898
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2576 155414 11898
rect 154794 -2812 154826 -2576
rect 155062 -2812 155146 -2576
rect 155382 -2812 155414 -2576
rect 154794 -2896 155414 -2812
rect 154794 -3132 154826 -2896
rect 155062 -3132 155146 -2896
rect 155382 -3132 155414 -2896
rect 154794 -7964 155414 -3132
rect 159294 268954 159914 298000
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 232954 159914 268398
rect 159294 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 159914 232954
rect 159294 232634 159914 232718
rect 159294 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 159914 232634
rect 159294 196954 159914 232398
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 159294 160954 159914 196398
rect 159294 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 159914 160954
rect 159294 160634 159914 160718
rect 159294 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 159914 160634
rect 159294 124954 159914 160398
rect 159294 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 159914 124954
rect 159294 124634 159914 124718
rect 159294 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 159914 124634
rect 159294 88954 159914 124398
rect 159294 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 159914 88954
rect 159294 88634 159914 88718
rect 159294 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 159914 88634
rect 159294 52954 159914 88398
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3536 159914 16398
rect 159294 -3772 159326 -3536
rect 159562 -3772 159646 -3536
rect 159882 -3772 159914 -3536
rect 159294 -3856 159914 -3772
rect 159294 -4092 159326 -3856
rect 159562 -4092 159646 -3856
rect 159882 -4092 159914 -3856
rect 159294 -7964 159914 -4092
rect 163794 273454 164414 298000
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4496 164414 20898
rect 163794 -4732 163826 -4496
rect 164062 -4732 164146 -4496
rect 164382 -4732 164414 -4496
rect 163794 -4816 164414 -4732
rect 163794 -5052 163826 -4816
rect 164062 -5052 164146 -4816
rect 164382 -5052 164414 -4816
rect 163794 -7964 164414 -5052
rect 168294 277954 168914 298000
rect 169526 297941 169586 301547
rect 169523 297940 169589 297941
rect 169523 297876 169524 297940
rect 169588 297876 169589 297940
rect 169523 297875 169589 297876
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 241954 168914 277398
rect 168294 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 168914 241954
rect 168294 241634 168914 241718
rect 168294 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 168914 241634
rect 168294 205954 168914 241398
rect 168294 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 168914 205954
rect 168294 205634 168914 205718
rect 168294 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 168914 205634
rect 168294 169954 168914 205398
rect 168294 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 168914 169954
rect 168294 169634 168914 169718
rect 168294 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 168914 169634
rect 168294 133954 168914 169398
rect 168294 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 168914 133954
rect 168294 133634 168914 133718
rect 168294 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 168914 133634
rect 168294 97954 168914 133398
rect 168294 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 168914 97954
rect 168294 97634 168914 97718
rect 168294 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 168914 97634
rect 168294 61954 168914 97398
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5456 168914 25398
rect 168294 -5692 168326 -5456
rect 168562 -5692 168646 -5456
rect 168882 -5692 168914 -5456
rect 168294 -5776 168914 -5692
rect 168294 -6012 168326 -5776
rect 168562 -6012 168646 -5776
rect 168882 -6012 168914 -5776
rect 168294 -7964 168914 -6012
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 246454 173414 281898
rect 172794 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 173414 246454
rect 172794 246134 173414 246218
rect 172794 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 173414 246134
rect 172794 210454 173414 245898
rect 172794 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 173414 210454
rect 172794 210134 173414 210218
rect 172794 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 173414 210134
rect 172794 174454 173414 209898
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 172794 138454 173414 173898
rect 172794 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 173414 138454
rect 172794 138134 173414 138218
rect 172794 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 173414 138134
rect 172794 102454 173414 137898
rect 172794 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 173414 102454
rect 172794 102134 173414 102218
rect 172794 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 173414 102134
rect 172794 66454 173414 101898
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6416 173414 29898
rect 172794 -6652 172826 -6416
rect 173062 -6652 173146 -6416
rect 173382 -6652 173414 -6416
rect 172794 -6736 173414 -6652
rect 172794 -6972 172826 -6736
rect 173062 -6972 173146 -6736
rect 173382 -6972 173414 -6736
rect 172794 -7964 173414 -6972
rect 177294 711868 177914 711900
rect 177294 711632 177326 711868
rect 177562 711632 177646 711868
rect 177882 711632 177914 711868
rect 177294 711548 177914 711632
rect 177294 711312 177326 711548
rect 177562 711312 177646 711548
rect 177882 711312 177914 711548
rect 177294 682954 177914 711312
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 214954 177914 250398
rect 177294 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 177914 214954
rect 177294 214634 177914 214718
rect 177294 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 177914 214634
rect 177294 178954 177914 214398
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 106954 177914 142398
rect 177294 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 177914 106954
rect 177294 106634 177914 106718
rect 177294 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 177914 106634
rect 177294 70954 177914 106398
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7376 177914 34398
rect 177294 -7612 177326 -7376
rect 177562 -7612 177646 -7376
rect 177882 -7612 177914 -7376
rect 177294 -7696 177914 -7612
rect 177294 -7932 177326 -7696
rect 177562 -7932 177646 -7696
rect 177882 -7932 177914 -7696
rect 177294 -7964 177914 -7932
rect 181794 705148 182414 711900
rect 181794 704912 181826 705148
rect 182062 704912 182146 705148
rect 182382 704912 182414 705148
rect 181794 704828 182414 704912
rect 181794 704592 181826 704828
rect 182062 704592 182146 704828
rect 182382 704592 182414 704828
rect 181794 687454 182414 704592
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -656 182414 2898
rect 181794 -892 181826 -656
rect 182062 -892 182146 -656
rect 182382 -892 182414 -656
rect 181794 -976 182414 -892
rect 181794 -1212 181826 -976
rect 182062 -1212 182146 -976
rect 182382 -1212 182414 -976
rect 181794 -7964 182414 -1212
rect 186294 706108 186914 711900
rect 186294 705872 186326 706108
rect 186562 705872 186646 706108
rect 186882 705872 186914 706108
rect 186294 705788 186914 705872
rect 186294 705552 186326 705788
rect 186562 705552 186646 705788
rect 186882 705552 186914 705788
rect 186294 691954 186914 705552
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 259954 186914 295398
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 223954 186914 259398
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 187954 186914 223398
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 115954 186914 151398
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 186294 79954 186914 115398
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 186294 79634 186914 79718
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1616 186914 7398
rect 186294 -1852 186326 -1616
rect 186562 -1852 186646 -1616
rect 186882 -1852 186914 -1616
rect 186294 -1936 186914 -1852
rect 186294 -2172 186326 -1936
rect 186562 -2172 186646 -1936
rect 186882 -2172 186914 -1936
rect 186294 -7964 186914 -2172
rect 190794 707068 191414 711900
rect 190794 706832 190826 707068
rect 191062 706832 191146 707068
rect 191382 706832 191414 707068
rect 190794 706748 191414 706832
rect 190794 706512 190826 706748
rect 191062 706512 191146 706748
rect 191382 706512 191414 706748
rect 190794 696454 191414 706512
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 228454 191414 263898
rect 190794 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 191414 228454
rect 190794 228134 191414 228218
rect 190794 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 191414 228134
rect 190794 192454 191414 227898
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 120454 191414 155898
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 84454 191414 119898
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2576 191414 11898
rect 190794 -2812 190826 -2576
rect 191062 -2812 191146 -2576
rect 191382 -2812 191414 -2576
rect 190794 -2896 191414 -2812
rect 190794 -3132 190826 -2896
rect 191062 -3132 191146 -2896
rect 191382 -3132 191414 -2896
rect 190794 -7964 191414 -3132
rect 195294 708028 195914 711900
rect 195294 707792 195326 708028
rect 195562 707792 195646 708028
rect 195882 707792 195914 708028
rect 195294 707708 195914 707792
rect 195294 707472 195326 707708
rect 195562 707472 195646 707708
rect 195882 707472 195914 707708
rect 195294 700954 195914 707472
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 195294 232954 195914 268398
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 196954 195914 232398
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3536 195914 16398
rect 195294 -3772 195326 -3536
rect 195562 -3772 195646 -3536
rect 195882 -3772 195914 -3536
rect 195294 -3856 195914 -3772
rect 195294 -4092 195326 -3856
rect 195562 -4092 195646 -3856
rect 195882 -4092 195914 -3856
rect 195294 -7964 195914 -4092
rect 199794 708988 200414 711900
rect 199794 708752 199826 708988
rect 200062 708752 200146 708988
rect 200382 708752 200414 708988
rect 199794 708668 200414 708752
rect 199794 708432 199826 708668
rect 200062 708432 200146 708668
rect 200382 708432 200414 708668
rect 199794 669454 200414 708432
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4496 200414 20898
rect 199794 -4732 199826 -4496
rect 200062 -4732 200146 -4496
rect 200382 -4732 200414 -4496
rect 199794 -4816 200414 -4732
rect 199794 -5052 199826 -4816
rect 200062 -5052 200146 -4816
rect 200382 -5052 200414 -4816
rect 199794 -7964 200414 -5052
rect 204294 709948 204914 711900
rect 204294 709712 204326 709948
rect 204562 709712 204646 709948
rect 204882 709712 204914 709948
rect 204294 709628 204914 709712
rect 204294 709392 204326 709628
rect 204562 709392 204646 709628
rect 204882 709392 204914 709628
rect 204294 673954 204914 709392
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 241954 204914 277398
rect 204294 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 204914 241954
rect 204294 241634 204914 241718
rect 204294 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 204914 241634
rect 204294 205954 204914 241398
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5456 204914 25398
rect 204294 -5692 204326 -5456
rect 204562 -5692 204646 -5456
rect 204882 -5692 204914 -5456
rect 204294 -5776 204914 -5692
rect 204294 -6012 204326 -5776
rect 204562 -6012 204646 -5776
rect 204882 -6012 204914 -5776
rect 204294 -7964 204914 -6012
rect 208794 710908 209414 711900
rect 208794 710672 208826 710908
rect 209062 710672 209146 710908
rect 209382 710672 209414 710908
rect 208794 710588 209414 710672
rect 208794 710352 208826 710588
rect 209062 710352 209146 710588
rect 209382 710352 209414 710588
rect 208794 678454 209414 710352
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 246454 209414 281898
rect 208794 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 209414 246454
rect 208794 246134 209414 246218
rect 208794 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 209414 246134
rect 208794 210454 209414 245898
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6416 209414 29898
rect 208794 -6652 208826 -6416
rect 209062 -6652 209146 -6416
rect 209382 -6652 209414 -6416
rect 208794 -6736 209414 -6652
rect 208794 -6972 208826 -6736
rect 209062 -6972 209146 -6736
rect 209382 -6972 209414 -6736
rect 208794 -7964 209414 -6972
rect 213294 711868 213914 711900
rect 213294 711632 213326 711868
rect 213562 711632 213646 711868
rect 213882 711632 213914 711868
rect 213294 711548 213914 711632
rect 213294 711312 213326 711548
rect 213562 711312 213646 711548
rect 213882 711312 213914 711548
rect 213294 682954 213914 711312
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 217794 705148 218414 711900
rect 217794 704912 217826 705148
rect 218062 704912 218146 705148
rect 218382 704912 218414 705148
rect 217794 704828 218414 704912
rect 217794 704592 217826 704828
rect 218062 704592 218146 704828
rect 218382 704592 218414 704828
rect 217794 687454 218414 704592
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 565308 218414 578898
rect 222294 706108 222914 711900
rect 222294 705872 222326 706108
rect 222562 705872 222646 706108
rect 222882 705872 222914 706108
rect 222294 705788 222914 705872
rect 222294 705552 222326 705788
rect 222562 705552 222646 705788
rect 222882 705552 222914 705788
rect 222294 691954 222914 705552
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 565308 222914 583398
rect 226794 707068 227414 711900
rect 226794 706832 226826 707068
rect 227062 706832 227146 707068
rect 227382 706832 227414 707068
rect 226794 706748 227414 706832
rect 226794 706512 226826 706748
rect 227062 706512 227146 706748
rect 227382 706512 227414 706748
rect 226794 696454 227414 706512
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 565308 227414 587898
rect 231294 708028 231914 711900
rect 231294 707792 231326 708028
rect 231562 707792 231646 708028
rect 231882 707792 231914 708028
rect 231294 707708 231914 707792
rect 231294 707472 231326 707708
rect 231562 707472 231646 707708
rect 231882 707472 231914 707708
rect 231294 700954 231914 707472
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 565308 231914 592398
rect 235794 708988 236414 711900
rect 235794 708752 235826 708988
rect 236062 708752 236146 708988
rect 236382 708752 236414 708988
rect 235794 708668 236414 708752
rect 235794 708432 235826 708668
rect 236062 708432 236146 708668
rect 236382 708432 236414 708668
rect 235794 669454 236414 708432
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 565308 236414 596898
rect 240294 709948 240914 711900
rect 240294 709712 240326 709948
rect 240562 709712 240646 709948
rect 240882 709712 240914 709948
rect 240294 709628 240914 709712
rect 240294 709392 240326 709628
rect 240562 709392 240646 709628
rect 240882 709392 240914 709628
rect 240294 673954 240914 709392
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 565308 240914 565398
rect 244794 710908 245414 711900
rect 244794 710672 244826 710908
rect 245062 710672 245146 710908
rect 245382 710672 245414 710908
rect 244794 710588 245414 710672
rect 244794 710352 244826 710588
rect 245062 710352 245146 710588
rect 245382 710352 245414 710588
rect 244794 678454 245414 710352
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 565308 245414 569898
rect 249294 711868 249914 711900
rect 249294 711632 249326 711868
rect 249562 711632 249646 711868
rect 249882 711632 249914 711868
rect 249294 711548 249914 711632
rect 249294 711312 249326 711548
rect 249562 711312 249646 711548
rect 249882 711312 249914 711548
rect 249294 682954 249914 711312
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 565308 249914 574398
rect 253794 705148 254414 711900
rect 253794 704912 253826 705148
rect 254062 704912 254146 705148
rect 254382 704912 254414 705148
rect 253794 704828 254414 704912
rect 253794 704592 253826 704828
rect 254062 704592 254146 704828
rect 254382 704592 254414 704828
rect 253794 687454 254414 704592
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 565308 254414 578898
rect 258294 706108 258914 711900
rect 258294 705872 258326 706108
rect 258562 705872 258646 706108
rect 258882 705872 258914 706108
rect 258294 705788 258914 705872
rect 258294 705552 258326 705788
rect 258562 705552 258646 705788
rect 258882 705552 258914 705788
rect 258294 691954 258914 705552
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 565308 258914 583398
rect 262794 707068 263414 711900
rect 262794 706832 262826 707068
rect 263062 706832 263146 707068
rect 263382 706832 263414 707068
rect 262794 706748 263414 706832
rect 262794 706512 262826 706748
rect 263062 706512 263146 706748
rect 263382 706512 263414 706748
rect 262794 696454 263414 706512
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 565308 263414 587898
rect 267294 708028 267914 711900
rect 267294 707792 267326 708028
rect 267562 707792 267646 708028
rect 267882 707792 267914 708028
rect 267294 707708 267914 707792
rect 267294 707472 267326 707708
rect 267562 707472 267646 707708
rect 267882 707472 267914 707708
rect 267294 700954 267914 707472
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 565308 267914 592398
rect 271794 708988 272414 711900
rect 271794 708752 271826 708988
rect 272062 708752 272146 708988
rect 272382 708752 272414 708988
rect 271794 708668 272414 708752
rect 271794 708432 271826 708668
rect 272062 708432 272146 708668
rect 272382 708432 272414 708668
rect 271794 669454 272414 708432
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 565308 272414 596898
rect 276294 709948 276914 711900
rect 276294 709712 276326 709948
rect 276562 709712 276646 709948
rect 276882 709712 276914 709948
rect 276294 709628 276914 709712
rect 276294 709392 276326 709628
rect 276562 709392 276646 709628
rect 276882 709392 276914 709628
rect 276294 673954 276914 709392
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 565308 276914 565398
rect 280794 710908 281414 711900
rect 280794 710672 280826 710908
rect 281062 710672 281146 710908
rect 281382 710672 281414 710908
rect 280794 710588 281414 710672
rect 280794 710352 280826 710588
rect 281062 710352 281146 710588
rect 281382 710352 281414 710588
rect 280794 678454 281414 710352
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 565308 281414 569898
rect 285294 711868 285914 711900
rect 285294 711632 285326 711868
rect 285562 711632 285646 711868
rect 285882 711632 285914 711868
rect 285294 711548 285914 711632
rect 285294 711312 285326 711548
rect 285562 711312 285646 711548
rect 285882 711312 285914 711548
rect 285294 682954 285914 711312
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 565308 285914 574398
rect 289794 705148 290414 711900
rect 289794 704912 289826 705148
rect 290062 704912 290146 705148
rect 290382 704912 290414 705148
rect 289794 704828 290414 704912
rect 289794 704592 289826 704828
rect 290062 704592 290146 704828
rect 290382 704592 290414 704828
rect 289794 687454 290414 704592
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 565308 290414 578898
rect 294294 706108 294914 711900
rect 294294 705872 294326 706108
rect 294562 705872 294646 706108
rect 294882 705872 294914 706108
rect 294294 705788 294914 705872
rect 294294 705552 294326 705788
rect 294562 705552 294646 705788
rect 294882 705552 294914 705788
rect 294294 691954 294914 705552
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 565308 294914 583398
rect 298794 707068 299414 711900
rect 298794 706832 298826 707068
rect 299062 706832 299146 707068
rect 299382 706832 299414 707068
rect 298794 706748 299414 706832
rect 298794 706512 298826 706748
rect 299062 706512 299146 706748
rect 299382 706512 299414 706748
rect 298794 696454 299414 706512
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 565308 299414 587898
rect 303294 708028 303914 711900
rect 303294 707792 303326 708028
rect 303562 707792 303646 708028
rect 303882 707792 303914 708028
rect 303294 707708 303914 707792
rect 303294 707472 303326 707708
rect 303562 707472 303646 707708
rect 303882 707472 303914 707708
rect 303294 700954 303914 707472
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 565308 303914 592398
rect 307794 708988 308414 711900
rect 307794 708752 307826 708988
rect 308062 708752 308146 708988
rect 308382 708752 308414 708988
rect 307794 708668 308414 708752
rect 307794 708432 307826 708668
rect 308062 708432 308146 708668
rect 308382 708432 308414 708668
rect 307794 669454 308414 708432
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 565308 308414 596898
rect 312294 709948 312914 711900
rect 312294 709712 312326 709948
rect 312562 709712 312646 709948
rect 312882 709712 312914 709948
rect 312294 709628 312914 709712
rect 312294 709392 312326 709628
rect 312562 709392 312646 709628
rect 312882 709392 312914 709628
rect 312294 673954 312914 709392
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 565308 312914 565398
rect 316794 710908 317414 711900
rect 316794 710672 316826 710908
rect 317062 710672 317146 710908
rect 317382 710672 317414 710908
rect 316794 710588 317414 710672
rect 316794 710352 316826 710588
rect 317062 710352 317146 710588
rect 317382 710352 317414 710588
rect 316794 678454 317414 710352
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 565308 317414 569898
rect 321294 711868 321914 711900
rect 321294 711632 321326 711868
rect 321562 711632 321646 711868
rect 321882 711632 321914 711868
rect 321294 711548 321914 711632
rect 321294 711312 321326 711548
rect 321562 711312 321646 711548
rect 321882 711312 321914 711548
rect 321294 682954 321914 711312
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 565308 321914 574398
rect 325794 705148 326414 711900
rect 325794 704912 325826 705148
rect 326062 704912 326146 705148
rect 326382 704912 326414 705148
rect 325794 704828 326414 704912
rect 325794 704592 325826 704828
rect 326062 704592 326146 704828
rect 326382 704592 326414 704828
rect 325794 687454 326414 704592
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 565308 326414 578898
rect 330294 706108 330914 711900
rect 330294 705872 330326 706108
rect 330562 705872 330646 706108
rect 330882 705872 330914 706108
rect 330294 705788 330914 705872
rect 330294 705552 330326 705788
rect 330562 705552 330646 705788
rect 330882 705552 330914 705788
rect 330294 691954 330914 705552
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 565308 330914 583398
rect 334794 707068 335414 711900
rect 334794 706832 334826 707068
rect 335062 706832 335146 707068
rect 335382 706832 335414 707068
rect 334794 706748 335414 706832
rect 334794 706512 334826 706748
rect 335062 706512 335146 706748
rect 335382 706512 335414 706748
rect 334794 696454 335414 706512
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 565308 335414 587898
rect 339294 708028 339914 711900
rect 339294 707792 339326 708028
rect 339562 707792 339646 708028
rect 339882 707792 339914 708028
rect 339294 707708 339914 707792
rect 339294 707472 339326 707708
rect 339562 707472 339646 707708
rect 339882 707472 339914 707708
rect 339294 700954 339914 707472
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 565308 339914 592398
rect 343794 708988 344414 711900
rect 343794 708752 343826 708988
rect 344062 708752 344146 708988
rect 344382 708752 344414 708988
rect 343794 708668 344414 708752
rect 343794 708432 343826 708668
rect 344062 708432 344146 708668
rect 344382 708432 344414 708668
rect 343794 669454 344414 708432
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 565308 344414 596898
rect 348294 709948 348914 711900
rect 348294 709712 348326 709948
rect 348562 709712 348646 709948
rect 348882 709712 348914 709948
rect 348294 709628 348914 709712
rect 348294 709392 348326 709628
rect 348562 709392 348646 709628
rect 348882 709392 348914 709628
rect 348294 673954 348914 709392
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 565308 348914 565398
rect 352794 710908 353414 711900
rect 352794 710672 352826 710908
rect 353062 710672 353146 710908
rect 353382 710672 353414 710908
rect 352794 710588 353414 710672
rect 352794 710352 352826 710588
rect 353062 710352 353146 710588
rect 353382 710352 353414 710588
rect 352794 678454 353414 710352
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 565308 353414 569898
rect 357294 711868 357914 711900
rect 357294 711632 357326 711868
rect 357562 711632 357646 711868
rect 357882 711632 357914 711868
rect 357294 711548 357914 711632
rect 357294 711312 357326 711548
rect 357562 711312 357646 711548
rect 357882 711312 357914 711548
rect 357294 682954 357914 711312
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 565308 357914 574398
rect 361794 705148 362414 711900
rect 361794 704912 361826 705148
rect 362062 704912 362146 705148
rect 362382 704912 362414 705148
rect 361794 704828 362414 704912
rect 361794 704592 361826 704828
rect 362062 704592 362146 704828
rect 362382 704592 362414 704828
rect 361794 687454 362414 704592
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 220272 547954 220620 547986
rect 220272 547718 220328 547954
rect 220564 547718 220620 547954
rect 220272 547634 220620 547718
rect 220272 547398 220328 547634
rect 220564 547398 220620 547634
rect 220272 547366 220620 547398
rect 356000 547954 356348 547986
rect 356000 547718 356056 547954
rect 356292 547718 356348 547954
rect 356000 547634 356348 547718
rect 356000 547398 356056 547634
rect 356292 547398 356348 547634
rect 356000 547366 356348 547398
rect 220952 543454 221300 543486
rect 220952 543218 221008 543454
rect 221244 543218 221300 543454
rect 220952 543134 221300 543218
rect 220952 542898 221008 543134
rect 221244 542898 221300 543134
rect 220952 542866 221300 542898
rect 355320 543454 355668 543486
rect 355320 543218 355376 543454
rect 355612 543218 355668 543454
rect 355320 543134 355668 543218
rect 355320 542898 355376 543134
rect 355612 542898 355668 543134
rect 355320 542866 355668 542898
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 220272 511954 220620 511986
rect 220272 511718 220328 511954
rect 220564 511718 220620 511954
rect 220272 511634 220620 511718
rect 220272 511398 220328 511634
rect 220564 511398 220620 511634
rect 220272 511366 220620 511398
rect 356000 511954 356348 511986
rect 356000 511718 356056 511954
rect 356292 511718 356348 511954
rect 356000 511634 356348 511718
rect 356000 511398 356056 511634
rect 356292 511398 356348 511634
rect 356000 511366 356348 511398
rect 220952 507454 221300 507486
rect 220952 507218 221008 507454
rect 221244 507218 221300 507454
rect 220952 507134 221300 507218
rect 220952 506898 221008 507134
rect 221244 506898 221300 507134
rect 220952 506866 221300 506898
rect 355320 507454 355668 507486
rect 355320 507218 355376 507454
rect 355612 507218 355668 507454
rect 355320 507134 355668 507218
rect 355320 506898 355376 507134
rect 355612 506898 355668 507134
rect 355320 506866 355668 506898
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 236056 479770 236116 480080
rect 237144 479770 237204 480080
rect 238232 479770 238292 480080
rect 239592 479770 239652 480080
rect 240544 479770 240604 480080
rect 241768 479770 241828 480080
rect 243128 479770 243188 480080
rect 236056 479710 236194 479770
rect 237144 479710 237298 479770
rect 238232 479710 238402 479770
rect 239592 479710 239690 479770
rect 240544 479710 240610 479770
rect 241768 479710 241898 479770
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 217794 471454 218414 478000
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 216075 444956 216141 444957
rect 216075 444892 216076 444956
rect 216140 444892 216141 444956
rect 216075 444891 216141 444892
rect 214603 444820 214669 444821
rect 214603 444756 214604 444820
rect 214668 444756 214669 444820
rect 214603 444755 214669 444756
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 214419 284884 214485 284885
rect 214419 284820 214420 284884
rect 214484 284820 214485 284884
rect 214419 284819 214485 284820
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 214954 213914 250398
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7376 213914 34398
rect 214422 3365 214482 284819
rect 214606 162893 214666 444755
rect 215891 441828 215957 441829
rect 215891 441764 215892 441828
rect 215956 441764 215957 441828
rect 215891 441763 215957 441764
rect 215155 303244 215221 303245
rect 215155 303180 215156 303244
rect 215220 303180 215221 303244
rect 215155 303179 215221 303180
rect 214603 162892 214669 162893
rect 214603 162828 214604 162892
rect 214668 162828 214669 162892
rect 214603 162827 214669 162828
rect 215158 3501 215218 303179
rect 215894 5677 215954 441763
rect 216078 214029 216138 444891
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217363 305828 217429 305829
rect 217363 305764 217364 305828
rect 217428 305764 217429 305828
rect 217363 305763 217429 305764
rect 217179 305692 217245 305693
rect 217179 305628 217180 305692
rect 217244 305628 217245 305692
rect 217179 305627 217245 305628
rect 216259 303380 216325 303381
rect 216259 303316 216260 303380
rect 216324 303316 216325 303380
rect 216259 303315 216325 303316
rect 216075 214028 216141 214029
rect 216075 213964 216076 214028
rect 216140 213964 216141 214028
rect 216075 213963 216141 213964
rect 216262 158269 216322 303315
rect 216995 297804 217061 297805
rect 216995 297740 216996 297804
rect 217060 297740 217061 297804
rect 216995 297739 217061 297740
rect 216443 255916 216509 255917
rect 216443 255852 216444 255916
rect 216508 255852 216509 255916
rect 216443 255851 216509 255852
rect 216259 158268 216325 158269
rect 216259 158204 216260 158268
rect 216324 158204 216325 158268
rect 216259 158203 216325 158204
rect 215891 5676 215957 5677
rect 215891 5612 215892 5676
rect 215956 5612 215957 5676
rect 215891 5611 215957 5612
rect 216446 3501 216506 255851
rect 216998 155413 217058 297739
rect 217182 157997 217242 305627
rect 217366 158133 217426 305763
rect 217794 291454 218414 326898
rect 222294 475954 222914 478000
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 218835 306236 218901 306237
rect 218835 306172 218836 306236
rect 218900 306172 218901 306236
rect 218835 306171 218901 306172
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217547 250476 217613 250477
rect 217547 250412 217548 250476
rect 217612 250412 217613 250476
rect 217547 250411 217613 250412
rect 217363 158132 217429 158133
rect 217363 158068 217364 158132
rect 217428 158068 217429 158132
rect 217363 158067 217429 158068
rect 217179 157996 217245 157997
rect 217179 157932 217180 157996
rect 217244 157932 217245 157996
rect 217179 157931 217245 157932
rect 216995 155412 217061 155413
rect 216995 155348 216996 155412
rect 217060 155348 217061 155412
rect 216995 155347 217061 155348
rect 217550 3501 217610 250411
rect 217794 245308 218414 254898
rect 218651 193220 218717 193221
rect 218651 193156 218652 193220
rect 218716 193156 218717 193220
rect 218651 193155 218717 193156
rect 217794 147454 218414 158000
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 215155 3500 215221 3501
rect 215155 3436 215156 3500
rect 215220 3436 215221 3500
rect 215155 3435 215221 3436
rect 216443 3500 216509 3501
rect 216443 3436 216444 3500
rect 216508 3436 216509 3500
rect 216443 3435 216509 3436
rect 217547 3500 217613 3501
rect 217547 3436 217548 3500
rect 217612 3436 217613 3500
rect 217547 3435 217613 3436
rect 217794 3454 218414 38898
rect 218654 3501 218714 193155
rect 218838 158677 218898 306171
rect 219019 306100 219085 306101
rect 219019 306036 219020 306100
rect 219084 306036 219085 306100
rect 219019 306035 219085 306036
rect 218835 158676 218901 158677
rect 218835 158612 218836 158676
rect 218900 158612 218901 158676
rect 218835 158611 218901 158612
rect 219022 158541 219082 306035
rect 219203 305964 219269 305965
rect 219203 305900 219204 305964
rect 219268 305900 219269 305964
rect 219203 305899 219269 305900
rect 219019 158540 219085 158541
rect 219019 158476 219020 158540
rect 219084 158476 219085 158540
rect 219019 158475 219085 158476
rect 219206 158405 219266 305899
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 245308 222914 259398
rect 226794 444454 227414 478000
rect 236134 476781 236194 479710
rect 236131 476780 236197 476781
rect 236131 476716 236132 476780
rect 236196 476716 236197 476780
rect 236131 476715 236197 476716
rect 237238 476237 237298 479710
rect 238342 477325 238402 479710
rect 238339 477324 238405 477325
rect 238339 477260 238340 477324
rect 238404 477260 238405 477324
rect 238339 477259 238405 477260
rect 239630 476917 239690 479710
rect 240550 476917 240610 479710
rect 241838 477189 241898 479710
rect 243126 479710 243188 479770
rect 244216 479770 244276 480080
rect 245440 479770 245500 480080
rect 246528 479770 246588 480080
rect 247616 479770 247676 480080
rect 248296 479770 248356 480080
rect 248704 479770 248764 480080
rect 244216 479710 244290 479770
rect 245440 479710 245578 479770
rect 246528 479710 246682 479770
rect 247616 479710 247786 479770
rect 241835 477188 241901 477189
rect 241835 477124 241836 477188
rect 241900 477124 241901 477188
rect 241835 477123 241901 477124
rect 239627 476916 239693 476917
rect 239627 476852 239628 476916
rect 239692 476852 239693 476916
rect 239627 476851 239693 476852
rect 240547 476916 240613 476917
rect 240547 476852 240548 476916
rect 240612 476852 240613 476916
rect 240547 476851 240613 476852
rect 243126 476237 243186 479710
rect 244230 476373 244290 479710
rect 244227 476372 244293 476373
rect 244227 476308 244228 476372
rect 244292 476308 244293 476372
rect 244227 476307 244293 476308
rect 245518 476237 245578 479710
rect 246622 476237 246682 479710
rect 247726 476373 247786 479710
rect 248278 479710 248356 479770
rect 248646 479710 248764 479770
rect 250064 479770 250124 480080
rect 250744 479770 250804 480080
rect 251288 479770 251348 480080
rect 252376 479770 252436 480080
rect 253464 479770 253524 480080
rect 250064 479710 250178 479770
rect 250744 479710 250914 479770
rect 251288 479710 251466 479770
rect 247723 476372 247789 476373
rect 247723 476308 247724 476372
rect 247788 476308 247789 476372
rect 247723 476307 247789 476308
rect 248278 476237 248338 479710
rect 248646 476237 248706 479710
rect 250118 476373 250178 479710
rect 250115 476372 250181 476373
rect 250115 476308 250116 476372
rect 250180 476308 250181 476372
rect 250115 476307 250181 476308
rect 250854 476237 250914 479710
rect 251406 476373 251466 479710
rect 252326 479710 252436 479770
rect 253430 479710 253524 479770
rect 253600 479770 253660 480080
rect 254552 479770 254612 480080
rect 255912 479770 255972 480080
rect 253600 479710 253674 479770
rect 251403 476372 251469 476373
rect 251403 476308 251404 476372
rect 251468 476308 251469 476372
rect 251403 476307 251469 476308
rect 252326 476237 252386 479710
rect 253430 477189 253490 479710
rect 253427 477188 253493 477189
rect 253427 477124 253428 477188
rect 253492 477124 253493 477188
rect 253427 477123 253493 477124
rect 253614 476237 253674 479710
rect 254534 479710 254612 479770
rect 255822 479710 255972 479770
rect 256048 479770 256108 480080
rect 257000 479770 257060 480080
rect 258088 479770 258148 480080
rect 256048 479710 256250 479770
rect 257000 479710 257170 479770
rect 254534 476237 254594 479710
rect 255822 476237 255882 479710
rect 256190 477053 256250 479710
rect 256187 477052 256253 477053
rect 256187 476988 256188 477052
rect 256252 476988 256253 477052
rect 256187 476987 256253 476988
rect 257110 476237 257170 479710
rect 257846 479710 258148 479770
rect 258496 479770 258556 480080
rect 259448 479770 259508 480080
rect 260672 479770 260732 480080
rect 258496 479710 258642 479770
rect 259448 479710 259562 479770
rect 257846 476778 257906 479710
rect 258027 476780 258093 476781
rect 258027 476778 258028 476780
rect 257846 476718 258028 476778
rect 258027 476716 258028 476718
rect 258092 476716 258093 476780
rect 258027 476715 258093 476716
rect 258582 476237 258642 479710
rect 259502 476373 259562 479710
rect 260606 479710 260732 479770
rect 261080 479770 261140 480080
rect 261760 479770 261820 480080
rect 262848 479770 262908 480080
rect 261080 479710 261218 479770
rect 259499 476372 259565 476373
rect 259499 476308 259500 476372
rect 259564 476308 259565 476372
rect 259499 476307 259565 476308
rect 260606 476237 260666 479710
rect 261158 476509 261218 479710
rect 261710 479710 261820 479770
rect 262814 479710 262908 479770
rect 263528 479770 263588 480080
rect 263936 479770 263996 480080
rect 263528 479710 263610 479770
rect 261155 476508 261221 476509
rect 261155 476444 261156 476508
rect 261220 476444 261221 476508
rect 261155 476443 261221 476444
rect 261710 476237 261770 479710
rect 262814 476237 262874 479710
rect 263550 476373 263610 479710
rect 263918 479710 263996 479770
rect 265296 479770 265356 480080
rect 265976 479770 266036 480080
rect 265296 479710 265450 479770
rect 263547 476372 263613 476373
rect 263547 476308 263548 476372
rect 263612 476308 263613 476372
rect 263547 476307 263613 476308
rect 263918 476237 263978 479710
rect 265390 476237 265450 479710
rect 265942 479710 266036 479770
rect 266384 479770 266444 480080
rect 267608 479770 267668 480080
rect 266384 479710 266554 479770
rect 265942 476645 266002 479710
rect 265939 476644 266005 476645
rect 265939 476580 265940 476644
rect 266004 476580 266005 476644
rect 265939 476579 266005 476580
rect 266494 476373 266554 479710
rect 267598 479710 267668 479770
rect 268288 479770 268348 480080
rect 268696 479770 268756 480080
rect 269784 479770 269844 480080
rect 271008 479770 271068 480080
rect 268288 479710 268394 479770
rect 268696 479710 268762 479770
rect 269784 479710 269866 479770
rect 266491 476372 266557 476373
rect 266491 476308 266492 476372
rect 266556 476308 266557 476372
rect 266491 476307 266557 476308
rect 267598 476237 267658 479710
rect 268334 476373 268394 479710
rect 268331 476372 268397 476373
rect 268331 476308 268332 476372
rect 268396 476308 268397 476372
rect 268331 476307 268397 476308
rect 268702 476237 268762 479710
rect 269806 476237 269866 479710
rect 270910 479710 271068 479770
rect 271144 479770 271204 480080
rect 272232 479770 272292 480080
rect 273320 479770 273380 480080
rect 271144 479710 271338 479770
rect 270910 476645 270970 479710
rect 270907 476644 270973 476645
rect 270907 476580 270908 476644
rect 270972 476580 270973 476644
rect 270907 476579 270973 476580
rect 271278 476237 271338 479710
rect 272198 479710 272292 479770
rect 273302 479710 273380 479770
rect 273592 479770 273652 480080
rect 274408 479770 274468 480080
rect 273592 479710 273730 479770
rect 272198 476237 272258 479710
rect 273302 476373 273362 479710
rect 273670 476509 273730 479710
rect 274406 479710 274468 479770
rect 275768 479770 275828 480080
rect 276040 479770 276100 480080
rect 276992 479770 277052 480080
rect 275768 479710 275938 479770
rect 276040 479710 276122 479770
rect 273667 476508 273733 476509
rect 273667 476444 273668 476508
rect 273732 476444 273733 476508
rect 273667 476443 273733 476444
rect 273299 476372 273365 476373
rect 273299 476308 273300 476372
rect 273364 476308 273365 476372
rect 273299 476307 273365 476308
rect 274406 476237 274466 479710
rect 275878 476237 275938 479710
rect 276062 476373 276122 479710
rect 276982 479710 277052 479770
rect 278080 479770 278140 480080
rect 278488 479770 278548 480080
rect 278080 479710 278146 479770
rect 276059 476372 276125 476373
rect 276059 476308 276060 476372
rect 276124 476308 276125 476372
rect 276059 476307 276125 476308
rect 276982 476237 277042 479710
rect 278086 476373 278146 479710
rect 278454 479710 278548 479770
rect 279168 479770 279228 480080
rect 280936 479770 280996 480080
rect 283520 479770 283580 480080
rect 285968 479770 286028 480080
rect 288280 479770 288340 480080
rect 291000 479770 291060 480080
rect 279168 479710 279250 479770
rect 280936 479710 281090 479770
rect 283520 479710 283666 479770
rect 285968 479710 286058 479770
rect 278083 476372 278149 476373
rect 278083 476308 278084 476372
rect 278148 476308 278149 476372
rect 278083 476307 278149 476308
rect 278454 476237 278514 479710
rect 279190 476237 279250 479710
rect 281030 476237 281090 479710
rect 283606 476237 283666 479710
rect 285998 476237 286058 479710
rect 288206 479710 288340 479770
rect 290966 479710 291060 479770
rect 293448 479770 293508 480080
rect 295896 479770 295956 480080
rect 298480 479770 298540 480080
rect 300928 479770 300988 480080
rect 303512 479770 303572 480080
rect 293448 479710 293602 479770
rect 295896 479710 295994 479770
rect 298480 479710 298570 479770
rect 288206 476237 288266 479710
rect 290966 476237 291026 479710
rect 293542 476237 293602 479710
rect 295934 476237 295994 479710
rect 298510 476237 298570 479710
rect 300902 479710 300988 479770
rect 303478 479710 303572 479770
rect 305960 479770 306020 480080
rect 308544 479770 308604 480080
rect 310992 479770 311052 480080
rect 313440 479770 313500 480080
rect 315888 479770 315948 480080
rect 305960 479710 306114 479770
rect 308544 479710 308690 479770
rect 310992 479710 311082 479770
rect 300902 476237 300962 479710
rect 303478 476237 303538 479710
rect 306054 476237 306114 479710
rect 308630 476781 308690 479710
rect 308627 476780 308693 476781
rect 308627 476716 308628 476780
rect 308692 476716 308693 476780
rect 308627 476715 308693 476716
rect 311022 476373 311082 479710
rect 313414 479710 313500 479770
rect 315806 479710 315948 479770
rect 318472 479770 318532 480080
rect 320920 479770 320980 480080
rect 323368 479770 323428 480080
rect 325952 479770 326012 480080
rect 318472 479710 318626 479770
rect 320920 479710 321018 479770
rect 313414 476781 313474 479710
rect 313411 476780 313477 476781
rect 313411 476716 313412 476780
rect 313476 476716 313477 476780
rect 313411 476715 313477 476716
rect 311019 476372 311085 476373
rect 311019 476308 311020 476372
rect 311084 476308 311085 476372
rect 311019 476307 311085 476308
rect 315806 476237 315866 479710
rect 318566 476509 318626 479710
rect 320958 477053 321018 479710
rect 323350 479710 323428 479770
rect 325926 479710 326012 479770
rect 320955 477052 321021 477053
rect 320955 476988 320956 477052
rect 321020 476988 321021 477052
rect 320955 476987 321021 476988
rect 323350 476509 323410 479710
rect 325926 476509 325986 479710
rect 318563 476508 318629 476509
rect 318563 476444 318564 476508
rect 318628 476444 318629 476508
rect 318563 476443 318629 476444
rect 323347 476508 323413 476509
rect 323347 476444 323348 476508
rect 323412 476444 323413 476508
rect 323347 476443 323413 476444
rect 325923 476508 325989 476509
rect 325923 476444 325924 476508
rect 325988 476444 325989 476508
rect 325923 476443 325989 476444
rect 237235 476236 237301 476237
rect 237235 476172 237236 476236
rect 237300 476172 237301 476236
rect 237235 476171 237301 476172
rect 243123 476236 243189 476237
rect 243123 476172 243124 476236
rect 243188 476172 243189 476236
rect 243123 476171 243189 476172
rect 245515 476236 245581 476237
rect 245515 476172 245516 476236
rect 245580 476172 245581 476236
rect 245515 476171 245581 476172
rect 246619 476236 246685 476237
rect 246619 476172 246620 476236
rect 246684 476172 246685 476236
rect 246619 476171 246685 476172
rect 248275 476236 248341 476237
rect 248275 476172 248276 476236
rect 248340 476172 248341 476236
rect 248275 476171 248341 476172
rect 248643 476236 248709 476237
rect 248643 476172 248644 476236
rect 248708 476172 248709 476236
rect 248643 476171 248709 476172
rect 250851 476236 250917 476237
rect 250851 476172 250852 476236
rect 250916 476172 250917 476236
rect 250851 476171 250917 476172
rect 252323 476236 252389 476237
rect 252323 476172 252324 476236
rect 252388 476172 252389 476236
rect 252323 476171 252389 476172
rect 253611 476236 253677 476237
rect 253611 476172 253612 476236
rect 253676 476172 253677 476236
rect 253611 476171 253677 476172
rect 254531 476236 254597 476237
rect 254531 476172 254532 476236
rect 254596 476172 254597 476236
rect 254531 476171 254597 476172
rect 255819 476236 255885 476237
rect 255819 476172 255820 476236
rect 255884 476172 255885 476236
rect 255819 476171 255885 476172
rect 257107 476236 257173 476237
rect 257107 476172 257108 476236
rect 257172 476172 257173 476236
rect 257107 476171 257173 476172
rect 258579 476236 258645 476237
rect 258579 476172 258580 476236
rect 258644 476172 258645 476236
rect 258579 476171 258645 476172
rect 260603 476236 260669 476237
rect 260603 476172 260604 476236
rect 260668 476172 260669 476236
rect 260603 476171 260669 476172
rect 261707 476236 261773 476237
rect 261707 476172 261708 476236
rect 261772 476172 261773 476236
rect 261707 476171 261773 476172
rect 262811 476236 262877 476237
rect 262811 476172 262812 476236
rect 262876 476172 262877 476236
rect 262811 476171 262877 476172
rect 263915 476236 263981 476237
rect 263915 476172 263916 476236
rect 263980 476172 263981 476236
rect 263915 476171 263981 476172
rect 265387 476236 265453 476237
rect 265387 476172 265388 476236
rect 265452 476172 265453 476236
rect 265387 476171 265453 476172
rect 267595 476236 267661 476237
rect 267595 476172 267596 476236
rect 267660 476172 267661 476236
rect 267595 476171 267661 476172
rect 268699 476236 268765 476237
rect 268699 476172 268700 476236
rect 268764 476172 268765 476236
rect 268699 476171 268765 476172
rect 269803 476236 269869 476237
rect 269803 476172 269804 476236
rect 269868 476172 269869 476236
rect 269803 476171 269869 476172
rect 271275 476236 271341 476237
rect 271275 476172 271276 476236
rect 271340 476172 271341 476236
rect 271275 476171 271341 476172
rect 272195 476236 272261 476237
rect 272195 476172 272196 476236
rect 272260 476172 272261 476236
rect 272195 476171 272261 476172
rect 274403 476236 274469 476237
rect 274403 476172 274404 476236
rect 274468 476172 274469 476236
rect 274403 476171 274469 476172
rect 275875 476236 275941 476237
rect 275875 476172 275876 476236
rect 275940 476172 275941 476236
rect 275875 476171 275941 476172
rect 276979 476236 277045 476237
rect 276979 476172 276980 476236
rect 277044 476172 277045 476236
rect 276979 476171 277045 476172
rect 278451 476236 278517 476237
rect 278451 476172 278452 476236
rect 278516 476172 278517 476236
rect 278451 476171 278517 476172
rect 279187 476236 279253 476237
rect 279187 476172 279188 476236
rect 279252 476172 279253 476236
rect 279187 476171 279253 476172
rect 281027 476236 281093 476237
rect 281027 476172 281028 476236
rect 281092 476172 281093 476236
rect 281027 476171 281093 476172
rect 283603 476236 283669 476237
rect 283603 476172 283604 476236
rect 283668 476172 283669 476236
rect 283603 476171 283669 476172
rect 285995 476236 286061 476237
rect 285995 476172 285996 476236
rect 286060 476172 286061 476236
rect 285995 476171 286061 476172
rect 288203 476236 288269 476237
rect 288203 476172 288204 476236
rect 288268 476172 288269 476236
rect 288203 476171 288269 476172
rect 290963 476236 291029 476237
rect 290963 476172 290964 476236
rect 291028 476172 291029 476236
rect 290963 476171 291029 476172
rect 293539 476236 293605 476237
rect 293539 476172 293540 476236
rect 293604 476172 293605 476236
rect 293539 476171 293605 476172
rect 295931 476236 295997 476237
rect 295931 476172 295932 476236
rect 295996 476172 295997 476236
rect 295931 476171 295997 476172
rect 298507 476236 298573 476237
rect 298507 476172 298508 476236
rect 298572 476172 298573 476236
rect 298507 476171 298573 476172
rect 300899 476236 300965 476237
rect 300899 476172 300900 476236
rect 300964 476172 300965 476236
rect 300899 476171 300965 476172
rect 303475 476236 303541 476237
rect 303475 476172 303476 476236
rect 303540 476172 303541 476236
rect 303475 476171 303541 476172
rect 306051 476236 306117 476237
rect 306051 476172 306052 476236
rect 306116 476172 306117 476236
rect 306051 476171 306117 476172
rect 315803 476236 315869 476237
rect 315803 476172 315804 476236
rect 315868 476172 315869 476236
rect 315803 476171 315869 476172
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 443544 362414 470898
rect 366294 706108 366914 711900
rect 366294 705872 366326 706108
rect 366562 705872 366646 706108
rect 366882 705872 366914 706108
rect 366294 705788 366914 705872
rect 366294 705552 366326 705788
rect 366562 705552 366646 705788
rect 366882 705552 366914 705788
rect 366294 691954 366914 705552
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 364931 444684 364997 444685
rect 364931 444620 364932 444684
rect 364996 444620 364997 444684
rect 364931 444619 364997 444620
rect 362539 443324 362605 443325
rect 362539 443260 362540 443324
rect 362604 443260 362605 443324
rect 362539 443259 362605 443260
rect 236608 435454 236928 435486
rect 236608 435218 236650 435454
rect 236886 435218 236928 435454
rect 236608 435134 236928 435218
rect 236608 434898 236650 435134
rect 236886 434898 236928 435134
rect 236608 434866 236928 434898
rect 267328 435454 267648 435486
rect 267328 435218 267370 435454
rect 267606 435218 267648 435454
rect 267328 435134 267648 435218
rect 267328 434898 267370 435134
rect 267606 434898 267648 435134
rect 267328 434866 267648 434898
rect 298048 435454 298368 435486
rect 298048 435218 298090 435454
rect 298326 435218 298368 435454
rect 298048 435134 298368 435218
rect 298048 434898 298090 435134
rect 298326 434898 298368 435134
rect 298048 434866 298368 434898
rect 328768 435454 329088 435486
rect 328768 435218 328810 435454
rect 329046 435218 329088 435454
rect 328768 435134 329088 435218
rect 328768 434898 328810 435134
rect 329046 434898 329088 435134
rect 328768 434866 329088 434898
rect 359488 435454 359808 435486
rect 359488 435218 359530 435454
rect 359766 435218 359808 435454
rect 359488 435134 359808 435218
rect 359488 434898 359530 435134
rect 359766 434898 359808 435134
rect 359488 434866 359808 434898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 251968 403954 252288 403986
rect 251968 403718 252010 403954
rect 252246 403718 252288 403954
rect 251968 403634 252288 403718
rect 251968 403398 252010 403634
rect 252246 403398 252288 403634
rect 251968 403366 252288 403398
rect 282688 403954 283008 403986
rect 282688 403718 282730 403954
rect 282966 403718 283008 403954
rect 282688 403634 283008 403718
rect 282688 403398 282730 403634
rect 282966 403398 283008 403634
rect 282688 403366 283008 403398
rect 313408 403954 313728 403986
rect 313408 403718 313450 403954
rect 313686 403718 313728 403954
rect 313408 403634 313728 403718
rect 313408 403398 313450 403634
rect 313686 403398 313728 403634
rect 313408 403366 313728 403398
rect 344128 403954 344448 403986
rect 344128 403718 344170 403954
rect 344406 403718 344448 403954
rect 344128 403634 344448 403718
rect 344128 403398 344170 403634
rect 344406 403398 344448 403634
rect 344128 403366 344448 403398
rect 236608 399454 236928 399486
rect 236608 399218 236650 399454
rect 236886 399218 236928 399454
rect 236608 399134 236928 399218
rect 236608 398898 236650 399134
rect 236886 398898 236928 399134
rect 236608 398866 236928 398898
rect 267328 399454 267648 399486
rect 267328 399218 267370 399454
rect 267606 399218 267648 399454
rect 267328 399134 267648 399218
rect 267328 398898 267370 399134
rect 267606 398898 267648 399134
rect 267328 398866 267648 398898
rect 298048 399454 298368 399486
rect 298048 399218 298090 399454
rect 298326 399218 298368 399454
rect 298048 399134 298368 399218
rect 298048 398898 298090 399134
rect 298326 398898 298368 399134
rect 298048 398866 298368 398898
rect 328768 399454 329088 399486
rect 328768 399218 328810 399454
rect 329046 399218 329088 399454
rect 328768 399134 329088 399218
rect 328768 398898 328810 399134
rect 329046 398898 329088 399134
rect 328768 398866 329088 398898
rect 359488 399454 359808 399486
rect 359488 399218 359530 399454
rect 359766 399218 359808 399454
rect 359488 399134 359808 399218
rect 359488 398898 359530 399134
rect 359766 398898 359808 399134
rect 359488 398866 359808 398898
rect 232083 374100 232149 374101
rect 232083 374036 232084 374100
rect 232148 374036 232149 374100
rect 232083 374035 232149 374036
rect 231899 373284 231965 373285
rect 231899 373220 231900 373284
rect 231964 373220 231965 373284
rect 231899 373219 231965 373220
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 231902 310317 231962 373219
rect 232086 364350 232146 374035
rect 251968 367954 252288 367986
rect 251968 367718 252010 367954
rect 252246 367718 252288 367954
rect 251968 367634 252288 367718
rect 251968 367398 252010 367634
rect 252246 367398 252288 367634
rect 251968 367366 252288 367398
rect 282688 367954 283008 367986
rect 282688 367718 282730 367954
rect 282966 367718 283008 367954
rect 282688 367634 283008 367718
rect 282688 367398 282730 367634
rect 282966 367398 283008 367634
rect 282688 367366 283008 367398
rect 313408 367954 313728 367986
rect 313408 367718 313450 367954
rect 313686 367718 313728 367954
rect 313408 367634 313728 367718
rect 313408 367398 313450 367634
rect 313686 367398 313728 367634
rect 313408 367366 313728 367398
rect 344128 367954 344448 367986
rect 344128 367718 344170 367954
rect 344406 367718 344448 367954
rect 344128 367634 344448 367718
rect 344128 367398 344170 367634
rect 344406 367398 344448 367634
rect 344128 367366 344448 367398
rect 232086 364290 232514 364350
rect 232083 311268 232149 311269
rect 232083 311204 232084 311268
rect 232148 311204 232149 311268
rect 232083 311203 232149 311204
rect 232086 310453 232146 311203
rect 232083 310452 232149 310453
rect 232083 310388 232084 310452
rect 232148 310388 232149 310452
rect 232083 310387 232149 310388
rect 231899 310316 231965 310317
rect 231899 310252 231900 310316
rect 231964 310252 231965 310316
rect 231899 310251 231965 310252
rect 232454 309773 232514 364290
rect 236608 363454 236928 363486
rect 236608 363218 236650 363454
rect 236886 363218 236928 363454
rect 236608 363134 236928 363218
rect 236608 362898 236650 363134
rect 236886 362898 236928 363134
rect 236608 362866 236928 362898
rect 267328 363454 267648 363486
rect 267328 363218 267370 363454
rect 267606 363218 267648 363454
rect 267328 363134 267648 363218
rect 267328 362898 267370 363134
rect 267606 362898 267648 363134
rect 267328 362866 267648 362898
rect 298048 363454 298368 363486
rect 298048 363218 298090 363454
rect 298326 363218 298368 363454
rect 298048 363134 298368 363218
rect 298048 362898 298090 363134
rect 298326 362898 298368 363134
rect 298048 362866 298368 362898
rect 328768 363454 329088 363486
rect 328768 363218 328810 363454
rect 329046 363218 329088 363454
rect 328768 363134 329088 363218
rect 328768 362898 328810 363134
rect 329046 362898 329088 363134
rect 328768 362866 329088 362898
rect 359488 363454 359808 363486
rect 359488 363218 359530 363454
rect 359766 363218 359808 363454
rect 359488 363134 359808 363218
rect 359488 362898 359530 363134
rect 359766 362898 359808 363134
rect 359488 362866 359808 362898
rect 251968 331954 252288 331986
rect 251968 331718 252010 331954
rect 252246 331718 252288 331954
rect 251968 331634 252288 331718
rect 251968 331398 252010 331634
rect 252246 331398 252288 331634
rect 251968 331366 252288 331398
rect 282688 331954 283008 331986
rect 282688 331718 282730 331954
rect 282966 331718 283008 331954
rect 282688 331634 283008 331718
rect 282688 331398 282730 331634
rect 282966 331398 283008 331634
rect 282688 331366 283008 331398
rect 313408 331954 313728 331986
rect 313408 331718 313450 331954
rect 313686 331718 313728 331954
rect 313408 331634 313728 331718
rect 313408 331398 313450 331634
rect 313686 331398 313728 331634
rect 313408 331366 313728 331398
rect 344128 331954 344448 331986
rect 344128 331718 344170 331954
rect 344406 331718 344448 331954
rect 344128 331634 344448 331718
rect 344128 331398 344170 331634
rect 344406 331398 344448 331634
rect 344128 331366 344448 331398
rect 236608 327454 236928 327486
rect 236608 327218 236650 327454
rect 236886 327218 236928 327454
rect 236608 327134 236928 327218
rect 236608 326898 236650 327134
rect 236886 326898 236928 327134
rect 236608 326866 236928 326898
rect 267328 327454 267648 327486
rect 267328 327218 267370 327454
rect 267606 327218 267648 327454
rect 267328 327134 267648 327218
rect 267328 326898 267370 327134
rect 267606 326898 267648 327134
rect 267328 326866 267648 326898
rect 298048 327454 298368 327486
rect 298048 327218 298090 327454
rect 298326 327218 298368 327454
rect 298048 327134 298368 327218
rect 298048 326898 298090 327134
rect 298326 326898 298368 327134
rect 298048 326866 298368 326898
rect 328768 327454 329088 327486
rect 328768 327218 328810 327454
rect 329046 327218 329088 327454
rect 328768 327134 329088 327218
rect 328768 326898 328810 327134
rect 329046 326898 329088 327134
rect 328768 326866 329088 326898
rect 359488 327454 359808 327486
rect 359488 327218 359530 327454
rect 359766 327218 359808 327454
rect 359488 327134 359808 327218
rect 359488 326898 359530 327134
rect 359766 326898 359808 327134
rect 359488 326866 359808 326898
rect 232451 309772 232517 309773
rect 232451 309708 232452 309772
rect 232516 309708 232517 309772
rect 232451 309707 232517 309708
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 245308 227414 263898
rect 231294 304954 231914 308400
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 245308 231914 268398
rect 244794 282454 245414 308400
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 246454 245414 281898
rect 244794 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 245414 246454
rect 244794 246134 245414 246218
rect 244794 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 245414 246134
rect 244794 245308 245414 245898
rect 249294 286954 249914 308400
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 245308 249914 250398
rect 253794 291454 254414 308400
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 245308 254414 254898
rect 258294 295954 258914 308400
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 245308 258914 259398
rect 262794 300454 263414 308400
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 245308 263414 263898
rect 267294 304954 267914 308400
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 245308 267914 268398
rect 280794 282454 281414 308400
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 246454 281414 281898
rect 280794 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 281414 246454
rect 280794 246134 281414 246218
rect 280794 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 281414 246134
rect 280794 245308 281414 245898
rect 285294 286954 285914 308400
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 245308 285914 250398
rect 289794 291454 290414 308400
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 245308 290414 254898
rect 294294 295954 294914 308400
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 245308 294914 259398
rect 298794 300454 299414 308400
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 245308 299414 263898
rect 303294 304954 303914 308400
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 245308 303914 268398
rect 316794 282454 317414 308400
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 246454 317414 281898
rect 316794 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 317414 246454
rect 316794 246134 317414 246218
rect 316794 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 317414 246134
rect 316794 245308 317414 245898
rect 321294 286954 321914 308400
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 245308 321914 250398
rect 325794 291454 326414 308400
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 245308 326414 254898
rect 330294 295954 330914 308400
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 245308 330914 259398
rect 334794 300454 335414 308400
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 245308 335414 263898
rect 339294 304954 339914 308400
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 245308 339914 268398
rect 352794 282454 353414 308400
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 245308 353414 245898
rect 357294 286954 357914 308400
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 361794 291454 362414 308400
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 358859 251972 358925 251973
rect 358859 251908 358860 251972
rect 358924 251908 358925 251972
rect 358859 251907 358925 251908
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 358123 250884 358189 250885
rect 358123 250820 358124 250884
rect 358188 250820 358189 250884
rect 358123 250819 358189 250820
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 245308 357914 250398
rect 220272 223954 220620 223986
rect 220272 223718 220328 223954
rect 220564 223718 220620 223954
rect 220272 223634 220620 223718
rect 220272 223398 220328 223634
rect 220564 223398 220620 223634
rect 220272 223366 220620 223398
rect 356000 223954 356348 223986
rect 356000 223718 356056 223954
rect 356292 223718 356348 223954
rect 356000 223634 356348 223718
rect 356000 223398 356056 223634
rect 356292 223398 356348 223634
rect 356000 223366 356348 223398
rect 220952 219454 221300 219486
rect 220952 219218 221008 219454
rect 221244 219218 221300 219454
rect 220952 219134 221300 219218
rect 220952 218898 221008 219134
rect 221244 218898 221300 219134
rect 220952 218866 221300 218898
rect 355320 219454 355668 219486
rect 355320 219218 355376 219454
rect 355612 219218 355668 219454
rect 355320 219134 355668 219218
rect 355320 218898 355376 219134
rect 355612 218898 355668 219134
rect 355320 218866 355668 218898
rect 220272 187954 220620 187986
rect 220272 187718 220328 187954
rect 220564 187718 220620 187954
rect 220272 187634 220620 187718
rect 220272 187398 220328 187634
rect 220564 187398 220620 187634
rect 220272 187366 220620 187398
rect 356000 187954 356348 187986
rect 356000 187718 356056 187954
rect 356292 187718 356348 187954
rect 356000 187634 356348 187718
rect 356000 187398 356056 187634
rect 356292 187398 356348 187634
rect 356000 187366 356348 187398
rect 220952 183454 221300 183486
rect 220952 183218 221008 183454
rect 221244 183218 221300 183454
rect 220952 183134 221300 183218
rect 220952 182898 221008 183134
rect 221244 182898 221300 183134
rect 220952 182866 221300 182898
rect 355320 183454 355668 183486
rect 355320 183218 355376 183454
rect 355612 183218 355668 183454
rect 355320 183134 355668 183218
rect 355320 182898 355376 183134
rect 355612 182898 355668 183134
rect 355320 182866 355668 182898
rect 236056 159490 236116 160106
rect 237144 159490 237204 160106
rect 238232 159490 238292 160106
rect 236056 159430 236194 159490
rect 237144 159430 237298 159490
rect 236134 158813 236194 159430
rect 236131 158812 236197 158813
rect 236131 158748 236132 158812
rect 236196 158748 236197 158812
rect 236131 158747 236197 158748
rect 219203 158404 219269 158405
rect 219203 158340 219204 158404
rect 219268 158340 219269 158404
rect 219203 158339 219269 158340
rect 222294 151954 222914 158000
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 214419 3364 214485 3365
rect 214419 3300 214420 3364
rect 214484 3300 214485 3364
rect 214419 3299 214485 3300
rect 213294 -7612 213326 -7376
rect 213562 -7612 213646 -7376
rect 213882 -7612 213914 -7376
rect 213294 -7696 213914 -7612
rect 213294 -7932 213326 -7696
rect 213562 -7932 213646 -7696
rect 213882 -7932 213914 -7696
rect 213294 -7964 213914 -7932
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 218651 3500 218717 3501
rect 218651 3436 218652 3500
rect 218716 3436 218717 3500
rect 218651 3435 218717 3436
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -656 218414 2898
rect 217794 -892 217826 -656
rect 218062 -892 218146 -656
rect 218382 -892 218414 -656
rect 217794 -976 218414 -892
rect 217794 -1212 217826 -976
rect 218062 -1212 218146 -976
rect 218382 -1212 218414 -976
rect 217794 -7964 218414 -1212
rect 222294 -1616 222914 7398
rect 222294 -1852 222326 -1616
rect 222562 -1852 222646 -1616
rect 222882 -1852 222914 -1616
rect 222294 -1936 222914 -1852
rect 222294 -2172 222326 -1936
rect 222562 -2172 222646 -1936
rect 222882 -2172 222914 -1936
rect 222294 -7964 222914 -2172
rect 226794 156454 227414 158000
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2576 227414 11898
rect 226794 -2812 226826 -2576
rect 227062 -2812 227146 -2576
rect 227382 -2812 227414 -2576
rect 226794 -2896 227414 -2812
rect 226794 -3132 226826 -2896
rect 227062 -3132 227146 -2896
rect 227382 -3132 227414 -2896
rect 226794 -7964 227414 -3132
rect 231294 124954 231914 158000
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3536 231914 16398
rect 231294 -3772 231326 -3536
rect 231562 -3772 231646 -3536
rect 231882 -3772 231914 -3536
rect 231294 -3856 231914 -3772
rect 231294 -4092 231326 -3856
rect 231562 -4092 231646 -3856
rect 231882 -4092 231914 -3856
rect 231294 -7964 231914 -4092
rect 235794 129454 236414 158000
rect 237238 157861 237298 159430
rect 238158 159430 238292 159490
rect 239592 159490 239652 160106
rect 240544 159490 240604 160106
rect 241768 159490 241828 160106
rect 243128 159490 243188 160106
rect 239592 159430 239690 159490
rect 240544 159430 240610 159490
rect 241768 159430 241898 159490
rect 238158 158677 238218 159430
rect 239630 158677 239690 159430
rect 240550 158677 240610 159430
rect 238155 158676 238221 158677
rect 238155 158612 238156 158676
rect 238220 158612 238221 158676
rect 238155 158611 238221 158612
rect 239627 158676 239693 158677
rect 239627 158612 239628 158676
rect 239692 158612 239693 158676
rect 239627 158611 239693 158612
rect 240547 158676 240613 158677
rect 240547 158612 240548 158676
rect 240612 158612 240613 158676
rect 240547 158611 240613 158612
rect 237235 157860 237301 157861
rect 237235 157796 237236 157860
rect 237300 157796 237301 157860
rect 237235 157795 237301 157796
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4496 236414 20898
rect 235794 -4732 235826 -4496
rect 236062 -4732 236146 -4496
rect 236382 -4732 236414 -4496
rect 235794 -4816 236414 -4732
rect 235794 -5052 235826 -4816
rect 236062 -5052 236146 -4816
rect 236382 -5052 236414 -4816
rect 235794 -7964 236414 -5052
rect 240294 133954 240914 158000
rect 241838 157453 241898 159430
rect 243126 159430 243188 159490
rect 244216 159490 244276 160106
rect 245440 159490 245500 160106
rect 246528 159490 246588 160106
rect 247616 159490 247676 160106
rect 248296 159490 248356 160106
rect 248704 159490 248764 160106
rect 244216 159430 244290 159490
rect 245440 159430 245578 159490
rect 246528 159430 246682 159490
rect 247616 159430 247786 159490
rect 243126 158949 243186 159430
rect 243123 158948 243189 158949
rect 243123 158884 243124 158948
rect 243188 158884 243189 158948
rect 243123 158883 243189 158884
rect 244230 158269 244290 159430
rect 244227 158268 244293 158269
rect 244227 158204 244228 158268
rect 244292 158204 244293 158268
rect 244227 158203 244293 158204
rect 241835 157452 241901 157453
rect 241835 157388 241836 157452
rect 241900 157388 241901 157452
rect 241835 157387 241901 157388
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5456 240914 25398
rect 240294 -5692 240326 -5456
rect 240562 -5692 240646 -5456
rect 240882 -5692 240914 -5456
rect 240294 -5776 240914 -5692
rect 240294 -6012 240326 -5776
rect 240562 -6012 240646 -5776
rect 240882 -6012 240914 -5776
rect 240294 -7964 240914 -6012
rect 244794 138454 245414 158000
rect 245518 157453 245578 159430
rect 246622 158133 246682 159430
rect 246619 158132 246685 158133
rect 246619 158068 246620 158132
rect 246684 158068 246685 158132
rect 246619 158067 246685 158068
rect 245515 157452 245581 157453
rect 245515 157388 245516 157452
rect 245580 157388 245581 157452
rect 245515 157387 245581 157388
rect 247726 157045 247786 159430
rect 248278 159430 248356 159490
rect 248646 159430 248764 159490
rect 250064 159490 250124 160106
rect 250744 159490 250804 160106
rect 251288 159490 251348 160106
rect 252376 159490 252436 160106
rect 253464 159490 253524 160106
rect 250064 159430 250178 159490
rect 250744 159430 250914 159490
rect 251288 159430 251466 159490
rect 248278 158677 248338 159430
rect 248275 158676 248341 158677
rect 248275 158612 248276 158676
rect 248340 158612 248341 158676
rect 248275 158611 248341 158612
rect 248646 157997 248706 159430
rect 250118 158677 250178 159430
rect 250854 159085 250914 159430
rect 250851 159084 250917 159085
rect 250851 159020 250852 159084
rect 250916 159020 250917 159084
rect 250851 159019 250917 159020
rect 250115 158676 250181 158677
rect 250115 158612 250116 158676
rect 250180 158612 250181 158676
rect 250115 158611 250181 158612
rect 248643 157996 248709 157997
rect 248643 157932 248644 157996
rect 248708 157932 248709 157996
rect 248643 157931 248709 157932
rect 247723 157044 247789 157045
rect 247723 156980 247724 157044
rect 247788 156980 247789 157044
rect 247723 156979 247789 156980
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6416 245414 29898
rect 244794 -6652 244826 -6416
rect 245062 -6652 245146 -6416
rect 245382 -6652 245414 -6416
rect 244794 -6736 245414 -6652
rect 244794 -6972 244826 -6736
rect 245062 -6972 245146 -6736
rect 245382 -6972 245414 -6736
rect 244794 -7964 245414 -6972
rect 249294 142954 249914 158000
rect 251406 157997 251466 159430
rect 252326 159430 252436 159490
rect 253430 159430 253524 159490
rect 253600 159490 253660 160106
rect 254552 159490 254612 160106
rect 255912 159629 255972 160106
rect 255909 159628 255975 159629
rect 255909 159564 255910 159628
rect 255974 159564 255975 159628
rect 255909 159563 255975 159564
rect 256048 159490 256108 160106
rect 253600 159430 253674 159490
rect 252326 158541 252386 159430
rect 252323 158540 252389 158541
rect 252323 158476 252324 158540
rect 252388 158476 252389 158540
rect 252323 158475 252389 158476
rect 253430 157997 253490 159430
rect 251403 157996 251469 157997
rect 251403 157932 251404 157996
rect 251468 157932 251469 157996
rect 251403 157931 251469 157932
rect 253427 157996 253493 157997
rect 253427 157932 253428 157996
rect 253492 157932 253493 157996
rect 253427 157931 253493 157932
rect 253614 157453 253674 159430
rect 254534 159430 254612 159490
rect 256006 159430 256108 159490
rect 257000 159490 257060 160106
rect 258088 159490 258148 160106
rect 258496 159901 258556 160106
rect 258493 159900 258559 159901
rect 258493 159836 258494 159900
rect 258558 159836 258559 159900
rect 258493 159835 258559 159836
rect 259448 159490 259508 160106
rect 260672 159490 260732 160106
rect 257000 159430 257170 159490
rect 258088 159430 258274 159490
rect 259448 159430 259562 159490
rect 254534 159221 254594 159430
rect 254531 159220 254597 159221
rect 254531 159156 254532 159220
rect 254596 159156 254597 159220
rect 254531 159155 254597 159156
rect 256006 158677 256066 159430
rect 257110 158677 257170 159430
rect 258214 158677 258274 159430
rect 259502 158677 259562 159430
rect 260606 159430 260732 159490
rect 261080 159490 261140 160106
rect 261760 159490 261820 160106
rect 262848 159490 262908 160106
rect 261080 159430 261218 159490
rect 256003 158676 256069 158677
rect 256003 158612 256004 158676
rect 256068 158612 256069 158676
rect 256003 158611 256069 158612
rect 257107 158676 257173 158677
rect 257107 158612 257108 158676
rect 257172 158612 257173 158676
rect 257107 158611 257173 158612
rect 258211 158676 258277 158677
rect 258211 158612 258212 158676
rect 258276 158612 258277 158676
rect 258211 158611 258277 158612
rect 259499 158676 259565 158677
rect 259499 158612 259500 158676
rect 259564 158612 259565 158676
rect 259499 158611 259565 158612
rect 260606 158541 260666 159430
rect 261158 158677 261218 159430
rect 261710 159430 261820 159490
rect 262814 159430 262908 159490
rect 263528 159490 263588 160106
rect 263936 159490 263996 160106
rect 263528 159430 263610 159490
rect 261155 158676 261221 158677
rect 261155 158612 261156 158676
rect 261220 158612 261221 158676
rect 261155 158611 261221 158612
rect 260603 158540 260669 158541
rect 260603 158476 260604 158540
rect 260668 158476 260669 158540
rect 260603 158475 260669 158476
rect 253611 157452 253677 157453
rect 253611 157388 253612 157452
rect 253676 157388 253677 157452
rect 253611 157387 253677 157388
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7376 249914 34398
rect 249294 -7612 249326 -7376
rect 249562 -7612 249646 -7376
rect 249882 -7612 249914 -7376
rect 249294 -7696 249914 -7612
rect 249294 -7932 249326 -7696
rect 249562 -7932 249646 -7696
rect 249882 -7932 249914 -7696
rect 249294 -7964 249914 -7932
rect 253794 147454 254414 158000
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -656 254414 2898
rect 253794 -892 253826 -656
rect 254062 -892 254146 -656
rect 254382 -892 254414 -656
rect 253794 -976 254414 -892
rect 253794 -1212 253826 -976
rect 254062 -1212 254146 -976
rect 254382 -1212 254414 -976
rect 253794 -7964 254414 -1212
rect 258294 151954 258914 158000
rect 261710 157997 261770 159430
rect 262814 158677 262874 159430
rect 262811 158676 262877 158677
rect 262811 158612 262812 158676
rect 262876 158612 262877 158676
rect 262811 158611 262877 158612
rect 261707 157996 261773 157997
rect 261707 157932 261708 157996
rect 261772 157932 261773 157996
rect 261707 157931 261773 157932
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1616 258914 7398
rect 258294 -1852 258326 -1616
rect 258562 -1852 258646 -1616
rect 258882 -1852 258914 -1616
rect 258294 -1936 258914 -1852
rect 258294 -2172 258326 -1936
rect 258562 -2172 258646 -1936
rect 258882 -2172 258914 -1936
rect 258294 -7964 258914 -2172
rect 262794 156454 263414 158000
rect 263550 157453 263610 159430
rect 263918 159430 263996 159490
rect 265296 159490 265356 160106
rect 265976 159490 266036 160106
rect 265296 159430 265450 159490
rect 263918 157725 263978 159430
rect 265390 157725 265450 159430
rect 265942 159430 266036 159490
rect 266384 159490 266444 160106
rect 267608 159490 267668 160106
rect 266384 159430 266554 159490
rect 265942 158677 266002 159430
rect 265939 158676 266005 158677
rect 265939 158612 265940 158676
rect 266004 158612 266005 158676
rect 265939 158611 266005 158612
rect 266494 157997 266554 159430
rect 267598 159430 267668 159490
rect 268288 159490 268348 160106
rect 268696 159490 268756 160106
rect 269784 159490 269844 160106
rect 271008 159629 271068 160106
rect 271005 159628 271071 159629
rect 271005 159564 271006 159628
rect 271070 159564 271071 159628
rect 271005 159563 271071 159564
rect 271144 159490 271204 160106
rect 272232 159490 272292 160106
rect 273320 159490 273380 160106
rect 268288 159430 268394 159490
rect 268696 159430 268762 159490
rect 269784 159430 269866 159490
rect 267598 158677 267658 159430
rect 267595 158676 267661 158677
rect 267595 158612 267596 158676
rect 267660 158612 267661 158676
rect 267595 158611 267661 158612
rect 266491 157996 266557 157997
rect 266491 157932 266492 157996
rect 266556 157932 266557 157996
rect 266491 157931 266557 157932
rect 263915 157724 263981 157725
rect 263915 157660 263916 157724
rect 263980 157660 263981 157724
rect 263915 157659 263981 157660
rect 265387 157724 265453 157725
rect 265387 157660 265388 157724
rect 265452 157660 265453 157724
rect 265387 157659 265453 157660
rect 263547 157452 263613 157453
rect 263547 157388 263548 157452
rect 263612 157388 263613 157452
rect 263547 157387 263613 157388
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2576 263414 11898
rect 262794 -2812 262826 -2576
rect 263062 -2812 263146 -2576
rect 263382 -2812 263414 -2576
rect 262794 -2896 263414 -2812
rect 262794 -3132 262826 -2896
rect 263062 -3132 263146 -2896
rect 263382 -3132 263414 -2896
rect 262794 -7964 263414 -3132
rect 267294 124954 267914 158000
rect 268334 157997 268394 159430
rect 268702 158677 268762 159430
rect 269806 158677 269866 159430
rect 271094 159430 271204 159490
rect 272198 159430 272292 159490
rect 273302 159430 273380 159490
rect 273592 159490 273652 160106
rect 274408 159629 274468 160106
rect 275768 159901 275828 160106
rect 275765 159900 275831 159901
rect 275765 159836 275766 159900
rect 275830 159836 275831 159900
rect 275765 159835 275831 159836
rect 274405 159628 274471 159629
rect 274405 159564 274406 159628
rect 274470 159564 274471 159628
rect 274405 159563 274471 159564
rect 276040 159490 276100 160106
rect 276992 159901 277052 160106
rect 278080 159901 278140 160106
rect 276989 159900 277055 159901
rect 276989 159836 276990 159900
rect 277054 159836 277055 159900
rect 276989 159835 277055 159836
rect 278077 159900 278143 159901
rect 278077 159836 278078 159900
rect 278142 159836 278143 159900
rect 278488 159898 278548 160106
rect 279168 159901 279228 160106
rect 278077 159835 278143 159836
rect 278454 159838 278548 159898
rect 279165 159900 279231 159901
rect 273592 159430 273730 159490
rect 276040 159430 276122 159490
rect 271094 158677 271154 159430
rect 272198 158677 272258 159430
rect 268699 158676 268765 158677
rect 268699 158612 268700 158676
rect 268764 158612 268765 158676
rect 268699 158611 268765 158612
rect 269803 158676 269869 158677
rect 269803 158612 269804 158676
rect 269868 158612 269869 158676
rect 269803 158611 269869 158612
rect 271091 158676 271157 158677
rect 271091 158612 271092 158676
rect 271156 158612 271157 158676
rect 271091 158611 271157 158612
rect 272195 158676 272261 158677
rect 272195 158612 272196 158676
rect 272260 158612 272261 158676
rect 272195 158611 272261 158612
rect 273302 158405 273362 159430
rect 273299 158404 273365 158405
rect 273299 158340 273300 158404
rect 273364 158340 273365 158404
rect 273299 158339 273365 158340
rect 268331 157996 268397 157997
rect 268331 157932 268332 157996
rect 268396 157932 268397 157996
rect 268331 157931 268397 157932
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3536 267914 16398
rect 267294 -3772 267326 -3536
rect 267562 -3772 267646 -3536
rect 267882 -3772 267914 -3536
rect 267294 -3856 267914 -3772
rect 267294 -4092 267326 -3856
rect 267562 -4092 267646 -3856
rect 267882 -4092 267914 -3856
rect 267294 -7964 267914 -4092
rect 271794 129454 272414 158000
rect 273670 157725 273730 159430
rect 276062 158541 276122 159430
rect 276059 158540 276125 158541
rect 276059 158476 276060 158540
rect 276124 158476 276125 158540
rect 276059 158475 276125 158476
rect 273667 157724 273733 157725
rect 273667 157660 273668 157724
rect 273732 157660 273733 157724
rect 273667 157659 273733 157660
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4496 272414 20898
rect 271794 -4732 271826 -4496
rect 272062 -4732 272146 -4496
rect 272382 -4732 272414 -4496
rect 271794 -4816 272414 -4732
rect 271794 -5052 271826 -4816
rect 272062 -5052 272146 -4816
rect 272382 -5052 272414 -4816
rect 271794 -7964 272414 -5052
rect 276294 133954 276914 158000
rect 278454 157725 278514 159838
rect 279165 159836 279166 159900
rect 279230 159836 279231 159900
rect 279165 159835 279231 159836
rect 280936 159490 280996 160106
rect 283520 159490 283580 160106
rect 285968 159898 286028 160106
rect 285968 159838 286058 159898
rect 280936 159430 281090 159490
rect 283520 159430 283666 159490
rect 281030 158541 281090 159430
rect 281027 158540 281093 158541
rect 281027 158476 281028 158540
rect 281092 158476 281093 158540
rect 281027 158475 281093 158476
rect 278451 157724 278517 157725
rect 278451 157660 278452 157724
rect 278516 157660 278517 157724
rect 278451 157659 278517 157660
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5456 276914 25398
rect 276294 -5692 276326 -5456
rect 276562 -5692 276646 -5456
rect 276882 -5692 276914 -5456
rect 276294 -5776 276914 -5692
rect 276294 -6012 276326 -5776
rect 276562 -6012 276646 -5776
rect 276882 -6012 276914 -5776
rect 276294 -7964 276914 -6012
rect 280794 138454 281414 158000
rect 283606 157725 283666 159430
rect 285998 158541 286058 159838
rect 288280 159490 288340 160106
rect 291000 159490 291060 160106
rect 288206 159430 288340 159490
rect 290966 159430 291060 159490
rect 293448 159490 293508 160106
rect 295896 159490 295956 160106
rect 298480 159490 298540 160106
rect 300928 159765 300988 160106
rect 300925 159764 300991 159765
rect 300925 159700 300926 159764
rect 300990 159700 300991 159764
rect 300925 159699 300991 159700
rect 303512 159490 303572 160106
rect 293448 159430 293602 159490
rect 295896 159430 295994 159490
rect 298480 159430 298570 159490
rect 285995 158540 286061 158541
rect 285995 158476 285996 158540
rect 286060 158476 286061 158540
rect 285995 158475 286061 158476
rect 283603 157724 283669 157725
rect 283603 157660 283604 157724
rect 283668 157660 283669 157724
rect 283603 157659 283669 157660
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6416 281414 29898
rect 280794 -6652 280826 -6416
rect 281062 -6652 281146 -6416
rect 281382 -6652 281414 -6416
rect 280794 -6736 281414 -6652
rect 280794 -6972 280826 -6736
rect 281062 -6972 281146 -6736
rect 281382 -6972 281414 -6736
rect 280794 -7964 281414 -6972
rect 285294 142954 285914 158000
rect 288206 157589 288266 159430
rect 290966 158405 291026 159430
rect 290963 158404 291029 158405
rect 290963 158340 290964 158404
rect 291028 158340 291029 158404
rect 290963 158339 291029 158340
rect 288203 157588 288269 157589
rect 288203 157524 288204 157588
rect 288268 157524 288269 157588
rect 288203 157523 288269 157524
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7376 285914 34398
rect 285294 -7612 285326 -7376
rect 285562 -7612 285646 -7376
rect 285882 -7612 285914 -7376
rect 285294 -7696 285914 -7612
rect 285294 -7932 285326 -7696
rect 285562 -7932 285646 -7696
rect 285882 -7932 285914 -7696
rect 285294 -7964 285914 -7932
rect 289794 147454 290414 158000
rect 293542 157589 293602 159430
rect 295934 158405 295994 159430
rect 298510 158677 298570 159430
rect 303478 159430 303572 159490
rect 305960 159490 306020 160106
rect 308544 159490 308604 160106
rect 310992 159490 311052 160106
rect 313440 159490 313500 160106
rect 315888 159490 315948 160106
rect 305960 159430 306114 159490
rect 308544 159430 308690 159490
rect 310992 159430 311082 159490
rect 303478 158677 303538 159430
rect 306054 158677 306114 159430
rect 308630 158677 308690 159430
rect 298507 158676 298573 158677
rect 298507 158612 298508 158676
rect 298572 158612 298573 158676
rect 298507 158611 298573 158612
rect 303475 158676 303541 158677
rect 303475 158612 303476 158676
rect 303540 158612 303541 158676
rect 303475 158611 303541 158612
rect 306051 158676 306117 158677
rect 306051 158612 306052 158676
rect 306116 158612 306117 158676
rect 306051 158611 306117 158612
rect 308627 158676 308693 158677
rect 308627 158612 308628 158676
rect 308692 158612 308693 158676
rect 308627 158611 308693 158612
rect 295931 158404 295997 158405
rect 295931 158340 295932 158404
rect 295996 158340 295997 158404
rect 295931 158339 295997 158340
rect 311022 158269 311082 159430
rect 313414 159430 313500 159490
rect 315806 159430 315948 159490
rect 318472 159490 318532 160106
rect 320920 159490 320980 160106
rect 323368 159490 323428 160106
rect 325952 159490 326012 160106
rect 318472 159430 318626 159490
rect 320920 159430 321018 159490
rect 313414 158677 313474 159430
rect 315806 158677 315866 159430
rect 318566 158677 318626 159430
rect 320958 158677 321018 159430
rect 323350 159430 323428 159490
rect 325926 159430 326012 159490
rect 323350 158677 323410 159430
rect 325926 158677 325986 159430
rect 313411 158676 313477 158677
rect 313411 158612 313412 158676
rect 313476 158612 313477 158676
rect 313411 158611 313477 158612
rect 315803 158676 315869 158677
rect 315803 158612 315804 158676
rect 315868 158612 315869 158676
rect 315803 158611 315869 158612
rect 318563 158676 318629 158677
rect 318563 158612 318564 158676
rect 318628 158612 318629 158676
rect 318563 158611 318629 158612
rect 320955 158676 321021 158677
rect 320955 158612 320956 158676
rect 321020 158612 321021 158676
rect 320955 158611 321021 158612
rect 323347 158676 323413 158677
rect 323347 158612 323348 158676
rect 323412 158612 323413 158676
rect 323347 158611 323413 158612
rect 325923 158676 325989 158677
rect 325923 158612 325924 158676
rect 325988 158612 325989 158676
rect 325923 158611 325989 158612
rect 311019 158268 311085 158269
rect 311019 158204 311020 158268
rect 311084 158204 311085 158268
rect 311019 158203 311085 158204
rect 293539 157588 293605 157589
rect 293539 157524 293540 157588
rect 293604 157524 293605 157588
rect 293539 157523 293605 157524
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -656 290414 2898
rect 289794 -892 289826 -656
rect 290062 -892 290146 -656
rect 290382 -892 290414 -656
rect 289794 -976 290414 -892
rect 289794 -1212 289826 -976
rect 290062 -1212 290146 -976
rect 290382 -1212 290414 -976
rect 289794 -7964 290414 -1212
rect 294294 151954 294914 158000
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1616 294914 7398
rect 294294 -1852 294326 -1616
rect 294562 -1852 294646 -1616
rect 294882 -1852 294914 -1616
rect 294294 -1936 294914 -1852
rect 294294 -2172 294326 -1936
rect 294562 -2172 294646 -1936
rect 294882 -2172 294914 -1936
rect 294294 -7964 294914 -2172
rect 298794 156454 299414 158000
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2576 299414 11898
rect 298794 -2812 298826 -2576
rect 299062 -2812 299146 -2576
rect 299382 -2812 299414 -2576
rect 298794 -2896 299414 -2812
rect 298794 -3132 298826 -2896
rect 299062 -3132 299146 -2896
rect 299382 -3132 299414 -2896
rect 298794 -7964 299414 -3132
rect 303294 124954 303914 158000
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3536 303914 16398
rect 303294 -3772 303326 -3536
rect 303562 -3772 303646 -3536
rect 303882 -3772 303914 -3536
rect 303294 -3856 303914 -3772
rect 303294 -4092 303326 -3856
rect 303562 -4092 303646 -3856
rect 303882 -4092 303914 -3856
rect 303294 -7964 303914 -4092
rect 307794 129454 308414 158000
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4496 308414 20898
rect 307794 -4732 307826 -4496
rect 308062 -4732 308146 -4496
rect 308382 -4732 308414 -4496
rect 307794 -4816 308414 -4732
rect 307794 -5052 307826 -4816
rect 308062 -5052 308146 -4816
rect 308382 -5052 308414 -4816
rect 307794 -7964 308414 -5052
rect 312294 133954 312914 158000
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5456 312914 25398
rect 312294 -5692 312326 -5456
rect 312562 -5692 312646 -5456
rect 312882 -5692 312914 -5456
rect 312294 -5776 312914 -5692
rect 312294 -6012 312326 -5776
rect 312562 -6012 312646 -5776
rect 312882 -6012 312914 -5776
rect 312294 -7964 312914 -6012
rect 316794 138454 317414 158000
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6416 317414 29898
rect 316794 -6652 316826 -6416
rect 317062 -6652 317146 -6416
rect 317382 -6652 317414 -6416
rect 316794 -6736 317414 -6652
rect 316794 -6972 316826 -6736
rect 317062 -6972 317146 -6736
rect 317382 -6972 317414 -6736
rect 316794 -7964 317414 -6972
rect 321294 142954 321914 158000
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7376 321914 34398
rect 321294 -7612 321326 -7376
rect 321562 -7612 321646 -7376
rect 321882 -7612 321914 -7376
rect 321294 -7696 321914 -7612
rect 321294 -7932 321326 -7696
rect 321562 -7932 321646 -7696
rect 321882 -7932 321914 -7696
rect 321294 -7964 321914 -7932
rect 325794 147454 326414 158000
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -656 326414 2898
rect 325794 -892 325826 -656
rect 326062 -892 326146 -656
rect 326382 -892 326414 -656
rect 325794 -976 326414 -892
rect 325794 -1212 325826 -976
rect 326062 -1212 326146 -976
rect 326382 -1212 326414 -976
rect 325794 -7964 326414 -1212
rect 330294 151954 330914 158000
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1616 330914 7398
rect 330294 -1852 330326 -1616
rect 330562 -1852 330646 -1616
rect 330882 -1852 330914 -1616
rect 330294 -1936 330914 -1852
rect 330294 -2172 330326 -1936
rect 330562 -2172 330646 -1936
rect 330882 -2172 330914 -1936
rect 330294 -7964 330914 -2172
rect 334794 156454 335414 158000
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2576 335414 11898
rect 334794 -2812 334826 -2576
rect 335062 -2812 335146 -2576
rect 335382 -2812 335414 -2576
rect 334794 -2896 335414 -2812
rect 334794 -3132 334826 -2896
rect 335062 -3132 335146 -2896
rect 335382 -3132 335414 -2896
rect 334794 -7964 335414 -3132
rect 339294 124954 339914 158000
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3536 339914 16398
rect 339294 -3772 339326 -3536
rect 339562 -3772 339646 -3536
rect 339882 -3772 339914 -3536
rect 339294 -3856 339914 -3772
rect 339294 -4092 339326 -3856
rect 339562 -4092 339646 -3856
rect 339882 -4092 339914 -3856
rect 339294 -7964 339914 -4092
rect 343794 129454 344414 158000
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4496 344414 20898
rect 343794 -4732 343826 -4496
rect 344062 -4732 344146 -4496
rect 344382 -4732 344414 -4496
rect 343794 -4816 344414 -4732
rect 343794 -5052 343826 -4816
rect 344062 -5052 344146 -4816
rect 344382 -5052 344414 -4816
rect 343794 -7964 344414 -5052
rect 348294 133954 348914 158000
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5456 348914 25398
rect 348294 -5692 348326 -5456
rect 348562 -5692 348646 -5456
rect 348882 -5692 348914 -5456
rect 348294 -5776 348914 -5692
rect 348294 -6012 348326 -5776
rect 348562 -6012 348646 -5776
rect 348882 -6012 348914 -5776
rect 348294 -7964 348914 -6012
rect 352794 138454 353414 158000
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6416 353414 29898
rect 352794 -6652 352826 -6416
rect 353062 -6652 353146 -6416
rect 353382 -6652 353414 -6416
rect 352794 -6736 353414 -6652
rect 352794 -6972 352826 -6736
rect 353062 -6972 353146 -6736
rect 353382 -6972 353414 -6736
rect 352794 -7964 353414 -6972
rect 357294 142954 357914 158000
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7376 357914 34398
rect 358126 6357 358186 250819
rect 358675 245580 358741 245581
rect 358675 245516 358676 245580
rect 358740 245516 358741 245580
rect 358675 245515 358741 245516
rect 358307 244764 358373 244765
rect 358307 244700 358308 244764
rect 358372 244700 358373 244764
rect 358307 244699 358373 244700
rect 358123 6356 358189 6357
rect 358123 6292 358124 6356
rect 358188 6292 358189 6356
rect 358123 6291 358189 6292
rect 358310 3501 358370 244699
rect 358491 243540 358557 243541
rect 358491 243476 358492 243540
rect 358556 243476 358557 243540
rect 358491 243475 358557 243476
rect 358494 3637 358554 243475
rect 358678 158813 358738 245515
rect 358675 158812 358741 158813
rect 358675 158748 358676 158812
rect 358740 158748 358741 158812
rect 358675 158747 358741 158748
rect 358491 3636 358557 3637
rect 358491 3572 358492 3636
rect 358556 3572 358557 3636
rect 358491 3571 358557 3572
rect 358862 3501 358922 251907
rect 360147 248300 360213 248301
rect 360147 248236 360148 248300
rect 360212 248236 360213 248300
rect 360147 248235 360213 248236
rect 359043 248164 359109 248165
rect 359043 248100 359044 248164
rect 359108 248100 359109 248164
rect 359043 248099 359109 248100
rect 359046 3773 359106 248099
rect 359411 245308 359477 245309
rect 359411 245244 359412 245308
rect 359476 245244 359477 245308
rect 359411 245243 359477 245244
rect 359227 245172 359293 245173
rect 359227 245108 359228 245172
rect 359292 245108 359293 245172
rect 359227 245107 359293 245108
rect 359043 3772 359109 3773
rect 359043 3708 359044 3772
rect 359108 3708 359109 3772
rect 359043 3707 359109 3708
rect 358307 3500 358373 3501
rect 358307 3436 358308 3500
rect 358372 3436 358373 3500
rect 358307 3435 358373 3436
rect 358859 3500 358925 3501
rect 358859 3436 358860 3500
rect 358924 3436 358925 3500
rect 358859 3435 358925 3436
rect 359230 3365 359290 245107
rect 359414 3909 359474 245243
rect 359411 3908 359477 3909
rect 359411 3844 359412 3908
rect 359476 3844 359477 3908
rect 359411 3843 359477 3844
rect 360150 3501 360210 248235
rect 360699 245444 360765 245445
rect 360699 245380 360700 245444
rect 360764 245380 360765 245444
rect 360699 245379 360765 245380
rect 360515 245036 360581 245037
rect 360515 244972 360516 245036
rect 360580 244972 360581 245036
rect 360515 244971 360581 244972
rect 360331 244900 360397 244901
rect 360331 244836 360332 244900
rect 360396 244836 360397 244900
rect 360331 244835 360397 244836
rect 360334 4045 360394 244835
rect 360331 4044 360397 4045
rect 360331 3980 360332 4044
rect 360396 3980 360397 4044
rect 360331 3979 360397 3980
rect 360147 3500 360213 3501
rect 360147 3436 360148 3500
rect 360212 3436 360213 3500
rect 360147 3435 360213 3436
rect 359227 3364 359293 3365
rect 359227 3300 359228 3364
rect 359292 3300 359293 3364
rect 359227 3299 359293 3300
rect 360518 3229 360578 244971
rect 360702 158813 360762 245379
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 360699 158812 360765 158813
rect 360699 158748 360700 158812
rect 360764 158748 360765 158812
rect 360699 158747 360765 158748
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 362542 71909 362602 443259
rect 362723 441692 362789 441693
rect 362723 441628 362724 441692
rect 362788 441628 362789 441692
rect 362723 441627 362789 441628
rect 362726 231981 362786 441627
rect 364379 258772 364445 258773
rect 364379 258708 364380 258772
rect 364444 258708 364445 258772
rect 364379 258707 364445 258708
rect 362907 251836 362973 251837
rect 362907 251772 362908 251836
rect 362972 251772 362973 251836
rect 362907 251771 362973 251772
rect 362723 231980 362789 231981
rect 362723 231916 362724 231980
rect 362788 231916 362789 231980
rect 362723 231915 362789 231916
rect 362539 71908 362605 71909
rect 362539 71844 362540 71908
rect 362604 71844 362605 71908
rect 362539 71843 362605 71844
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 362910 3501 362970 251771
rect 363091 250748 363157 250749
rect 363091 250684 363092 250748
rect 363156 250684 363157 250748
rect 363091 250683 363157 250684
rect 363094 6493 363154 250683
rect 363275 250612 363341 250613
rect 363275 250548 363276 250612
rect 363340 250548 363341 250612
rect 363275 250547 363341 250548
rect 363278 6629 363338 250547
rect 363459 248028 363525 248029
rect 363459 247964 363460 248028
rect 363524 247964 363525 248028
rect 363459 247963 363525 247964
rect 363462 6901 363522 247963
rect 363459 6900 363525 6901
rect 363459 6836 363460 6900
rect 363524 6836 363525 6900
rect 363459 6835 363525 6836
rect 363275 6628 363341 6629
rect 363275 6564 363276 6628
rect 363340 6564 363341 6628
rect 363275 6563 363341 6564
rect 363091 6492 363157 6493
rect 363091 6428 363092 6492
rect 363156 6428 363157 6492
rect 363091 6427 363157 6428
rect 364382 3501 364442 258707
rect 364747 247892 364813 247893
rect 364747 247828 364748 247892
rect 364812 247828 364813 247892
rect 364747 247827 364813 247828
rect 364563 247756 364629 247757
rect 364563 247692 364564 247756
rect 364628 247692 364629 247756
rect 364563 247691 364629 247692
rect 360515 3228 360581 3229
rect 360515 3164 360516 3228
rect 360580 3164 360581 3228
rect 360515 3163 360581 3164
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 362907 3500 362973 3501
rect 362907 3436 362908 3500
rect 362972 3436 362973 3500
rect 362907 3435 362973 3436
rect 364379 3500 364445 3501
rect 364379 3436 364380 3500
rect 364444 3436 364445 3500
rect 364379 3435 364445 3436
rect 357294 -7612 357326 -7376
rect 357562 -7612 357646 -7376
rect 357882 -7612 357914 -7376
rect 357294 -7696 357914 -7612
rect 357294 -7932 357326 -7696
rect 357562 -7932 357646 -7696
rect 357882 -7932 357914 -7696
rect 357294 -7964 357914 -7932
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 364566 3093 364626 247691
rect 364750 158813 364810 247827
rect 364747 158812 364813 158813
rect 364747 158748 364748 158812
rect 364812 158748 364813 158812
rect 364747 158747 364813 158748
rect 364934 45661 364994 444619
rect 366294 439954 366914 475398
rect 370794 707068 371414 711900
rect 370794 706832 370826 707068
rect 371062 706832 371146 707068
rect 371382 706832 371414 707068
rect 370794 706748 371414 706832
rect 370794 706512 370826 706748
rect 371062 706512 371146 706748
rect 371382 706512 371414 706748
rect 370794 696454 371414 706512
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 369347 445908 369413 445909
rect 369347 445844 369348 445908
rect 369412 445844 369413 445908
rect 369347 445843 369413 445844
rect 367875 445772 367941 445773
rect 367875 445708 367876 445772
rect 367940 445708 367941 445772
rect 367875 445707 367941 445708
rect 367691 444412 367757 444413
rect 367691 444348 367692 444412
rect 367756 444348 367757 444412
rect 367691 444347 367757 444348
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 367139 286380 367205 286381
rect 367139 286316 367140 286380
rect 367204 286316 367205 286380
rect 367139 286315 367205 286316
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 365667 254692 365733 254693
rect 365667 254628 365668 254692
rect 365732 254628 365733 254692
rect 365667 254627 365733 254628
rect 364931 45660 364997 45661
rect 364931 45596 364932 45660
rect 364996 45596 364997 45660
rect 364931 45595 364997 45596
rect 365670 3637 365730 254627
rect 365851 253196 365917 253197
rect 365851 253132 365852 253196
rect 365916 253132 365917 253196
rect 365851 253131 365917 253132
rect 365667 3636 365733 3637
rect 365667 3572 365668 3636
rect 365732 3572 365733 3636
rect 365667 3571 365733 3572
rect 365854 3501 365914 253131
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 365851 3500 365917 3501
rect 365851 3436 365852 3500
rect 365916 3436 365917 3500
rect 365851 3435 365917 3436
rect 364563 3092 364629 3093
rect 364563 3028 364564 3092
rect 364628 3028 364629 3092
rect 364563 3027 364629 3028
rect 361794 -656 362414 2898
rect 361794 -892 361826 -656
rect 362062 -892 362146 -656
rect 362382 -892 362414 -656
rect 361794 -976 362414 -892
rect 361794 -1212 361826 -976
rect 362062 -1212 362146 -976
rect 362382 -1212 362414 -976
rect 361794 -7964 362414 -1212
rect 366294 -1616 366914 7398
rect 367142 3501 367202 286315
rect 367323 250476 367389 250477
rect 367323 250412 367324 250476
rect 367388 250412 367389 250476
rect 367323 250411 367389 250412
rect 367326 6221 367386 250411
rect 367694 85645 367754 444347
rect 367878 99517 367938 445707
rect 368979 444548 369045 444549
rect 368979 444484 368980 444548
rect 369044 444484 369045 444548
rect 368979 444483 369045 444484
rect 368427 300116 368493 300117
rect 368427 300052 368428 300116
rect 368492 300052 368493 300116
rect 368427 300051 368493 300052
rect 368430 155413 368490 300051
rect 368427 155412 368493 155413
rect 368427 155348 368428 155412
rect 368492 155348 368493 155412
rect 368427 155347 368493 155348
rect 368982 125629 369042 444483
rect 369163 254556 369229 254557
rect 369163 254492 369164 254556
rect 369228 254492 369229 254556
rect 369163 254491 369229 254492
rect 368979 125628 369045 125629
rect 368979 125564 368980 125628
rect 369044 125564 369045 125628
rect 368979 125563 369045 125564
rect 367875 99516 367941 99517
rect 367875 99452 367876 99516
rect 367940 99452 367941 99516
rect 367875 99451 367941 99452
rect 367691 85644 367757 85645
rect 367691 85580 367692 85644
rect 367756 85580 367757 85644
rect 367691 85579 367757 85580
rect 367323 6220 367389 6221
rect 367323 6156 367324 6220
rect 367388 6156 367389 6220
rect 367323 6155 367389 6156
rect 367139 3500 367205 3501
rect 367139 3436 367140 3500
rect 367204 3436 367205 3500
rect 367139 3435 367205 3436
rect 369166 3365 369226 254491
rect 369350 218109 369410 445843
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 369899 303516 369965 303517
rect 369899 303452 369900 303516
rect 369964 303452 369965 303516
rect 369899 303451 369965 303452
rect 369347 218108 369413 218109
rect 369347 218044 369348 218108
rect 369412 218044 369413 218108
rect 369347 218043 369413 218044
rect 369902 3501 369962 303451
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 369899 3500 369965 3501
rect 369899 3436 369900 3500
rect 369964 3436 369965 3500
rect 369899 3435 369965 3436
rect 369163 3364 369229 3365
rect 369163 3300 369164 3364
rect 369228 3300 369229 3364
rect 369163 3299 369229 3300
rect 366294 -1852 366326 -1616
rect 366562 -1852 366646 -1616
rect 366882 -1852 366914 -1616
rect 366294 -1936 366914 -1852
rect 366294 -2172 366326 -1936
rect 366562 -2172 366646 -1936
rect 366882 -2172 366914 -1936
rect 366294 -7964 366914 -2172
rect 370794 -2576 371414 11898
rect 370794 -2812 370826 -2576
rect 371062 -2812 371146 -2576
rect 371382 -2812 371414 -2576
rect 370794 -2896 371414 -2812
rect 370794 -3132 370826 -2896
rect 371062 -3132 371146 -2896
rect 371382 -3132 371414 -2896
rect 370794 -7964 371414 -3132
rect 375294 708028 375914 711900
rect 375294 707792 375326 708028
rect 375562 707792 375646 708028
rect 375882 707792 375914 708028
rect 375294 707708 375914 707792
rect 375294 707472 375326 707708
rect 375562 707472 375646 707708
rect 375882 707472 375914 707708
rect 375294 700954 375914 707472
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3536 375914 16398
rect 375294 -3772 375326 -3536
rect 375562 -3772 375646 -3536
rect 375882 -3772 375914 -3536
rect 375294 -3856 375914 -3772
rect 375294 -4092 375326 -3856
rect 375562 -4092 375646 -3856
rect 375882 -4092 375914 -3856
rect 375294 -7964 375914 -4092
rect 379794 708988 380414 711900
rect 379794 708752 379826 708988
rect 380062 708752 380146 708988
rect 380382 708752 380414 708988
rect 379794 708668 380414 708752
rect 379794 708432 379826 708668
rect 380062 708432 380146 708668
rect 380382 708432 380414 708668
rect 379794 669454 380414 708432
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4496 380414 20898
rect 379794 -4732 379826 -4496
rect 380062 -4732 380146 -4496
rect 380382 -4732 380414 -4496
rect 379794 -4816 380414 -4732
rect 379794 -5052 379826 -4816
rect 380062 -5052 380146 -4816
rect 380382 -5052 380414 -4816
rect 379794 -7964 380414 -5052
rect 384294 709948 384914 711900
rect 384294 709712 384326 709948
rect 384562 709712 384646 709948
rect 384882 709712 384914 709948
rect 384294 709628 384914 709712
rect 384294 709392 384326 709628
rect 384562 709392 384646 709628
rect 384882 709392 384914 709628
rect 384294 673954 384914 709392
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5456 384914 25398
rect 384294 -5692 384326 -5456
rect 384562 -5692 384646 -5456
rect 384882 -5692 384914 -5456
rect 384294 -5776 384914 -5692
rect 384294 -6012 384326 -5776
rect 384562 -6012 384646 -5776
rect 384882 -6012 384914 -5776
rect 384294 -7964 384914 -6012
rect 388794 710908 389414 711900
rect 388794 710672 388826 710908
rect 389062 710672 389146 710908
rect 389382 710672 389414 710908
rect 388794 710588 389414 710672
rect 388794 710352 388826 710588
rect 389062 710352 389146 710588
rect 389382 710352 389414 710588
rect 388794 678454 389414 710352
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 210454 389414 245898
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6416 389414 29898
rect 388794 -6652 388826 -6416
rect 389062 -6652 389146 -6416
rect 389382 -6652 389414 -6416
rect 388794 -6736 389414 -6652
rect 388794 -6972 388826 -6736
rect 389062 -6972 389146 -6736
rect 389382 -6972 389414 -6736
rect 388794 -7964 389414 -6972
rect 393294 711868 393914 711900
rect 393294 711632 393326 711868
rect 393562 711632 393646 711868
rect 393882 711632 393914 711868
rect 393294 711548 393914 711632
rect 393294 711312 393326 711548
rect 393562 711312 393646 711548
rect 393882 711312 393914 711548
rect 393294 682954 393914 711312
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 214954 393914 250398
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7376 393914 34398
rect 393294 -7612 393326 -7376
rect 393562 -7612 393646 -7376
rect 393882 -7612 393914 -7376
rect 393294 -7696 393914 -7612
rect 393294 -7932 393326 -7696
rect 393562 -7932 393646 -7696
rect 393882 -7932 393914 -7696
rect 393294 -7964 393914 -7932
rect 397794 705148 398414 711900
rect 397794 704912 397826 705148
rect 398062 704912 398146 705148
rect 398382 704912 398414 705148
rect 397794 704828 398414 704912
rect 397794 704592 397826 704828
rect 398062 704592 398146 704828
rect 398382 704592 398414 704828
rect 397794 687454 398414 704592
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -656 398414 2898
rect 397794 -892 397826 -656
rect 398062 -892 398146 -656
rect 398382 -892 398414 -656
rect 397794 -976 398414 -892
rect 397794 -1212 397826 -976
rect 398062 -1212 398146 -976
rect 398382 -1212 398414 -976
rect 397794 -7964 398414 -1212
rect 402294 706108 402914 711900
rect 402294 705872 402326 706108
rect 402562 705872 402646 706108
rect 402882 705872 402914 706108
rect 402294 705788 402914 705872
rect 402294 705552 402326 705788
rect 402562 705552 402646 705788
rect 402882 705552 402914 705788
rect 402294 691954 402914 705552
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1616 402914 7398
rect 402294 -1852 402326 -1616
rect 402562 -1852 402646 -1616
rect 402882 -1852 402914 -1616
rect 402294 -1936 402914 -1852
rect 402294 -2172 402326 -1936
rect 402562 -2172 402646 -1936
rect 402882 -2172 402914 -1936
rect 402294 -7964 402914 -2172
rect 406794 707068 407414 711900
rect 406794 706832 406826 707068
rect 407062 706832 407146 707068
rect 407382 706832 407414 707068
rect 406794 706748 407414 706832
rect 406794 706512 406826 706748
rect 407062 706512 407146 706748
rect 407382 706512 407414 706748
rect 406794 696454 407414 706512
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2576 407414 11898
rect 406794 -2812 406826 -2576
rect 407062 -2812 407146 -2576
rect 407382 -2812 407414 -2576
rect 406794 -2896 407414 -2812
rect 406794 -3132 406826 -2896
rect 407062 -3132 407146 -2896
rect 407382 -3132 407414 -2896
rect 406794 -7964 407414 -3132
rect 411294 708028 411914 711900
rect 411294 707792 411326 708028
rect 411562 707792 411646 708028
rect 411882 707792 411914 708028
rect 411294 707708 411914 707792
rect 411294 707472 411326 707708
rect 411562 707472 411646 707708
rect 411882 707472 411914 707708
rect 411294 700954 411914 707472
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3536 411914 16398
rect 411294 -3772 411326 -3536
rect 411562 -3772 411646 -3536
rect 411882 -3772 411914 -3536
rect 411294 -3856 411914 -3772
rect 411294 -4092 411326 -3856
rect 411562 -4092 411646 -3856
rect 411882 -4092 411914 -3856
rect 411294 -7964 411914 -4092
rect 415794 708988 416414 711900
rect 415794 708752 415826 708988
rect 416062 708752 416146 708988
rect 416382 708752 416414 708988
rect 415794 708668 416414 708752
rect 415794 708432 415826 708668
rect 416062 708432 416146 708668
rect 416382 708432 416414 708668
rect 415794 669454 416414 708432
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4496 416414 20898
rect 415794 -4732 415826 -4496
rect 416062 -4732 416146 -4496
rect 416382 -4732 416414 -4496
rect 415794 -4816 416414 -4732
rect 415794 -5052 415826 -4816
rect 416062 -5052 416146 -4816
rect 416382 -5052 416414 -4816
rect 415794 -7964 416414 -5052
rect 420294 709948 420914 711900
rect 420294 709712 420326 709948
rect 420562 709712 420646 709948
rect 420882 709712 420914 709948
rect 420294 709628 420914 709712
rect 420294 709392 420326 709628
rect 420562 709392 420646 709628
rect 420882 709392 420914 709628
rect 420294 673954 420914 709392
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5456 420914 25398
rect 420294 -5692 420326 -5456
rect 420562 -5692 420646 -5456
rect 420882 -5692 420914 -5456
rect 420294 -5776 420914 -5692
rect 420294 -6012 420326 -5776
rect 420562 -6012 420646 -5776
rect 420882 -6012 420914 -5776
rect 420294 -7964 420914 -6012
rect 424794 710908 425414 711900
rect 424794 710672 424826 710908
rect 425062 710672 425146 710908
rect 425382 710672 425414 710908
rect 424794 710588 425414 710672
rect 424794 710352 424826 710588
rect 425062 710352 425146 710588
rect 425382 710352 425414 710588
rect 424794 678454 425414 710352
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6416 425414 29898
rect 424794 -6652 424826 -6416
rect 425062 -6652 425146 -6416
rect 425382 -6652 425414 -6416
rect 424794 -6736 425414 -6652
rect 424794 -6972 424826 -6736
rect 425062 -6972 425146 -6736
rect 425382 -6972 425414 -6736
rect 424794 -7964 425414 -6972
rect 429294 711868 429914 711900
rect 429294 711632 429326 711868
rect 429562 711632 429646 711868
rect 429882 711632 429914 711868
rect 429294 711548 429914 711632
rect 429294 711312 429326 711548
rect 429562 711312 429646 711548
rect 429882 711312 429914 711548
rect 429294 682954 429914 711312
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7376 429914 34398
rect 429294 -7612 429326 -7376
rect 429562 -7612 429646 -7376
rect 429882 -7612 429914 -7376
rect 429294 -7696 429914 -7612
rect 429294 -7932 429326 -7696
rect 429562 -7932 429646 -7696
rect 429882 -7932 429914 -7696
rect 429294 -7964 429914 -7932
rect 433794 705148 434414 711900
rect 433794 704912 433826 705148
rect 434062 704912 434146 705148
rect 434382 704912 434414 705148
rect 433794 704828 434414 704912
rect 433794 704592 433826 704828
rect 434062 704592 434146 704828
rect 434382 704592 434414 704828
rect 433794 687454 434414 704592
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -656 434414 2898
rect 433794 -892 433826 -656
rect 434062 -892 434146 -656
rect 434382 -892 434414 -656
rect 433794 -976 434414 -892
rect 433794 -1212 433826 -976
rect 434062 -1212 434146 -976
rect 434382 -1212 434414 -976
rect 433794 -7964 434414 -1212
rect 438294 706108 438914 711900
rect 438294 705872 438326 706108
rect 438562 705872 438646 706108
rect 438882 705872 438914 706108
rect 438294 705788 438914 705872
rect 438294 705552 438326 705788
rect 438562 705552 438646 705788
rect 438882 705552 438914 705788
rect 438294 691954 438914 705552
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1616 438914 7398
rect 438294 -1852 438326 -1616
rect 438562 -1852 438646 -1616
rect 438882 -1852 438914 -1616
rect 438294 -1936 438914 -1852
rect 438294 -2172 438326 -1936
rect 438562 -2172 438646 -1936
rect 438882 -2172 438914 -1936
rect 438294 -7964 438914 -2172
rect 442794 707068 443414 711900
rect 442794 706832 442826 707068
rect 443062 706832 443146 707068
rect 443382 706832 443414 707068
rect 442794 706748 443414 706832
rect 442794 706512 442826 706748
rect 443062 706512 443146 706748
rect 443382 706512 443414 706748
rect 442794 696454 443414 706512
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2576 443414 11898
rect 442794 -2812 442826 -2576
rect 443062 -2812 443146 -2576
rect 443382 -2812 443414 -2576
rect 442794 -2896 443414 -2812
rect 442794 -3132 442826 -2896
rect 443062 -3132 443146 -2896
rect 443382 -3132 443414 -2896
rect 442794 -7964 443414 -3132
rect 447294 708028 447914 711900
rect 447294 707792 447326 708028
rect 447562 707792 447646 708028
rect 447882 707792 447914 708028
rect 447294 707708 447914 707792
rect 447294 707472 447326 707708
rect 447562 707472 447646 707708
rect 447882 707472 447914 707708
rect 447294 700954 447914 707472
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3536 447914 16398
rect 447294 -3772 447326 -3536
rect 447562 -3772 447646 -3536
rect 447882 -3772 447914 -3536
rect 447294 -3856 447914 -3772
rect 447294 -4092 447326 -3856
rect 447562 -4092 447646 -3856
rect 447882 -4092 447914 -3856
rect 447294 -7964 447914 -4092
rect 451794 708988 452414 711900
rect 451794 708752 451826 708988
rect 452062 708752 452146 708988
rect 452382 708752 452414 708988
rect 451794 708668 452414 708752
rect 451794 708432 451826 708668
rect 452062 708432 452146 708668
rect 452382 708432 452414 708668
rect 451794 669454 452414 708432
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4496 452414 20898
rect 451794 -4732 451826 -4496
rect 452062 -4732 452146 -4496
rect 452382 -4732 452414 -4496
rect 451794 -4816 452414 -4732
rect 451794 -5052 451826 -4816
rect 452062 -5052 452146 -4816
rect 452382 -5052 452414 -4816
rect 451794 -7964 452414 -5052
rect 456294 709948 456914 711900
rect 456294 709712 456326 709948
rect 456562 709712 456646 709948
rect 456882 709712 456914 709948
rect 456294 709628 456914 709712
rect 456294 709392 456326 709628
rect 456562 709392 456646 709628
rect 456882 709392 456914 709628
rect 456294 673954 456914 709392
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5456 456914 25398
rect 456294 -5692 456326 -5456
rect 456562 -5692 456646 -5456
rect 456882 -5692 456914 -5456
rect 456294 -5776 456914 -5692
rect 456294 -6012 456326 -5776
rect 456562 -6012 456646 -5776
rect 456882 -6012 456914 -5776
rect 456294 -7964 456914 -6012
rect 460794 710908 461414 711900
rect 460794 710672 460826 710908
rect 461062 710672 461146 710908
rect 461382 710672 461414 710908
rect 460794 710588 461414 710672
rect 460794 710352 460826 710588
rect 461062 710352 461146 710588
rect 461382 710352 461414 710588
rect 460794 678454 461414 710352
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6416 461414 29898
rect 460794 -6652 460826 -6416
rect 461062 -6652 461146 -6416
rect 461382 -6652 461414 -6416
rect 460794 -6736 461414 -6652
rect 460794 -6972 460826 -6736
rect 461062 -6972 461146 -6736
rect 461382 -6972 461414 -6736
rect 460794 -7964 461414 -6972
rect 465294 711868 465914 711900
rect 465294 711632 465326 711868
rect 465562 711632 465646 711868
rect 465882 711632 465914 711868
rect 465294 711548 465914 711632
rect 465294 711312 465326 711548
rect 465562 711312 465646 711548
rect 465882 711312 465914 711548
rect 465294 682954 465914 711312
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7376 465914 34398
rect 465294 -7612 465326 -7376
rect 465562 -7612 465646 -7376
rect 465882 -7612 465914 -7376
rect 465294 -7696 465914 -7612
rect 465294 -7932 465326 -7696
rect 465562 -7932 465646 -7696
rect 465882 -7932 465914 -7696
rect 465294 -7964 465914 -7932
rect 469794 705148 470414 711900
rect 469794 704912 469826 705148
rect 470062 704912 470146 705148
rect 470382 704912 470414 705148
rect 469794 704828 470414 704912
rect 469794 704592 469826 704828
rect 470062 704592 470146 704828
rect 470382 704592 470414 704828
rect 469794 687454 470414 704592
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -656 470414 2898
rect 469794 -892 469826 -656
rect 470062 -892 470146 -656
rect 470382 -892 470414 -656
rect 469794 -976 470414 -892
rect 469794 -1212 469826 -976
rect 470062 -1212 470146 -976
rect 470382 -1212 470414 -976
rect 469794 -7964 470414 -1212
rect 474294 706108 474914 711900
rect 474294 705872 474326 706108
rect 474562 705872 474646 706108
rect 474882 705872 474914 706108
rect 474294 705788 474914 705872
rect 474294 705552 474326 705788
rect 474562 705552 474646 705788
rect 474882 705552 474914 705788
rect 474294 691954 474914 705552
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1616 474914 7398
rect 474294 -1852 474326 -1616
rect 474562 -1852 474646 -1616
rect 474882 -1852 474914 -1616
rect 474294 -1936 474914 -1852
rect 474294 -2172 474326 -1936
rect 474562 -2172 474646 -1936
rect 474882 -2172 474914 -1936
rect 474294 -7964 474914 -2172
rect 478794 707068 479414 711900
rect 478794 706832 478826 707068
rect 479062 706832 479146 707068
rect 479382 706832 479414 707068
rect 478794 706748 479414 706832
rect 478794 706512 478826 706748
rect 479062 706512 479146 706748
rect 479382 706512 479414 706748
rect 478794 696454 479414 706512
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2576 479414 11898
rect 478794 -2812 478826 -2576
rect 479062 -2812 479146 -2576
rect 479382 -2812 479414 -2576
rect 478794 -2896 479414 -2812
rect 478794 -3132 478826 -2896
rect 479062 -3132 479146 -2896
rect 479382 -3132 479414 -2896
rect 478794 -7964 479414 -3132
rect 483294 708028 483914 711900
rect 483294 707792 483326 708028
rect 483562 707792 483646 708028
rect 483882 707792 483914 708028
rect 483294 707708 483914 707792
rect 483294 707472 483326 707708
rect 483562 707472 483646 707708
rect 483882 707472 483914 707708
rect 483294 700954 483914 707472
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3536 483914 16398
rect 483294 -3772 483326 -3536
rect 483562 -3772 483646 -3536
rect 483882 -3772 483914 -3536
rect 483294 -3856 483914 -3772
rect 483294 -4092 483326 -3856
rect 483562 -4092 483646 -3856
rect 483882 -4092 483914 -3856
rect 483294 -7964 483914 -4092
rect 487794 708988 488414 711900
rect 487794 708752 487826 708988
rect 488062 708752 488146 708988
rect 488382 708752 488414 708988
rect 487794 708668 488414 708752
rect 487794 708432 487826 708668
rect 488062 708432 488146 708668
rect 488382 708432 488414 708668
rect 487794 669454 488414 708432
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4496 488414 20898
rect 487794 -4732 487826 -4496
rect 488062 -4732 488146 -4496
rect 488382 -4732 488414 -4496
rect 487794 -4816 488414 -4732
rect 487794 -5052 487826 -4816
rect 488062 -5052 488146 -4816
rect 488382 -5052 488414 -4816
rect 487794 -7964 488414 -5052
rect 492294 709948 492914 711900
rect 492294 709712 492326 709948
rect 492562 709712 492646 709948
rect 492882 709712 492914 709948
rect 492294 709628 492914 709712
rect 492294 709392 492326 709628
rect 492562 709392 492646 709628
rect 492882 709392 492914 709628
rect 492294 673954 492914 709392
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5456 492914 25398
rect 492294 -5692 492326 -5456
rect 492562 -5692 492646 -5456
rect 492882 -5692 492914 -5456
rect 492294 -5776 492914 -5692
rect 492294 -6012 492326 -5776
rect 492562 -6012 492646 -5776
rect 492882 -6012 492914 -5776
rect 492294 -7964 492914 -6012
rect 496794 710908 497414 711900
rect 496794 710672 496826 710908
rect 497062 710672 497146 710908
rect 497382 710672 497414 710908
rect 496794 710588 497414 710672
rect 496794 710352 496826 710588
rect 497062 710352 497146 710588
rect 497382 710352 497414 710588
rect 496794 678454 497414 710352
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6416 497414 29898
rect 496794 -6652 496826 -6416
rect 497062 -6652 497146 -6416
rect 497382 -6652 497414 -6416
rect 496794 -6736 497414 -6652
rect 496794 -6972 496826 -6736
rect 497062 -6972 497146 -6736
rect 497382 -6972 497414 -6736
rect 496794 -7964 497414 -6972
rect 501294 711868 501914 711900
rect 501294 711632 501326 711868
rect 501562 711632 501646 711868
rect 501882 711632 501914 711868
rect 501294 711548 501914 711632
rect 501294 711312 501326 711548
rect 501562 711312 501646 711548
rect 501882 711312 501914 711548
rect 501294 682954 501914 711312
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7376 501914 34398
rect 501294 -7612 501326 -7376
rect 501562 -7612 501646 -7376
rect 501882 -7612 501914 -7376
rect 501294 -7696 501914 -7612
rect 501294 -7932 501326 -7696
rect 501562 -7932 501646 -7696
rect 501882 -7932 501914 -7696
rect 501294 -7964 501914 -7932
rect 505794 705148 506414 711900
rect 505794 704912 505826 705148
rect 506062 704912 506146 705148
rect 506382 704912 506414 705148
rect 505794 704828 506414 704912
rect 505794 704592 505826 704828
rect 506062 704592 506146 704828
rect 506382 704592 506414 704828
rect 505794 687454 506414 704592
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -656 506414 2898
rect 505794 -892 505826 -656
rect 506062 -892 506146 -656
rect 506382 -892 506414 -656
rect 505794 -976 506414 -892
rect 505794 -1212 505826 -976
rect 506062 -1212 506146 -976
rect 506382 -1212 506414 -976
rect 505794 -7964 506414 -1212
rect 510294 706108 510914 711900
rect 510294 705872 510326 706108
rect 510562 705872 510646 706108
rect 510882 705872 510914 706108
rect 510294 705788 510914 705872
rect 510294 705552 510326 705788
rect 510562 705552 510646 705788
rect 510882 705552 510914 705788
rect 510294 691954 510914 705552
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1616 510914 7398
rect 510294 -1852 510326 -1616
rect 510562 -1852 510646 -1616
rect 510882 -1852 510914 -1616
rect 510294 -1936 510914 -1852
rect 510294 -2172 510326 -1936
rect 510562 -2172 510646 -1936
rect 510882 -2172 510914 -1936
rect 510294 -7964 510914 -2172
rect 514794 707068 515414 711900
rect 514794 706832 514826 707068
rect 515062 706832 515146 707068
rect 515382 706832 515414 707068
rect 514794 706748 515414 706832
rect 514794 706512 514826 706748
rect 515062 706512 515146 706748
rect 515382 706512 515414 706748
rect 514794 696454 515414 706512
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2576 515414 11898
rect 514794 -2812 514826 -2576
rect 515062 -2812 515146 -2576
rect 515382 -2812 515414 -2576
rect 514794 -2896 515414 -2812
rect 514794 -3132 514826 -2896
rect 515062 -3132 515146 -2896
rect 515382 -3132 515414 -2896
rect 514794 -7964 515414 -3132
rect 519294 708028 519914 711900
rect 519294 707792 519326 708028
rect 519562 707792 519646 708028
rect 519882 707792 519914 708028
rect 519294 707708 519914 707792
rect 519294 707472 519326 707708
rect 519562 707472 519646 707708
rect 519882 707472 519914 707708
rect 519294 700954 519914 707472
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3536 519914 16398
rect 519294 -3772 519326 -3536
rect 519562 -3772 519646 -3536
rect 519882 -3772 519914 -3536
rect 519294 -3856 519914 -3772
rect 519294 -4092 519326 -3856
rect 519562 -4092 519646 -3856
rect 519882 -4092 519914 -3856
rect 519294 -7964 519914 -4092
rect 523794 708988 524414 711900
rect 523794 708752 523826 708988
rect 524062 708752 524146 708988
rect 524382 708752 524414 708988
rect 523794 708668 524414 708752
rect 523794 708432 523826 708668
rect 524062 708432 524146 708668
rect 524382 708432 524414 708668
rect 523794 669454 524414 708432
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4496 524414 20898
rect 523794 -4732 523826 -4496
rect 524062 -4732 524146 -4496
rect 524382 -4732 524414 -4496
rect 523794 -4816 524414 -4732
rect 523794 -5052 523826 -4816
rect 524062 -5052 524146 -4816
rect 524382 -5052 524414 -4816
rect 523794 -7964 524414 -5052
rect 528294 709948 528914 711900
rect 528294 709712 528326 709948
rect 528562 709712 528646 709948
rect 528882 709712 528914 709948
rect 528294 709628 528914 709712
rect 528294 709392 528326 709628
rect 528562 709392 528646 709628
rect 528882 709392 528914 709628
rect 528294 673954 528914 709392
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5456 528914 25398
rect 528294 -5692 528326 -5456
rect 528562 -5692 528646 -5456
rect 528882 -5692 528914 -5456
rect 528294 -5776 528914 -5692
rect 528294 -6012 528326 -5776
rect 528562 -6012 528646 -5776
rect 528882 -6012 528914 -5776
rect 528294 -7964 528914 -6012
rect 532794 710908 533414 711900
rect 532794 710672 532826 710908
rect 533062 710672 533146 710908
rect 533382 710672 533414 710908
rect 532794 710588 533414 710672
rect 532794 710352 532826 710588
rect 533062 710352 533146 710588
rect 533382 710352 533414 710588
rect 532794 678454 533414 710352
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6416 533414 29898
rect 532794 -6652 532826 -6416
rect 533062 -6652 533146 -6416
rect 533382 -6652 533414 -6416
rect 532794 -6736 533414 -6652
rect 532794 -6972 532826 -6736
rect 533062 -6972 533146 -6736
rect 533382 -6972 533414 -6736
rect 532794 -7964 533414 -6972
rect 537294 711868 537914 711900
rect 537294 711632 537326 711868
rect 537562 711632 537646 711868
rect 537882 711632 537914 711868
rect 537294 711548 537914 711632
rect 537294 711312 537326 711548
rect 537562 711312 537646 711548
rect 537882 711312 537914 711548
rect 537294 682954 537914 711312
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7376 537914 34398
rect 537294 -7612 537326 -7376
rect 537562 -7612 537646 -7376
rect 537882 -7612 537914 -7376
rect 537294 -7696 537914 -7612
rect 537294 -7932 537326 -7696
rect 537562 -7932 537646 -7696
rect 537882 -7932 537914 -7696
rect 537294 -7964 537914 -7932
rect 541794 705148 542414 711900
rect 541794 704912 541826 705148
rect 542062 704912 542146 705148
rect 542382 704912 542414 705148
rect 541794 704828 542414 704912
rect 541794 704592 541826 704828
rect 542062 704592 542146 704828
rect 542382 704592 542414 704828
rect 541794 687454 542414 704592
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -656 542414 2898
rect 541794 -892 541826 -656
rect 542062 -892 542146 -656
rect 542382 -892 542414 -656
rect 541794 -976 542414 -892
rect 541794 -1212 541826 -976
rect 542062 -1212 542146 -976
rect 542382 -1212 542414 -976
rect 541794 -7964 542414 -1212
rect 546294 706108 546914 711900
rect 546294 705872 546326 706108
rect 546562 705872 546646 706108
rect 546882 705872 546914 706108
rect 546294 705788 546914 705872
rect 546294 705552 546326 705788
rect 546562 705552 546646 705788
rect 546882 705552 546914 705788
rect 546294 691954 546914 705552
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1616 546914 7398
rect 546294 -1852 546326 -1616
rect 546562 -1852 546646 -1616
rect 546882 -1852 546914 -1616
rect 546294 -1936 546914 -1852
rect 546294 -2172 546326 -1936
rect 546562 -2172 546646 -1936
rect 546882 -2172 546914 -1936
rect 546294 -7964 546914 -2172
rect 550794 707068 551414 711900
rect 550794 706832 550826 707068
rect 551062 706832 551146 707068
rect 551382 706832 551414 707068
rect 550794 706748 551414 706832
rect 550794 706512 550826 706748
rect 551062 706512 551146 706748
rect 551382 706512 551414 706748
rect 550794 696454 551414 706512
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2576 551414 11898
rect 550794 -2812 550826 -2576
rect 551062 -2812 551146 -2576
rect 551382 -2812 551414 -2576
rect 550794 -2896 551414 -2812
rect 550794 -3132 550826 -2896
rect 551062 -3132 551146 -2896
rect 551382 -3132 551414 -2896
rect 550794 -7964 551414 -3132
rect 555294 708028 555914 711900
rect 555294 707792 555326 708028
rect 555562 707792 555646 708028
rect 555882 707792 555914 708028
rect 555294 707708 555914 707792
rect 555294 707472 555326 707708
rect 555562 707472 555646 707708
rect 555882 707472 555914 707708
rect 555294 700954 555914 707472
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3536 555914 16398
rect 555294 -3772 555326 -3536
rect 555562 -3772 555646 -3536
rect 555882 -3772 555914 -3536
rect 555294 -3856 555914 -3772
rect 555294 -4092 555326 -3856
rect 555562 -4092 555646 -3856
rect 555882 -4092 555914 -3856
rect 555294 -7964 555914 -4092
rect 559794 708988 560414 711900
rect 559794 708752 559826 708988
rect 560062 708752 560146 708988
rect 560382 708752 560414 708988
rect 559794 708668 560414 708752
rect 559794 708432 559826 708668
rect 560062 708432 560146 708668
rect 560382 708432 560414 708668
rect 559794 669454 560414 708432
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4496 560414 20898
rect 559794 -4732 559826 -4496
rect 560062 -4732 560146 -4496
rect 560382 -4732 560414 -4496
rect 559794 -4816 560414 -4732
rect 559794 -5052 559826 -4816
rect 560062 -5052 560146 -4816
rect 560382 -5052 560414 -4816
rect 559794 -7964 560414 -5052
rect 564294 709948 564914 711900
rect 564294 709712 564326 709948
rect 564562 709712 564646 709948
rect 564882 709712 564914 709948
rect 564294 709628 564914 709712
rect 564294 709392 564326 709628
rect 564562 709392 564646 709628
rect 564882 709392 564914 709628
rect 564294 673954 564914 709392
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5456 564914 25398
rect 564294 -5692 564326 -5456
rect 564562 -5692 564646 -5456
rect 564882 -5692 564914 -5456
rect 564294 -5776 564914 -5692
rect 564294 -6012 564326 -5776
rect 564562 -6012 564646 -5776
rect 564882 -6012 564914 -5776
rect 564294 -7964 564914 -6012
rect 568794 710908 569414 711900
rect 568794 710672 568826 710908
rect 569062 710672 569146 710908
rect 569382 710672 569414 710908
rect 568794 710588 569414 710672
rect 568794 710352 568826 710588
rect 569062 710352 569146 710588
rect 569382 710352 569414 710588
rect 568794 678454 569414 710352
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6416 569414 29898
rect 568794 -6652 568826 -6416
rect 569062 -6652 569146 -6416
rect 569382 -6652 569414 -6416
rect 568794 -6736 569414 -6652
rect 568794 -6972 568826 -6736
rect 569062 -6972 569146 -6736
rect 569382 -6972 569414 -6736
rect 568794 -7964 569414 -6972
rect 573294 711868 573914 711900
rect 573294 711632 573326 711868
rect 573562 711632 573646 711868
rect 573882 711632 573914 711868
rect 573294 711548 573914 711632
rect 573294 711312 573326 711548
rect 573562 711312 573646 711548
rect 573882 711312 573914 711548
rect 573294 682954 573914 711312
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7376 573914 34398
rect 573294 -7612 573326 -7376
rect 573562 -7612 573646 -7376
rect 573882 -7612 573914 -7376
rect 573294 -7696 573914 -7612
rect 573294 -7932 573326 -7696
rect 573562 -7932 573646 -7696
rect 573882 -7932 573914 -7696
rect 573294 -7964 573914 -7932
rect 577794 705148 578414 711900
rect 577794 704912 577826 705148
rect 578062 704912 578146 705148
rect 578382 704912 578414 705148
rect 577794 704828 578414 704912
rect 577794 704592 577826 704828
rect 578062 704592 578146 704828
rect 578382 704592 578414 704828
rect 577794 687454 578414 704592
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -656 578414 2898
rect 577794 -892 577826 -656
rect 578062 -892 578146 -656
rect 578382 -892 578414 -656
rect 577794 -976 578414 -892
rect 577794 -1212 577826 -976
rect 578062 -1212 578146 -976
rect 578382 -1212 578414 -976
rect 577794 -7964 578414 -1212
rect 582294 706108 582914 711900
rect 592340 711868 592960 711900
rect 592340 711632 592372 711868
rect 592608 711632 592692 711868
rect 592928 711632 592960 711868
rect 592340 711548 592960 711632
rect 592340 711312 592372 711548
rect 592608 711312 592692 711548
rect 592928 711312 592960 711548
rect 591380 710908 592000 710940
rect 591380 710672 591412 710908
rect 591648 710672 591732 710908
rect 591968 710672 592000 710908
rect 591380 710588 592000 710672
rect 591380 710352 591412 710588
rect 591648 710352 591732 710588
rect 591968 710352 592000 710588
rect 590420 709948 591040 709980
rect 590420 709712 590452 709948
rect 590688 709712 590772 709948
rect 591008 709712 591040 709948
rect 590420 709628 591040 709712
rect 590420 709392 590452 709628
rect 590688 709392 590772 709628
rect 591008 709392 591040 709628
rect 589460 708988 590080 709020
rect 589460 708752 589492 708988
rect 589728 708752 589812 708988
rect 590048 708752 590080 708988
rect 589460 708668 590080 708752
rect 589460 708432 589492 708668
rect 589728 708432 589812 708668
rect 590048 708432 590080 708668
rect 588500 708028 589120 708060
rect 588500 707792 588532 708028
rect 588768 707792 588852 708028
rect 589088 707792 589120 708028
rect 588500 707708 589120 707792
rect 588500 707472 588532 707708
rect 588768 707472 588852 707708
rect 589088 707472 589120 707708
rect 587540 707068 588160 707100
rect 587540 706832 587572 707068
rect 587808 706832 587892 707068
rect 588128 706832 588160 707068
rect 587540 706748 588160 706832
rect 587540 706512 587572 706748
rect 587808 706512 587892 706748
rect 588128 706512 588160 706748
rect 582294 705872 582326 706108
rect 582562 705872 582646 706108
rect 582882 705872 582914 706108
rect 582294 705788 582914 705872
rect 582294 705552 582326 705788
rect 582562 705552 582646 705788
rect 582882 705552 582914 705788
rect 582294 691954 582914 705552
rect 586580 706108 587200 706140
rect 586580 705872 586612 706108
rect 586848 705872 586932 706108
rect 587168 705872 587200 706108
rect 586580 705788 587200 705872
rect 586580 705552 586612 705788
rect 586848 705552 586932 705788
rect 587168 705552 587200 705788
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1616 582914 7398
rect 585620 705148 586240 705180
rect 585620 704912 585652 705148
rect 585888 704912 585972 705148
rect 586208 704912 586240 705148
rect 585620 704828 586240 704912
rect 585620 704592 585652 704828
rect 585888 704592 585972 704828
rect 586208 704592 586240 704828
rect 585620 687454 586240 704592
rect 585620 687218 585652 687454
rect 585888 687218 585972 687454
rect 586208 687218 586240 687454
rect 585620 687134 586240 687218
rect 585620 686898 585652 687134
rect 585888 686898 585972 687134
rect 586208 686898 586240 687134
rect 585620 651454 586240 686898
rect 585620 651218 585652 651454
rect 585888 651218 585972 651454
rect 586208 651218 586240 651454
rect 585620 651134 586240 651218
rect 585620 650898 585652 651134
rect 585888 650898 585972 651134
rect 586208 650898 586240 651134
rect 585620 615454 586240 650898
rect 585620 615218 585652 615454
rect 585888 615218 585972 615454
rect 586208 615218 586240 615454
rect 585620 615134 586240 615218
rect 585620 614898 585652 615134
rect 585888 614898 585972 615134
rect 586208 614898 586240 615134
rect 585620 579454 586240 614898
rect 585620 579218 585652 579454
rect 585888 579218 585972 579454
rect 586208 579218 586240 579454
rect 585620 579134 586240 579218
rect 585620 578898 585652 579134
rect 585888 578898 585972 579134
rect 586208 578898 586240 579134
rect 585620 543454 586240 578898
rect 585620 543218 585652 543454
rect 585888 543218 585972 543454
rect 586208 543218 586240 543454
rect 585620 543134 586240 543218
rect 585620 542898 585652 543134
rect 585888 542898 585972 543134
rect 586208 542898 586240 543134
rect 585620 507454 586240 542898
rect 585620 507218 585652 507454
rect 585888 507218 585972 507454
rect 586208 507218 586240 507454
rect 585620 507134 586240 507218
rect 585620 506898 585652 507134
rect 585888 506898 585972 507134
rect 586208 506898 586240 507134
rect 585620 471454 586240 506898
rect 585620 471218 585652 471454
rect 585888 471218 585972 471454
rect 586208 471218 586240 471454
rect 585620 471134 586240 471218
rect 585620 470898 585652 471134
rect 585888 470898 585972 471134
rect 586208 470898 586240 471134
rect 585620 435454 586240 470898
rect 585620 435218 585652 435454
rect 585888 435218 585972 435454
rect 586208 435218 586240 435454
rect 585620 435134 586240 435218
rect 585620 434898 585652 435134
rect 585888 434898 585972 435134
rect 586208 434898 586240 435134
rect 585620 399454 586240 434898
rect 585620 399218 585652 399454
rect 585888 399218 585972 399454
rect 586208 399218 586240 399454
rect 585620 399134 586240 399218
rect 585620 398898 585652 399134
rect 585888 398898 585972 399134
rect 586208 398898 586240 399134
rect 585620 363454 586240 398898
rect 585620 363218 585652 363454
rect 585888 363218 585972 363454
rect 586208 363218 586240 363454
rect 585620 363134 586240 363218
rect 585620 362898 585652 363134
rect 585888 362898 585972 363134
rect 586208 362898 586240 363134
rect 585620 327454 586240 362898
rect 585620 327218 585652 327454
rect 585888 327218 585972 327454
rect 586208 327218 586240 327454
rect 585620 327134 586240 327218
rect 585620 326898 585652 327134
rect 585888 326898 585972 327134
rect 586208 326898 586240 327134
rect 585620 291454 586240 326898
rect 585620 291218 585652 291454
rect 585888 291218 585972 291454
rect 586208 291218 586240 291454
rect 585620 291134 586240 291218
rect 585620 290898 585652 291134
rect 585888 290898 585972 291134
rect 586208 290898 586240 291134
rect 585620 255454 586240 290898
rect 585620 255218 585652 255454
rect 585888 255218 585972 255454
rect 586208 255218 586240 255454
rect 585620 255134 586240 255218
rect 585620 254898 585652 255134
rect 585888 254898 585972 255134
rect 586208 254898 586240 255134
rect 585620 219454 586240 254898
rect 585620 219218 585652 219454
rect 585888 219218 585972 219454
rect 586208 219218 586240 219454
rect 585620 219134 586240 219218
rect 585620 218898 585652 219134
rect 585888 218898 585972 219134
rect 586208 218898 586240 219134
rect 585620 183454 586240 218898
rect 585620 183218 585652 183454
rect 585888 183218 585972 183454
rect 586208 183218 586240 183454
rect 585620 183134 586240 183218
rect 585620 182898 585652 183134
rect 585888 182898 585972 183134
rect 586208 182898 586240 183134
rect 585620 147454 586240 182898
rect 585620 147218 585652 147454
rect 585888 147218 585972 147454
rect 586208 147218 586240 147454
rect 585620 147134 586240 147218
rect 585620 146898 585652 147134
rect 585888 146898 585972 147134
rect 586208 146898 586240 147134
rect 585620 111454 586240 146898
rect 585620 111218 585652 111454
rect 585888 111218 585972 111454
rect 586208 111218 586240 111454
rect 585620 111134 586240 111218
rect 585620 110898 585652 111134
rect 585888 110898 585972 111134
rect 586208 110898 586240 111134
rect 585620 75454 586240 110898
rect 585620 75218 585652 75454
rect 585888 75218 585972 75454
rect 586208 75218 586240 75454
rect 585620 75134 586240 75218
rect 585620 74898 585652 75134
rect 585888 74898 585972 75134
rect 586208 74898 586240 75134
rect 585620 39454 586240 74898
rect 585620 39218 585652 39454
rect 585888 39218 585972 39454
rect 586208 39218 586240 39454
rect 585620 39134 586240 39218
rect 585620 38898 585652 39134
rect 585888 38898 585972 39134
rect 586208 38898 586240 39134
rect 585620 3454 586240 38898
rect 585620 3218 585652 3454
rect 585888 3218 585972 3454
rect 586208 3218 586240 3454
rect 585620 3134 586240 3218
rect 585620 2898 585652 3134
rect 585888 2898 585972 3134
rect 586208 2898 586240 3134
rect 585620 -656 586240 2898
rect 585620 -892 585652 -656
rect 585888 -892 585972 -656
rect 586208 -892 586240 -656
rect 585620 -976 586240 -892
rect 585620 -1212 585652 -976
rect 585888 -1212 585972 -976
rect 586208 -1212 586240 -976
rect 585620 -1244 586240 -1212
rect 586580 691954 587200 705552
rect 586580 691718 586612 691954
rect 586848 691718 586932 691954
rect 587168 691718 587200 691954
rect 586580 691634 587200 691718
rect 586580 691398 586612 691634
rect 586848 691398 586932 691634
rect 587168 691398 587200 691634
rect 586580 655954 587200 691398
rect 586580 655718 586612 655954
rect 586848 655718 586932 655954
rect 587168 655718 587200 655954
rect 586580 655634 587200 655718
rect 586580 655398 586612 655634
rect 586848 655398 586932 655634
rect 587168 655398 587200 655634
rect 586580 619954 587200 655398
rect 586580 619718 586612 619954
rect 586848 619718 586932 619954
rect 587168 619718 587200 619954
rect 586580 619634 587200 619718
rect 586580 619398 586612 619634
rect 586848 619398 586932 619634
rect 587168 619398 587200 619634
rect 586580 583954 587200 619398
rect 586580 583718 586612 583954
rect 586848 583718 586932 583954
rect 587168 583718 587200 583954
rect 586580 583634 587200 583718
rect 586580 583398 586612 583634
rect 586848 583398 586932 583634
rect 587168 583398 587200 583634
rect 586580 547954 587200 583398
rect 586580 547718 586612 547954
rect 586848 547718 586932 547954
rect 587168 547718 587200 547954
rect 586580 547634 587200 547718
rect 586580 547398 586612 547634
rect 586848 547398 586932 547634
rect 587168 547398 587200 547634
rect 586580 511954 587200 547398
rect 586580 511718 586612 511954
rect 586848 511718 586932 511954
rect 587168 511718 587200 511954
rect 586580 511634 587200 511718
rect 586580 511398 586612 511634
rect 586848 511398 586932 511634
rect 587168 511398 587200 511634
rect 586580 475954 587200 511398
rect 586580 475718 586612 475954
rect 586848 475718 586932 475954
rect 587168 475718 587200 475954
rect 586580 475634 587200 475718
rect 586580 475398 586612 475634
rect 586848 475398 586932 475634
rect 587168 475398 587200 475634
rect 586580 439954 587200 475398
rect 586580 439718 586612 439954
rect 586848 439718 586932 439954
rect 587168 439718 587200 439954
rect 586580 439634 587200 439718
rect 586580 439398 586612 439634
rect 586848 439398 586932 439634
rect 587168 439398 587200 439634
rect 586580 403954 587200 439398
rect 586580 403718 586612 403954
rect 586848 403718 586932 403954
rect 587168 403718 587200 403954
rect 586580 403634 587200 403718
rect 586580 403398 586612 403634
rect 586848 403398 586932 403634
rect 587168 403398 587200 403634
rect 586580 367954 587200 403398
rect 586580 367718 586612 367954
rect 586848 367718 586932 367954
rect 587168 367718 587200 367954
rect 586580 367634 587200 367718
rect 586580 367398 586612 367634
rect 586848 367398 586932 367634
rect 587168 367398 587200 367634
rect 586580 331954 587200 367398
rect 586580 331718 586612 331954
rect 586848 331718 586932 331954
rect 587168 331718 587200 331954
rect 586580 331634 587200 331718
rect 586580 331398 586612 331634
rect 586848 331398 586932 331634
rect 587168 331398 587200 331634
rect 586580 295954 587200 331398
rect 586580 295718 586612 295954
rect 586848 295718 586932 295954
rect 587168 295718 587200 295954
rect 586580 295634 587200 295718
rect 586580 295398 586612 295634
rect 586848 295398 586932 295634
rect 587168 295398 587200 295634
rect 586580 259954 587200 295398
rect 586580 259718 586612 259954
rect 586848 259718 586932 259954
rect 587168 259718 587200 259954
rect 586580 259634 587200 259718
rect 586580 259398 586612 259634
rect 586848 259398 586932 259634
rect 587168 259398 587200 259634
rect 586580 223954 587200 259398
rect 586580 223718 586612 223954
rect 586848 223718 586932 223954
rect 587168 223718 587200 223954
rect 586580 223634 587200 223718
rect 586580 223398 586612 223634
rect 586848 223398 586932 223634
rect 587168 223398 587200 223634
rect 586580 187954 587200 223398
rect 586580 187718 586612 187954
rect 586848 187718 586932 187954
rect 587168 187718 587200 187954
rect 586580 187634 587200 187718
rect 586580 187398 586612 187634
rect 586848 187398 586932 187634
rect 587168 187398 587200 187634
rect 586580 151954 587200 187398
rect 586580 151718 586612 151954
rect 586848 151718 586932 151954
rect 587168 151718 587200 151954
rect 586580 151634 587200 151718
rect 586580 151398 586612 151634
rect 586848 151398 586932 151634
rect 587168 151398 587200 151634
rect 586580 115954 587200 151398
rect 586580 115718 586612 115954
rect 586848 115718 586932 115954
rect 587168 115718 587200 115954
rect 586580 115634 587200 115718
rect 586580 115398 586612 115634
rect 586848 115398 586932 115634
rect 587168 115398 587200 115634
rect 586580 79954 587200 115398
rect 586580 79718 586612 79954
rect 586848 79718 586932 79954
rect 587168 79718 587200 79954
rect 586580 79634 587200 79718
rect 586580 79398 586612 79634
rect 586848 79398 586932 79634
rect 587168 79398 587200 79634
rect 586580 43954 587200 79398
rect 586580 43718 586612 43954
rect 586848 43718 586932 43954
rect 587168 43718 587200 43954
rect 586580 43634 587200 43718
rect 586580 43398 586612 43634
rect 586848 43398 586932 43634
rect 587168 43398 587200 43634
rect 586580 7954 587200 43398
rect 586580 7718 586612 7954
rect 586848 7718 586932 7954
rect 587168 7718 587200 7954
rect 586580 7634 587200 7718
rect 586580 7398 586612 7634
rect 586848 7398 586932 7634
rect 587168 7398 587200 7634
rect 582294 -1852 582326 -1616
rect 582562 -1852 582646 -1616
rect 582882 -1852 582914 -1616
rect 582294 -1936 582914 -1852
rect 582294 -2172 582326 -1936
rect 582562 -2172 582646 -1936
rect 582882 -2172 582914 -1936
rect 582294 -7964 582914 -2172
rect 586580 -1616 587200 7398
rect 586580 -1852 586612 -1616
rect 586848 -1852 586932 -1616
rect 587168 -1852 587200 -1616
rect 586580 -1936 587200 -1852
rect 586580 -2172 586612 -1936
rect 586848 -2172 586932 -1936
rect 587168 -2172 587200 -1936
rect 586580 -2204 587200 -2172
rect 587540 696454 588160 706512
rect 587540 696218 587572 696454
rect 587808 696218 587892 696454
rect 588128 696218 588160 696454
rect 587540 696134 588160 696218
rect 587540 695898 587572 696134
rect 587808 695898 587892 696134
rect 588128 695898 588160 696134
rect 587540 660454 588160 695898
rect 587540 660218 587572 660454
rect 587808 660218 587892 660454
rect 588128 660218 588160 660454
rect 587540 660134 588160 660218
rect 587540 659898 587572 660134
rect 587808 659898 587892 660134
rect 588128 659898 588160 660134
rect 587540 624454 588160 659898
rect 587540 624218 587572 624454
rect 587808 624218 587892 624454
rect 588128 624218 588160 624454
rect 587540 624134 588160 624218
rect 587540 623898 587572 624134
rect 587808 623898 587892 624134
rect 588128 623898 588160 624134
rect 587540 588454 588160 623898
rect 587540 588218 587572 588454
rect 587808 588218 587892 588454
rect 588128 588218 588160 588454
rect 587540 588134 588160 588218
rect 587540 587898 587572 588134
rect 587808 587898 587892 588134
rect 588128 587898 588160 588134
rect 587540 552454 588160 587898
rect 587540 552218 587572 552454
rect 587808 552218 587892 552454
rect 588128 552218 588160 552454
rect 587540 552134 588160 552218
rect 587540 551898 587572 552134
rect 587808 551898 587892 552134
rect 588128 551898 588160 552134
rect 587540 516454 588160 551898
rect 587540 516218 587572 516454
rect 587808 516218 587892 516454
rect 588128 516218 588160 516454
rect 587540 516134 588160 516218
rect 587540 515898 587572 516134
rect 587808 515898 587892 516134
rect 588128 515898 588160 516134
rect 587540 480454 588160 515898
rect 587540 480218 587572 480454
rect 587808 480218 587892 480454
rect 588128 480218 588160 480454
rect 587540 480134 588160 480218
rect 587540 479898 587572 480134
rect 587808 479898 587892 480134
rect 588128 479898 588160 480134
rect 587540 444454 588160 479898
rect 587540 444218 587572 444454
rect 587808 444218 587892 444454
rect 588128 444218 588160 444454
rect 587540 444134 588160 444218
rect 587540 443898 587572 444134
rect 587808 443898 587892 444134
rect 588128 443898 588160 444134
rect 587540 408454 588160 443898
rect 587540 408218 587572 408454
rect 587808 408218 587892 408454
rect 588128 408218 588160 408454
rect 587540 408134 588160 408218
rect 587540 407898 587572 408134
rect 587808 407898 587892 408134
rect 588128 407898 588160 408134
rect 587540 372454 588160 407898
rect 587540 372218 587572 372454
rect 587808 372218 587892 372454
rect 588128 372218 588160 372454
rect 587540 372134 588160 372218
rect 587540 371898 587572 372134
rect 587808 371898 587892 372134
rect 588128 371898 588160 372134
rect 587540 336454 588160 371898
rect 587540 336218 587572 336454
rect 587808 336218 587892 336454
rect 588128 336218 588160 336454
rect 587540 336134 588160 336218
rect 587540 335898 587572 336134
rect 587808 335898 587892 336134
rect 588128 335898 588160 336134
rect 587540 300454 588160 335898
rect 587540 300218 587572 300454
rect 587808 300218 587892 300454
rect 588128 300218 588160 300454
rect 587540 300134 588160 300218
rect 587540 299898 587572 300134
rect 587808 299898 587892 300134
rect 588128 299898 588160 300134
rect 587540 264454 588160 299898
rect 587540 264218 587572 264454
rect 587808 264218 587892 264454
rect 588128 264218 588160 264454
rect 587540 264134 588160 264218
rect 587540 263898 587572 264134
rect 587808 263898 587892 264134
rect 588128 263898 588160 264134
rect 587540 228454 588160 263898
rect 587540 228218 587572 228454
rect 587808 228218 587892 228454
rect 588128 228218 588160 228454
rect 587540 228134 588160 228218
rect 587540 227898 587572 228134
rect 587808 227898 587892 228134
rect 588128 227898 588160 228134
rect 587540 192454 588160 227898
rect 587540 192218 587572 192454
rect 587808 192218 587892 192454
rect 588128 192218 588160 192454
rect 587540 192134 588160 192218
rect 587540 191898 587572 192134
rect 587808 191898 587892 192134
rect 588128 191898 588160 192134
rect 587540 156454 588160 191898
rect 587540 156218 587572 156454
rect 587808 156218 587892 156454
rect 588128 156218 588160 156454
rect 587540 156134 588160 156218
rect 587540 155898 587572 156134
rect 587808 155898 587892 156134
rect 588128 155898 588160 156134
rect 587540 120454 588160 155898
rect 587540 120218 587572 120454
rect 587808 120218 587892 120454
rect 588128 120218 588160 120454
rect 587540 120134 588160 120218
rect 587540 119898 587572 120134
rect 587808 119898 587892 120134
rect 588128 119898 588160 120134
rect 587540 84454 588160 119898
rect 587540 84218 587572 84454
rect 587808 84218 587892 84454
rect 588128 84218 588160 84454
rect 587540 84134 588160 84218
rect 587540 83898 587572 84134
rect 587808 83898 587892 84134
rect 588128 83898 588160 84134
rect 587540 48454 588160 83898
rect 587540 48218 587572 48454
rect 587808 48218 587892 48454
rect 588128 48218 588160 48454
rect 587540 48134 588160 48218
rect 587540 47898 587572 48134
rect 587808 47898 587892 48134
rect 588128 47898 588160 48134
rect 587540 12454 588160 47898
rect 587540 12218 587572 12454
rect 587808 12218 587892 12454
rect 588128 12218 588160 12454
rect 587540 12134 588160 12218
rect 587540 11898 587572 12134
rect 587808 11898 587892 12134
rect 588128 11898 588160 12134
rect 587540 -2576 588160 11898
rect 587540 -2812 587572 -2576
rect 587808 -2812 587892 -2576
rect 588128 -2812 588160 -2576
rect 587540 -2896 588160 -2812
rect 587540 -3132 587572 -2896
rect 587808 -3132 587892 -2896
rect 588128 -3132 588160 -2896
rect 587540 -3164 588160 -3132
rect 588500 700954 589120 707472
rect 588500 700718 588532 700954
rect 588768 700718 588852 700954
rect 589088 700718 589120 700954
rect 588500 700634 589120 700718
rect 588500 700398 588532 700634
rect 588768 700398 588852 700634
rect 589088 700398 589120 700634
rect 588500 664954 589120 700398
rect 588500 664718 588532 664954
rect 588768 664718 588852 664954
rect 589088 664718 589120 664954
rect 588500 664634 589120 664718
rect 588500 664398 588532 664634
rect 588768 664398 588852 664634
rect 589088 664398 589120 664634
rect 588500 628954 589120 664398
rect 588500 628718 588532 628954
rect 588768 628718 588852 628954
rect 589088 628718 589120 628954
rect 588500 628634 589120 628718
rect 588500 628398 588532 628634
rect 588768 628398 588852 628634
rect 589088 628398 589120 628634
rect 588500 592954 589120 628398
rect 588500 592718 588532 592954
rect 588768 592718 588852 592954
rect 589088 592718 589120 592954
rect 588500 592634 589120 592718
rect 588500 592398 588532 592634
rect 588768 592398 588852 592634
rect 589088 592398 589120 592634
rect 588500 556954 589120 592398
rect 588500 556718 588532 556954
rect 588768 556718 588852 556954
rect 589088 556718 589120 556954
rect 588500 556634 589120 556718
rect 588500 556398 588532 556634
rect 588768 556398 588852 556634
rect 589088 556398 589120 556634
rect 588500 520954 589120 556398
rect 588500 520718 588532 520954
rect 588768 520718 588852 520954
rect 589088 520718 589120 520954
rect 588500 520634 589120 520718
rect 588500 520398 588532 520634
rect 588768 520398 588852 520634
rect 589088 520398 589120 520634
rect 588500 484954 589120 520398
rect 588500 484718 588532 484954
rect 588768 484718 588852 484954
rect 589088 484718 589120 484954
rect 588500 484634 589120 484718
rect 588500 484398 588532 484634
rect 588768 484398 588852 484634
rect 589088 484398 589120 484634
rect 588500 448954 589120 484398
rect 588500 448718 588532 448954
rect 588768 448718 588852 448954
rect 589088 448718 589120 448954
rect 588500 448634 589120 448718
rect 588500 448398 588532 448634
rect 588768 448398 588852 448634
rect 589088 448398 589120 448634
rect 588500 412954 589120 448398
rect 588500 412718 588532 412954
rect 588768 412718 588852 412954
rect 589088 412718 589120 412954
rect 588500 412634 589120 412718
rect 588500 412398 588532 412634
rect 588768 412398 588852 412634
rect 589088 412398 589120 412634
rect 588500 376954 589120 412398
rect 588500 376718 588532 376954
rect 588768 376718 588852 376954
rect 589088 376718 589120 376954
rect 588500 376634 589120 376718
rect 588500 376398 588532 376634
rect 588768 376398 588852 376634
rect 589088 376398 589120 376634
rect 588500 340954 589120 376398
rect 588500 340718 588532 340954
rect 588768 340718 588852 340954
rect 589088 340718 589120 340954
rect 588500 340634 589120 340718
rect 588500 340398 588532 340634
rect 588768 340398 588852 340634
rect 589088 340398 589120 340634
rect 588500 304954 589120 340398
rect 588500 304718 588532 304954
rect 588768 304718 588852 304954
rect 589088 304718 589120 304954
rect 588500 304634 589120 304718
rect 588500 304398 588532 304634
rect 588768 304398 588852 304634
rect 589088 304398 589120 304634
rect 588500 268954 589120 304398
rect 588500 268718 588532 268954
rect 588768 268718 588852 268954
rect 589088 268718 589120 268954
rect 588500 268634 589120 268718
rect 588500 268398 588532 268634
rect 588768 268398 588852 268634
rect 589088 268398 589120 268634
rect 588500 232954 589120 268398
rect 588500 232718 588532 232954
rect 588768 232718 588852 232954
rect 589088 232718 589120 232954
rect 588500 232634 589120 232718
rect 588500 232398 588532 232634
rect 588768 232398 588852 232634
rect 589088 232398 589120 232634
rect 588500 196954 589120 232398
rect 588500 196718 588532 196954
rect 588768 196718 588852 196954
rect 589088 196718 589120 196954
rect 588500 196634 589120 196718
rect 588500 196398 588532 196634
rect 588768 196398 588852 196634
rect 589088 196398 589120 196634
rect 588500 160954 589120 196398
rect 588500 160718 588532 160954
rect 588768 160718 588852 160954
rect 589088 160718 589120 160954
rect 588500 160634 589120 160718
rect 588500 160398 588532 160634
rect 588768 160398 588852 160634
rect 589088 160398 589120 160634
rect 588500 124954 589120 160398
rect 588500 124718 588532 124954
rect 588768 124718 588852 124954
rect 589088 124718 589120 124954
rect 588500 124634 589120 124718
rect 588500 124398 588532 124634
rect 588768 124398 588852 124634
rect 589088 124398 589120 124634
rect 588500 88954 589120 124398
rect 588500 88718 588532 88954
rect 588768 88718 588852 88954
rect 589088 88718 589120 88954
rect 588500 88634 589120 88718
rect 588500 88398 588532 88634
rect 588768 88398 588852 88634
rect 589088 88398 589120 88634
rect 588500 52954 589120 88398
rect 588500 52718 588532 52954
rect 588768 52718 588852 52954
rect 589088 52718 589120 52954
rect 588500 52634 589120 52718
rect 588500 52398 588532 52634
rect 588768 52398 588852 52634
rect 589088 52398 589120 52634
rect 588500 16954 589120 52398
rect 588500 16718 588532 16954
rect 588768 16718 588852 16954
rect 589088 16718 589120 16954
rect 588500 16634 589120 16718
rect 588500 16398 588532 16634
rect 588768 16398 588852 16634
rect 589088 16398 589120 16634
rect 588500 -3536 589120 16398
rect 588500 -3772 588532 -3536
rect 588768 -3772 588852 -3536
rect 589088 -3772 589120 -3536
rect 588500 -3856 589120 -3772
rect 588500 -4092 588532 -3856
rect 588768 -4092 588852 -3856
rect 589088 -4092 589120 -3856
rect 588500 -4124 589120 -4092
rect 589460 669454 590080 708432
rect 589460 669218 589492 669454
rect 589728 669218 589812 669454
rect 590048 669218 590080 669454
rect 589460 669134 590080 669218
rect 589460 668898 589492 669134
rect 589728 668898 589812 669134
rect 590048 668898 590080 669134
rect 589460 633454 590080 668898
rect 589460 633218 589492 633454
rect 589728 633218 589812 633454
rect 590048 633218 590080 633454
rect 589460 633134 590080 633218
rect 589460 632898 589492 633134
rect 589728 632898 589812 633134
rect 590048 632898 590080 633134
rect 589460 597454 590080 632898
rect 589460 597218 589492 597454
rect 589728 597218 589812 597454
rect 590048 597218 590080 597454
rect 589460 597134 590080 597218
rect 589460 596898 589492 597134
rect 589728 596898 589812 597134
rect 590048 596898 590080 597134
rect 589460 561454 590080 596898
rect 589460 561218 589492 561454
rect 589728 561218 589812 561454
rect 590048 561218 590080 561454
rect 589460 561134 590080 561218
rect 589460 560898 589492 561134
rect 589728 560898 589812 561134
rect 590048 560898 590080 561134
rect 589460 525454 590080 560898
rect 589460 525218 589492 525454
rect 589728 525218 589812 525454
rect 590048 525218 590080 525454
rect 589460 525134 590080 525218
rect 589460 524898 589492 525134
rect 589728 524898 589812 525134
rect 590048 524898 590080 525134
rect 589460 489454 590080 524898
rect 589460 489218 589492 489454
rect 589728 489218 589812 489454
rect 590048 489218 590080 489454
rect 589460 489134 590080 489218
rect 589460 488898 589492 489134
rect 589728 488898 589812 489134
rect 590048 488898 590080 489134
rect 589460 453454 590080 488898
rect 589460 453218 589492 453454
rect 589728 453218 589812 453454
rect 590048 453218 590080 453454
rect 589460 453134 590080 453218
rect 589460 452898 589492 453134
rect 589728 452898 589812 453134
rect 590048 452898 590080 453134
rect 589460 417454 590080 452898
rect 589460 417218 589492 417454
rect 589728 417218 589812 417454
rect 590048 417218 590080 417454
rect 589460 417134 590080 417218
rect 589460 416898 589492 417134
rect 589728 416898 589812 417134
rect 590048 416898 590080 417134
rect 589460 381454 590080 416898
rect 589460 381218 589492 381454
rect 589728 381218 589812 381454
rect 590048 381218 590080 381454
rect 589460 381134 590080 381218
rect 589460 380898 589492 381134
rect 589728 380898 589812 381134
rect 590048 380898 590080 381134
rect 589460 345454 590080 380898
rect 589460 345218 589492 345454
rect 589728 345218 589812 345454
rect 590048 345218 590080 345454
rect 589460 345134 590080 345218
rect 589460 344898 589492 345134
rect 589728 344898 589812 345134
rect 590048 344898 590080 345134
rect 589460 309454 590080 344898
rect 589460 309218 589492 309454
rect 589728 309218 589812 309454
rect 590048 309218 590080 309454
rect 589460 309134 590080 309218
rect 589460 308898 589492 309134
rect 589728 308898 589812 309134
rect 590048 308898 590080 309134
rect 589460 273454 590080 308898
rect 589460 273218 589492 273454
rect 589728 273218 589812 273454
rect 590048 273218 590080 273454
rect 589460 273134 590080 273218
rect 589460 272898 589492 273134
rect 589728 272898 589812 273134
rect 590048 272898 590080 273134
rect 589460 237454 590080 272898
rect 589460 237218 589492 237454
rect 589728 237218 589812 237454
rect 590048 237218 590080 237454
rect 589460 237134 590080 237218
rect 589460 236898 589492 237134
rect 589728 236898 589812 237134
rect 590048 236898 590080 237134
rect 589460 201454 590080 236898
rect 589460 201218 589492 201454
rect 589728 201218 589812 201454
rect 590048 201218 590080 201454
rect 589460 201134 590080 201218
rect 589460 200898 589492 201134
rect 589728 200898 589812 201134
rect 590048 200898 590080 201134
rect 589460 165454 590080 200898
rect 589460 165218 589492 165454
rect 589728 165218 589812 165454
rect 590048 165218 590080 165454
rect 589460 165134 590080 165218
rect 589460 164898 589492 165134
rect 589728 164898 589812 165134
rect 590048 164898 590080 165134
rect 589460 129454 590080 164898
rect 589460 129218 589492 129454
rect 589728 129218 589812 129454
rect 590048 129218 590080 129454
rect 589460 129134 590080 129218
rect 589460 128898 589492 129134
rect 589728 128898 589812 129134
rect 590048 128898 590080 129134
rect 589460 93454 590080 128898
rect 589460 93218 589492 93454
rect 589728 93218 589812 93454
rect 590048 93218 590080 93454
rect 589460 93134 590080 93218
rect 589460 92898 589492 93134
rect 589728 92898 589812 93134
rect 590048 92898 590080 93134
rect 589460 57454 590080 92898
rect 589460 57218 589492 57454
rect 589728 57218 589812 57454
rect 590048 57218 590080 57454
rect 589460 57134 590080 57218
rect 589460 56898 589492 57134
rect 589728 56898 589812 57134
rect 590048 56898 590080 57134
rect 589460 21454 590080 56898
rect 589460 21218 589492 21454
rect 589728 21218 589812 21454
rect 590048 21218 590080 21454
rect 589460 21134 590080 21218
rect 589460 20898 589492 21134
rect 589728 20898 589812 21134
rect 590048 20898 590080 21134
rect 589460 -4496 590080 20898
rect 589460 -4732 589492 -4496
rect 589728 -4732 589812 -4496
rect 590048 -4732 590080 -4496
rect 589460 -4816 590080 -4732
rect 589460 -5052 589492 -4816
rect 589728 -5052 589812 -4816
rect 590048 -5052 590080 -4816
rect 589460 -5084 590080 -5052
rect 590420 673954 591040 709392
rect 590420 673718 590452 673954
rect 590688 673718 590772 673954
rect 591008 673718 591040 673954
rect 590420 673634 591040 673718
rect 590420 673398 590452 673634
rect 590688 673398 590772 673634
rect 591008 673398 591040 673634
rect 590420 637954 591040 673398
rect 590420 637718 590452 637954
rect 590688 637718 590772 637954
rect 591008 637718 591040 637954
rect 590420 637634 591040 637718
rect 590420 637398 590452 637634
rect 590688 637398 590772 637634
rect 591008 637398 591040 637634
rect 590420 601954 591040 637398
rect 590420 601718 590452 601954
rect 590688 601718 590772 601954
rect 591008 601718 591040 601954
rect 590420 601634 591040 601718
rect 590420 601398 590452 601634
rect 590688 601398 590772 601634
rect 591008 601398 591040 601634
rect 590420 565954 591040 601398
rect 590420 565718 590452 565954
rect 590688 565718 590772 565954
rect 591008 565718 591040 565954
rect 590420 565634 591040 565718
rect 590420 565398 590452 565634
rect 590688 565398 590772 565634
rect 591008 565398 591040 565634
rect 590420 529954 591040 565398
rect 590420 529718 590452 529954
rect 590688 529718 590772 529954
rect 591008 529718 591040 529954
rect 590420 529634 591040 529718
rect 590420 529398 590452 529634
rect 590688 529398 590772 529634
rect 591008 529398 591040 529634
rect 590420 493954 591040 529398
rect 590420 493718 590452 493954
rect 590688 493718 590772 493954
rect 591008 493718 591040 493954
rect 590420 493634 591040 493718
rect 590420 493398 590452 493634
rect 590688 493398 590772 493634
rect 591008 493398 591040 493634
rect 590420 457954 591040 493398
rect 590420 457718 590452 457954
rect 590688 457718 590772 457954
rect 591008 457718 591040 457954
rect 590420 457634 591040 457718
rect 590420 457398 590452 457634
rect 590688 457398 590772 457634
rect 591008 457398 591040 457634
rect 590420 421954 591040 457398
rect 590420 421718 590452 421954
rect 590688 421718 590772 421954
rect 591008 421718 591040 421954
rect 590420 421634 591040 421718
rect 590420 421398 590452 421634
rect 590688 421398 590772 421634
rect 591008 421398 591040 421634
rect 590420 385954 591040 421398
rect 590420 385718 590452 385954
rect 590688 385718 590772 385954
rect 591008 385718 591040 385954
rect 590420 385634 591040 385718
rect 590420 385398 590452 385634
rect 590688 385398 590772 385634
rect 591008 385398 591040 385634
rect 590420 349954 591040 385398
rect 590420 349718 590452 349954
rect 590688 349718 590772 349954
rect 591008 349718 591040 349954
rect 590420 349634 591040 349718
rect 590420 349398 590452 349634
rect 590688 349398 590772 349634
rect 591008 349398 591040 349634
rect 590420 313954 591040 349398
rect 590420 313718 590452 313954
rect 590688 313718 590772 313954
rect 591008 313718 591040 313954
rect 590420 313634 591040 313718
rect 590420 313398 590452 313634
rect 590688 313398 590772 313634
rect 591008 313398 591040 313634
rect 590420 277954 591040 313398
rect 590420 277718 590452 277954
rect 590688 277718 590772 277954
rect 591008 277718 591040 277954
rect 590420 277634 591040 277718
rect 590420 277398 590452 277634
rect 590688 277398 590772 277634
rect 591008 277398 591040 277634
rect 590420 241954 591040 277398
rect 590420 241718 590452 241954
rect 590688 241718 590772 241954
rect 591008 241718 591040 241954
rect 590420 241634 591040 241718
rect 590420 241398 590452 241634
rect 590688 241398 590772 241634
rect 591008 241398 591040 241634
rect 590420 205954 591040 241398
rect 590420 205718 590452 205954
rect 590688 205718 590772 205954
rect 591008 205718 591040 205954
rect 590420 205634 591040 205718
rect 590420 205398 590452 205634
rect 590688 205398 590772 205634
rect 591008 205398 591040 205634
rect 590420 169954 591040 205398
rect 590420 169718 590452 169954
rect 590688 169718 590772 169954
rect 591008 169718 591040 169954
rect 590420 169634 591040 169718
rect 590420 169398 590452 169634
rect 590688 169398 590772 169634
rect 591008 169398 591040 169634
rect 590420 133954 591040 169398
rect 590420 133718 590452 133954
rect 590688 133718 590772 133954
rect 591008 133718 591040 133954
rect 590420 133634 591040 133718
rect 590420 133398 590452 133634
rect 590688 133398 590772 133634
rect 591008 133398 591040 133634
rect 590420 97954 591040 133398
rect 590420 97718 590452 97954
rect 590688 97718 590772 97954
rect 591008 97718 591040 97954
rect 590420 97634 591040 97718
rect 590420 97398 590452 97634
rect 590688 97398 590772 97634
rect 591008 97398 591040 97634
rect 590420 61954 591040 97398
rect 590420 61718 590452 61954
rect 590688 61718 590772 61954
rect 591008 61718 591040 61954
rect 590420 61634 591040 61718
rect 590420 61398 590452 61634
rect 590688 61398 590772 61634
rect 591008 61398 591040 61634
rect 590420 25954 591040 61398
rect 590420 25718 590452 25954
rect 590688 25718 590772 25954
rect 591008 25718 591040 25954
rect 590420 25634 591040 25718
rect 590420 25398 590452 25634
rect 590688 25398 590772 25634
rect 591008 25398 591040 25634
rect 590420 -5456 591040 25398
rect 590420 -5692 590452 -5456
rect 590688 -5692 590772 -5456
rect 591008 -5692 591040 -5456
rect 590420 -5776 591040 -5692
rect 590420 -6012 590452 -5776
rect 590688 -6012 590772 -5776
rect 591008 -6012 591040 -5776
rect 590420 -6044 591040 -6012
rect 591380 678454 592000 710352
rect 591380 678218 591412 678454
rect 591648 678218 591732 678454
rect 591968 678218 592000 678454
rect 591380 678134 592000 678218
rect 591380 677898 591412 678134
rect 591648 677898 591732 678134
rect 591968 677898 592000 678134
rect 591380 642454 592000 677898
rect 591380 642218 591412 642454
rect 591648 642218 591732 642454
rect 591968 642218 592000 642454
rect 591380 642134 592000 642218
rect 591380 641898 591412 642134
rect 591648 641898 591732 642134
rect 591968 641898 592000 642134
rect 591380 606454 592000 641898
rect 591380 606218 591412 606454
rect 591648 606218 591732 606454
rect 591968 606218 592000 606454
rect 591380 606134 592000 606218
rect 591380 605898 591412 606134
rect 591648 605898 591732 606134
rect 591968 605898 592000 606134
rect 591380 570454 592000 605898
rect 591380 570218 591412 570454
rect 591648 570218 591732 570454
rect 591968 570218 592000 570454
rect 591380 570134 592000 570218
rect 591380 569898 591412 570134
rect 591648 569898 591732 570134
rect 591968 569898 592000 570134
rect 591380 534454 592000 569898
rect 591380 534218 591412 534454
rect 591648 534218 591732 534454
rect 591968 534218 592000 534454
rect 591380 534134 592000 534218
rect 591380 533898 591412 534134
rect 591648 533898 591732 534134
rect 591968 533898 592000 534134
rect 591380 498454 592000 533898
rect 591380 498218 591412 498454
rect 591648 498218 591732 498454
rect 591968 498218 592000 498454
rect 591380 498134 592000 498218
rect 591380 497898 591412 498134
rect 591648 497898 591732 498134
rect 591968 497898 592000 498134
rect 591380 462454 592000 497898
rect 591380 462218 591412 462454
rect 591648 462218 591732 462454
rect 591968 462218 592000 462454
rect 591380 462134 592000 462218
rect 591380 461898 591412 462134
rect 591648 461898 591732 462134
rect 591968 461898 592000 462134
rect 591380 426454 592000 461898
rect 591380 426218 591412 426454
rect 591648 426218 591732 426454
rect 591968 426218 592000 426454
rect 591380 426134 592000 426218
rect 591380 425898 591412 426134
rect 591648 425898 591732 426134
rect 591968 425898 592000 426134
rect 591380 390454 592000 425898
rect 591380 390218 591412 390454
rect 591648 390218 591732 390454
rect 591968 390218 592000 390454
rect 591380 390134 592000 390218
rect 591380 389898 591412 390134
rect 591648 389898 591732 390134
rect 591968 389898 592000 390134
rect 591380 354454 592000 389898
rect 591380 354218 591412 354454
rect 591648 354218 591732 354454
rect 591968 354218 592000 354454
rect 591380 354134 592000 354218
rect 591380 353898 591412 354134
rect 591648 353898 591732 354134
rect 591968 353898 592000 354134
rect 591380 318454 592000 353898
rect 591380 318218 591412 318454
rect 591648 318218 591732 318454
rect 591968 318218 592000 318454
rect 591380 318134 592000 318218
rect 591380 317898 591412 318134
rect 591648 317898 591732 318134
rect 591968 317898 592000 318134
rect 591380 282454 592000 317898
rect 591380 282218 591412 282454
rect 591648 282218 591732 282454
rect 591968 282218 592000 282454
rect 591380 282134 592000 282218
rect 591380 281898 591412 282134
rect 591648 281898 591732 282134
rect 591968 281898 592000 282134
rect 591380 246454 592000 281898
rect 591380 246218 591412 246454
rect 591648 246218 591732 246454
rect 591968 246218 592000 246454
rect 591380 246134 592000 246218
rect 591380 245898 591412 246134
rect 591648 245898 591732 246134
rect 591968 245898 592000 246134
rect 591380 210454 592000 245898
rect 591380 210218 591412 210454
rect 591648 210218 591732 210454
rect 591968 210218 592000 210454
rect 591380 210134 592000 210218
rect 591380 209898 591412 210134
rect 591648 209898 591732 210134
rect 591968 209898 592000 210134
rect 591380 174454 592000 209898
rect 591380 174218 591412 174454
rect 591648 174218 591732 174454
rect 591968 174218 592000 174454
rect 591380 174134 592000 174218
rect 591380 173898 591412 174134
rect 591648 173898 591732 174134
rect 591968 173898 592000 174134
rect 591380 138454 592000 173898
rect 591380 138218 591412 138454
rect 591648 138218 591732 138454
rect 591968 138218 592000 138454
rect 591380 138134 592000 138218
rect 591380 137898 591412 138134
rect 591648 137898 591732 138134
rect 591968 137898 592000 138134
rect 591380 102454 592000 137898
rect 591380 102218 591412 102454
rect 591648 102218 591732 102454
rect 591968 102218 592000 102454
rect 591380 102134 592000 102218
rect 591380 101898 591412 102134
rect 591648 101898 591732 102134
rect 591968 101898 592000 102134
rect 591380 66454 592000 101898
rect 591380 66218 591412 66454
rect 591648 66218 591732 66454
rect 591968 66218 592000 66454
rect 591380 66134 592000 66218
rect 591380 65898 591412 66134
rect 591648 65898 591732 66134
rect 591968 65898 592000 66134
rect 591380 30454 592000 65898
rect 591380 30218 591412 30454
rect 591648 30218 591732 30454
rect 591968 30218 592000 30454
rect 591380 30134 592000 30218
rect 591380 29898 591412 30134
rect 591648 29898 591732 30134
rect 591968 29898 592000 30134
rect 591380 -6416 592000 29898
rect 591380 -6652 591412 -6416
rect 591648 -6652 591732 -6416
rect 591968 -6652 592000 -6416
rect 591380 -6736 592000 -6652
rect 591380 -6972 591412 -6736
rect 591648 -6972 591732 -6736
rect 591968 -6972 592000 -6736
rect 591380 -7004 592000 -6972
rect 592340 682954 592960 711312
rect 592340 682718 592372 682954
rect 592608 682718 592692 682954
rect 592928 682718 592960 682954
rect 592340 682634 592960 682718
rect 592340 682398 592372 682634
rect 592608 682398 592692 682634
rect 592928 682398 592960 682634
rect 592340 646954 592960 682398
rect 592340 646718 592372 646954
rect 592608 646718 592692 646954
rect 592928 646718 592960 646954
rect 592340 646634 592960 646718
rect 592340 646398 592372 646634
rect 592608 646398 592692 646634
rect 592928 646398 592960 646634
rect 592340 610954 592960 646398
rect 592340 610718 592372 610954
rect 592608 610718 592692 610954
rect 592928 610718 592960 610954
rect 592340 610634 592960 610718
rect 592340 610398 592372 610634
rect 592608 610398 592692 610634
rect 592928 610398 592960 610634
rect 592340 574954 592960 610398
rect 592340 574718 592372 574954
rect 592608 574718 592692 574954
rect 592928 574718 592960 574954
rect 592340 574634 592960 574718
rect 592340 574398 592372 574634
rect 592608 574398 592692 574634
rect 592928 574398 592960 574634
rect 592340 538954 592960 574398
rect 592340 538718 592372 538954
rect 592608 538718 592692 538954
rect 592928 538718 592960 538954
rect 592340 538634 592960 538718
rect 592340 538398 592372 538634
rect 592608 538398 592692 538634
rect 592928 538398 592960 538634
rect 592340 502954 592960 538398
rect 592340 502718 592372 502954
rect 592608 502718 592692 502954
rect 592928 502718 592960 502954
rect 592340 502634 592960 502718
rect 592340 502398 592372 502634
rect 592608 502398 592692 502634
rect 592928 502398 592960 502634
rect 592340 466954 592960 502398
rect 592340 466718 592372 466954
rect 592608 466718 592692 466954
rect 592928 466718 592960 466954
rect 592340 466634 592960 466718
rect 592340 466398 592372 466634
rect 592608 466398 592692 466634
rect 592928 466398 592960 466634
rect 592340 430954 592960 466398
rect 592340 430718 592372 430954
rect 592608 430718 592692 430954
rect 592928 430718 592960 430954
rect 592340 430634 592960 430718
rect 592340 430398 592372 430634
rect 592608 430398 592692 430634
rect 592928 430398 592960 430634
rect 592340 394954 592960 430398
rect 592340 394718 592372 394954
rect 592608 394718 592692 394954
rect 592928 394718 592960 394954
rect 592340 394634 592960 394718
rect 592340 394398 592372 394634
rect 592608 394398 592692 394634
rect 592928 394398 592960 394634
rect 592340 358954 592960 394398
rect 592340 358718 592372 358954
rect 592608 358718 592692 358954
rect 592928 358718 592960 358954
rect 592340 358634 592960 358718
rect 592340 358398 592372 358634
rect 592608 358398 592692 358634
rect 592928 358398 592960 358634
rect 592340 322954 592960 358398
rect 592340 322718 592372 322954
rect 592608 322718 592692 322954
rect 592928 322718 592960 322954
rect 592340 322634 592960 322718
rect 592340 322398 592372 322634
rect 592608 322398 592692 322634
rect 592928 322398 592960 322634
rect 592340 286954 592960 322398
rect 592340 286718 592372 286954
rect 592608 286718 592692 286954
rect 592928 286718 592960 286954
rect 592340 286634 592960 286718
rect 592340 286398 592372 286634
rect 592608 286398 592692 286634
rect 592928 286398 592960 286634
rect 592340 250954 592960 286398
rect 592340 250718 592372 250954
rect 592608 250718 592692 250954
rect 592928 250718 592960 250954
rect 592340 250634 592960 250718
rect 592340 250398 592372 250634
rect 592608 250398 592692 250634
rect 592928 250398 592960 250634
rect 592340 214954 592960 250398
rect 592340 214718 592372 214954
rect 592608 214718 592692 214954
rect 592928 214718 592960 214954
rect 592340 214634 592960 214718
rect 592340 214398 592372 214634
rect 592608 214398 592692 214634
rect 592928 214398 592960 214634
rect 592340 178954 592960 214398
rect 592340 178718 592372 178954
rect 592608 178718 592692 178954
rect 592928 178718 592960 178954
rect 592340 178634 592960 178718
rect 592340 178398 592372 178634
rect 592608 178398 592692 178634
rect 592928 178398 592960 178634
rect 592340 142954 592960 178398
rect 592340 142718 592372 142954
rect 592608 142718 592692 142954
rect 592928 142718 592960 142954
rect 592340 142634 592960 142718
rect 592340 142398 592372 142634
rect 592608 142398 592692 142634
rect 592928 142398 592960 142634
rect 592340 106954 592960 142398
rect 592340 106718 592372 106954
rect 592608 106718 592692 106954
rect 592928 106718 592960 106954
rect 592340 106634 592960 106718
rect 592340 106398 592372 106634
rect 592608 106398 592692 106634
rect 592928 106398 592960 106634
rect 592340 70954 592960 106398
rect 592340 70718 592372 70954
rect 592608 70718 592692 70954
rect 592928 70718 592960 70954
rect 592340 70634 592960 70718
rect 592340 70398 592372 70634
rect 592608 70398 592692 70634
rect 592928 70398 592960 70634
rect 592340 34954 592960 70398
rect 592340 34718 592372 34954
rect 592608 34718 592692 34954
rect 592928 34718 592960 34954
rect 592340 34634 592960 34718
rect 592340 34398 592372 34634
rect 592608 34398 592692 34634
rect 592928 34398 592960 34634
rect 592340 -7376 592960 34398
rect 592340 -7612 592372 -7376
rect 592608 -7612 592692 -7376
rect 592928 -7612 592960 -7376
rect 592340 -7696 592960 -7612
rect 592340 -7932 592372 -7696
rect 592608 -7932 592692 -7696
rect 592928 -7932 592960 -7696
rect 592340 -7964 592960 -7932
<< via4 >>
rect -9004 711632 -8768 711868
rect -8684 711632 -8448 711868
rect -9004 711312 -8768 711548
rect -8684 711312 -8448 711548
rect -9004 682718 -8768 682954
rect -8684 682718 -8448 682954
rect -9004 682398 -8768 682634
rect -8684 682398 -8448 682634
rect -9004 646718 -8768 646954
rect -8684 646718 -8448 646954
rect -9004 646398 -8768 646634
rect -8684 646398 -8448 646634
rect -9004 610718 -8768 610954
rect -8684 610718 -8448 610954
rect -9004 610398 -8768 610634
rect -8684 610398 -8448 610634
rect -9004 574718 -8768 574954
rect -8684 574718 -8448 574954
rect -9004 574398 -8768 574634
rect -8684 574398 -8448 574634
rect -9004 538718 -8768 538954
rect -8684 538718 -8448 538954
rect -9004 538398 -8768 538634
rect -8684 538398 -8448 538634
rect -9004 502718 -8768 502954
rect -8684 502718 -8448 502954
rect -9004 502398 -8768 502634
rect -8684 502398 -8448 502634
rect -9004 466718 -8768 466954
rect -8684 466718 -8448 466954
rect -9004 466398 -8768 466634
rect -8684 466398 -8448 466634
rect -9004 430718 -8768 430954
rect -8684 430718 -8448 430954
rect -9004 430398 -8768 430634
rect -8684 430398 -8448 430634
rect -9004 394718 -8768 394954
rect -8684 394718 -8448 394954
rect -9004 394398 -8768 394634
rect -8684 394398 -8448 394634
rect -9004 358718 -8768 358954
rect -8684 358718 -8448 358954
rect -9004 358398 -8768 358634
rect -8684 358398 -8448 358634
rect -9004 322718 -8768 322954
rect -8684 322718 -8448 322954
rect -9004 322398 -8768 322634
rect -8684 322398 -8448 322634
rect -9004 286718 -8768 286954
rect -8684 286718 -8448 286954
rect -9004 286398 -8768 286634
rect -8684 286398 -8448 286634
rect -9004 250718 -8768 250954
rect -8684 250718 -8448 250954
rect -9004 250398 -8768 250634
rect -8684 250398 -8448 250634
rect -9004 214718 -8768 214954
rect -8684 214718 -8448 214954
rect -9004 214398 -8768 214634
rect -8684 214398 -8448 214634
rect -9004 178718 -8768 178954
rect -8684 178718 -8448 178954
rect -9004 178398 -8768 178634
rect -8684 178398 -8448 178634
rect -9004 142718 -8768 142954
rect -8684 142718 -8448 142954
rect -9004 142398 -8768 142634
rect -8684 142398 -8448 142634
rect -9004 106718 -8768 106954
rect -8684 106718 -8448 106954
rect -9004 106398 -8768 106634
rect -8684 106398 -8448 106634
rect -9004 70718 -8768 70954
rect -8684 70718 -8448 70954
rect -9004 70398 -8768 70634
rect -8684 70398 -8448 70634
rect -9004 34718 -8768 34954
rect -8684 34718 -8448 34954
rect -9004 34398 -8768 34634
rect -8684 34398 -8448 34634
rect -8044 710672 -7808 710908
rect -7724 710672 -7488 710908
rect -8044 710352 -7808 710588
rect -7724 710352 -7488 710588
rect -8044 678218 -7808 678454
rect -7724 678218 -7488 678454
rect -8044 677898 -7808 678134
rect -7724 677898 -7488 678134
rect -8044 642218 -7808 642454
rect -7724 642218 -7488 642454
rect -8044 641898 -7808 642134
rect -7724 641898 -7488 642134
rect -8044 606218 -7808 606454
rect -7724 606218 -7488 606454
rect -8044 605898 -7808 606134
rect -7724 605898 -7488 606134
rect -8044 570218 -7808 570454
rect -7724 570218 -7488 570454
rect -8044 569898 -7808 570134
rect -7724 569898 -7488 570134
rect -8044 534218 -7808 534454
rect -7724 534218 -7488 534454
rect -8044 533898 -7808 534134
rect -7724 533898 -7488 534134
rect -8044 498218 -7808 498454
rect -7724 498218 -7488 498454
rect -8044 497898 -7808 498134
rect -7724 497898 -7488 498134
rect -8044 462218 -7808 462454
rect -7724 462218 -7488 462454
rect -8044 461898 -7808 462134
rect -7724 461898 -7488 462134
rect -8044 426218 -7808 426454
rect -7724 426218 -7488 426454
rect -8044 425898 -7808 426134
rect -7724 425898 -7488 426134
rect -8044 390218 -7808 390454
rect -7724 390218 -7488 390454
rect -8044 389898 -7808 390134
rect -7724 389898 -7488 390134
rect -8044 354218 -7808 354454
rect -7724 354218 -7488 354454
rect -8044 353898 -7808 354134
rect -7724 353898 -7488 354134
rect -8044 318218 -7808 318454
rect -7724 318218 -7488 318454
rect -8044 317898 -7808 318134
rect -7724 317898 -7488 318134
rect -8044 282218 -7808 282454
rect -7724 282218 -7488 282454
rect -8044 281898 -7808 282134
rect -7724 281898 -7488 282134
rect -8044 246218 -7808 246454
rect -7724 246218 -7488 246454
rect -8044 245898 -7808 246134
rect -7724 245898 -7488 246134
rect -8044 210218 -7808 210454
rect -7724 210218 -7488 210454
rect -8044 209898 -7808 210134
rect -7724 209898 -7488 210134
rect -8044 174218 -7808 174454
rect -7724 174218 -7488 174454
rect -8044 173898 -7808 174134
rect -7724 173898 -7488 174134
rect -8044 138218 -7808 138454
rect -7724 138218 -7488 138454
rect -8044 137898 -7808 138134
rect -7724 137898 -7488 138134
rect -8044 102218 -7808 102454
rect -7724 102218 -7488 102454
rect -8044 101898 -7808 102134
rect -7724 101898 -7488 102134
rect -8044 66218 -7808 66454
rect -7724 66218 -7488 66454
rect -8044 65898 -7808 66134
rect -7724 65898 -7488 66134
rect -8044 30218 -7808 30454
rect -7724 30218 -7488 30454
rect -8044 29898 -7808 30134
rect -7724 29898 -7488 30134
rect -7084 709712 -6848 709948
rect -6764 709712 -6528 709948
rect -7084 709392 -6848 709628
rect -6764 709392 -6528 709628
rect -7084 673718 -6848 673954
rect -6764 673718 -6528 673954
rect -7084 673398 -6848 673634
rect -6764 673398 -6528 673634
rect -7084 637718 -6848 637954
rect -6764 637718 -6528 637954
rect -7084 637398 -6848 637634
rect -6764 637398 -6528 637634
rect -7084 601718 -6848 601954
rect -6764 601718 -6528 601954
rect -7084 601398 -6848 601634
rect -6764 601398 -6528 601634
rect -7084 565718 -6848 565954
rect -6764 565718 -6528 565954
rect -7084 565398 -6848 565634
rect -6764 565398 -6528 565634
rect -7084 529718 -6848 529954
rect -6764 529718 -6528 529954
rect -7084 529398 -6848 529634
rect -6764 529398 -6528 529634
rect -7084 493718 -6848 493954
rect -6764 493718 -6528 493954
rect -7084 493398 -6848 493634
rect -6764 493398 -6528 493634
rect -7084 457718 -6848 457954
rect -6764 457718 -6528 457954
rect -7084 457398 -6848 457634
rect -6764 457398 -6528 457634
rect -7084 421718 -6848 421954
rect -6764 421718 -6528 421954
rect -7084 421398 -6848 421634
rect -6764 421398 -6528 421634
rect -7084 385718 -6848 385954
rect -6764 385718 -6528 385954
rect -7084 385398 -6848 385634
rect -6764 385398 -6528 385634
rect -7084 349718 -6848 349954
rect -6764 349718 -6528 349954
rect -7084 349398 -6848 349634
rect -6764 349398 -6528 349634
rect -7084 313718 -6848 313954
rect -6764 313718 -6528 313954
rect -7084 313398 -6848 313634
rect -6764 313398 -6528 313634
rect -7084 277718 -6848 277954
rect -6764 277718 -6528 277954
rect -7084 277398 -6848 277634
rect -6764 277398 -6528 277634
rect -7084 241718 -6848 241954
rect -6764 241718 -6528 241954
rect -7084 241398 -6848 241634
rect -6764 241398 -6528 241634
rect -7084 205718 -6848 205954
rect -6764 205718 -6528 205954
rect -7084 205398 -6848 205634
rect -6764 205398 -6528 205634
rect -7084 169718 -6848 169954
rect -6764 169718 -6528 169954
rect -7084 169398 -6848 169634
rect -6764 169398 -6528 169634
rect -7084 133718 -6848 133954
rect -6764 133718 -6528 133954
rect -7084 133398 -6848 133634
rect -6764 133398 -6528 133634
rect -7084 97718 -6848 97954
rect -6764 97718 -6528 97954
rect -7084 97398 -6848 97634
rect -6764 97398 -6528 97634
rect -7084 61718 -6848 61954
rect -6764 61718 -6528 61954
rect -7084 61398 -6848 61634
rect -6764 61398 -6528 61634
rect -7084 25718 -6848 25954
rect -6764 25718 -6528 25954
rect -7084 25398 -6848 25634
rect -6764 25398 -6528 25634
rect -6124 708752 -5888 708988
rect -5804 708752 -5568 708988
rect -6124 708432 -5888 708668
rect -5804 708432 -5568 708668
rect -6124 669218 -5888 669454
rect -5804 669218 -5568 669454
rect -6124 668898 -5888 669134
rect -5804 668898 -5568 669134
rect -6124 633218 -5888 633454
rect -5804 633218 -5568 633454
rect -6124 632898 -5888 633134
rect -5804 632898 -5568 633134
rect -6124 597218 -5888 597454
rect -5804 597218 -5568 597454
rect -6124 596898 -5888 597134
rect -5804 596898 -5568 597134
rect -6124 561218 -5888 561454
rect -5804 561218 -5568 561454
rect -6124 560898 -5888 561134
rect -5804 560898 -5568 561134
rect -6124 525218 -5888 525454
rect -5804 525218 -5568 525454
rect -6124 524898 -5888 525134
rect -5804 524898 -5568 525134
rect -6124 489218 -5888 489454
rect -5804 489218 -5568 489454
rect -6124 488898 -5888 489134
rect -5804 488898 -5568 489134
rect -6124 453218 -5888 453454
rect -5804 453218 -5568 453454
rect -6124 452898 -5888 453134
rect -5804 452898 -5568 453134
rect -6124 417218 -5888 417454
rect -5804 417218 -5568 417454
rect -6124 416898 -5888 417134
rect -5804 416898 -5568 417134
rect -6124 381218 -5888 381454
rect -5804 381218 -5568 381454
rect -6124 380898 -5888 381134
rect -5804 380898 -5568 381134
rect -6124 345218 -5888 345454
rect -5804 345218 -5568 345454
rect -6124 344898 -5888 345134
rect -5804 344898 -5568 345134
rect -6124 309218 -5888 309454
rect -5804 309218 -5568 309454
rect -6124 308898 -5888 309134
rect -5804 308898 -5568 309134
rect -6124 273218 -5888 273454
rect -5804 273218 -5568 273454
rect -6124 272898 -5888 273134
rect -5804 272898 -5568 273134
rect -6124 237218 -5888 237454
rect -5804 237218 -5568 237454
rect -6124 236898 -5888 237134
rect -5804 236898 -5568 237134
rect -6124 201218 -5888 201454
rect -5804 201218 -5568 201454
rect -6124 200898 -5888 201134
rect -5804 200898 -5568 201134
rect -6124 165218 -5888 165454
rect -5804 165218 -5568 165454
rect -6124 164898 -5888 165134
rect -5804 164898 -5568 165134
rect -6124 129218 -5888 129454
rect -5804 129218 -5568 129454
rect -6124 128898 -5888 129134
rect -5804 128898 -5568 129134
rect -6124 93218 -5888 93454
rect -5804 93218 -5568 93454
rect -6124 92898 -5888 93134
rect -5804 92898 -5568 93134
rect -6124 57218 -5888 57454
rect -5804 57218 -5568 57454
rect -6124 56898 -5888 57134
rect -5804 56898 -5568 57134
rect -6124 21218 -5888 21454
rect -5804 21218 -5568 21454
rect -6124 20898 -5888 21134
rect -5804 20898 -5568 21134
rect -5164 707792 -4928 708028
rect -4844 707792 -4608 708028
rect -5164 707472 -4928 707708
rect -4844 707472 -4608 707708
rect -5164 700718 -4928 700954
rect -4844 700718 -4608 700954
rect -5164 700398 -4928 700634
rect -4844 700398 -4608 700634
rect -5164 664718 -4928 664954
rect -4844 664718 -4608 664954
rect -5164 664398 -4928 664634
rect -4844 664398 -4608 664634
rect -5164 628718 -4928 628954
rect -4844 628718 -4608 628954
rect -5164 628398 -4928 628634
rect -4844 628398 -4608 628634
rect -5164 592718 -4928 592954
rect -4844 592718 -4608 592954
rect -5164 592398 -4928 592634
rect -4844 592398 -4608 592634
rect -5164 556718 -4928 556954
rect -4844 556718 -4608 556954
rect -5164 556398 -4928 556634
rect -4844 556398 -4608 556634
rect -5164 520718 -4928 520954
rect -4844 520718 -4608 520954
rect -5164 520398 -4928 520634
rect -4844 520398 -4608 520634
rect -5164 484718 -4928 484954
rect -4844 484718 -4608 484954
rect -5164 484398 -4928 484634
rect -4844 484398 -4608 484634
rect -5164 448718 -4928 448954
rect -4844 448718 -4608 448954
rect -5164 448398 -4928 448634
rect -4844 448398 -4608 448634
rect -5164 412718 -4928 412954
rect -4844 412718 -4608 412954
rect -5164 412398 -4928 412634
rect -4844 412398 -4608 412634
rect -5164 376718 -4928 376954
rect -4844 376718 -4608 376954
rect -5164 376398 -4928 376634
rect -4844 376398 -4608 376634
rect -5164 340718 -4928 340954
rect -4844 340718 -4608 340954
rect -5164 340398 -4928 340634
rect -4844 340398 -4608 340634
rect -5164 304718 -4928 304954
rect -4844 304718 -4608 304954
rect -5164 304398 -4928 304634
rect -4844 304398 -4608 304634
rect -5164 268718 -4928 268954
rect -4844 268718 -4608 268954
rect -5164 268398 -4928 268634
rect -4844 268398 -4608 268634
rect -5164 232718 -4928 232954
rect -4844 232718 -4608 232954
rect -5164 232398 -4928 232634
rect -4844 232398 -4608 232634
rect -5164 196718 -4928 196954
rect -4844 196718 -4608 196954
rect -5164 196398 -4928 196634
rect -4844 196398 -4608 196634
rect -5164 160718 -4928 160954
rect -4844 160718 -4608 160954
rect -5164 160398 -4928 160634
rect -4844 160398 -4608 160634
rect -5164 124718 -4928 124954
rect -4844 124718 -4608 124954
rect -5164 124398 -4928 124634
rect -4844 124398 -4608 124634
rect -5164 88718 -4928 88954
rect -4844 88718 -4608 88954
rect -5164 88398 -4928 88634
rect -4844 88398 -4608 88634
rect -5164 52718 -4928 52954
rect -4844 52718 -4608 52954
rect -5164 52398 -4928 52634
rect -4844 52398 -4608 52634
rect -5164 16718 -4928 16954
rect -4844 16718 -4608 16954
rect -5164 16398 -4928 16634
rect -4844 16398 -4608 16634
rect -4204 706832 -3968 707068
rect -3884 706832 -3648 707068
rect -4204 706512 -3968 706748
rect -3884 706512 -3648 706748
rect -4204 696218 -3968 696454
rect -3884 696218 -3648 696454
rect -4204 695898 -3968 696134
rect -3884 695898 -3648 696134
rect -4204 660218 -3968 660454
rect -3884 660218 -3648 660454
rect -4204 659898 -3968 660134
rect -3884 659898 -3648 660134
rect -4204 624218 -3968 624454
rect -3884 624218 -3648 624454
rect -4204 623898 -3968 624134
rect -3884 623898 -3648 624134
rect -4204 588218 -3968 588454
rect -3884 588218 -3648 588454
rect -4204 587898 -3968 588134
rect -3884 587898 -3648 588134
rect -4204 552218 -3968 552454
rect -3884 552218 -3648 552454
rect -4204 551898 -3968 552134
rect -3884 551898 -3648 552134
rect -4204 516218 -3968 516454
rect -3884 516218 -3648 516454
rect -4204 515898 -3968 516134
rect -3884 515898 -3648 516134
rect -4204 480218 -3968 480454
rect -3884 480218 -3648 480454
rect -4204 479898 -3968 480134
rect -3884 479898 -3648 480134
rect -4204 444218 -3968 444454
rect -3884 444218 -3648 444454
rect -4204 443898 -3968 444134
rect -3884 443898 -3648 444134
rect -4204 408218 -3968 408454
rect -3884 408218 -3648 408454
rect -4204 407898 -3968 408134
rect -3884 407898 -3648 408134
rect -4204 372218 -3968 372454
rect -3884 372218 -3648 372454
rect -4204 371898 -3968 372134
rect -3884 371898 -3648 372134
rect -4204 336218 -3968 336454
rect -3884 336218 -3648 336454
rect -4204 335898 -3968 336134
rect -3884 335898 -3648 336134
rect -4204 300218 -3968 300454
rect -3884 300218 -3648 300454
rect -4204 299898 -3968 300134
rect -3884 299898 -3648 300134
rect -4204 264218 -3968 264454
rect -3884 264218 -3648 264454
rect -4204 263898 -3968 264134
rect -3884 263898 -3648 264134
rect -4204 228218 -3968 228454
rect -3884 228218 -3648 228454
rect -4204 227898 -3968 228134
rect -3884 227898 -3648 228134
rect -4204 192218 -3968 192454
rect -3884 192218 -3648 192454
rect -4204 191898 -3968 192134
rect -3884 191898 -3648 192134
rect -4204 156218 -3968 156454
rect -3884 156218 -3648 156454
rect -4204 155898 -3968 156134
rect -3884 155898 -3648 156134
rect -4204 120218 -3968 120454
rect -3884 120218 -3648 120454
rect -4204 119898 -3968 120134
rect -3884 119898 -3648 120134
rect -4204 84218 -3968 84454
rect -3884 84218 -3648 84454
rect -4204 83898 -3968 84134
rect -3884 83898 -3648 84134
rect -4204 48218 -3968 48454
rect -3884 48218 -3648 48454
rect -4204 47898 -3968 48134
rect -3884 47898 -3648 48134
rect -4204 12218 -3968 12454
rect -3884 12218 -3648 12454
rect -4204 11898 -3968 12134
rect -3884 11898 -3648 12134
rect -3244 705872 -3008 706108
rect -2924 705872 -2688 706108
rect -3244 705552 -3008 705788
rect -2924 705552 -2688 705788
rect -3244 691718 -3008 691954
rect -2924 691718 -2688 691954
rect -3244 691398 -3008 691634
rect -2924 691398 -2688 691634
rect -3244 655718 -3008 655954
rect -2924 655718 -2688 655954
rect -3244 655398 -3008 655634
rect -2924 655398 -2688 655634
rect -3244 619718 -3008 619954
rect -2924 619718 -2688 619954
rect -3244 619398 -3008 619634
rect -2924 619398 -2688 619634
rect -3244 583718 -3008 583954
rect -2924 583718 -2688 583954
rect -3244 583398 -3008 583634
rect -2924 583398 -2688 583634
rect -3244 547718 -3008 547954
rect -2924 547718 -2688 547954
rect -3244 547398 -3008 547634
rect -2924 547398 -2688 547634
rect -3244 511718 -3008 511954
rect -2924 511718 -2688 511954
rect -3244 511398 -3008 511634
rect -2924 511398 -2688 511634
rect -3244 475718 -3008 475954
rect -2924 475718 -2688 475954
rect -3244 475398 -3008 475634
rect -2924 475398 -2688 475634
rect -3244 439718 -3008 439954
rect -2924 439718 -2688 439954
rect -3244 439398 -3008 439634
rect -2924 439398 -2688 439634
rect -3244 403718 -3008 403954
rect -2924 403718 -2688 403954
rect -3244 403398 -3008 403634
rect -2924 403398 -2688 403634
rect -3244 367718 -3008 367954
rect -2924 367718 -2688 367954
rect -3244 367398 -3008 367634
rect -2924 367398 -2688 367634
rect -3244 331718 -3008 331954
rect -2924 331718 -2688 331954
rect -3244 331398 -3008 331634
rect -2924 331398 -2688 331634
rect -3244 295718 -3008 295954
rect -2924 295718 -2688 295954
rect -3244 295398 -3008 295634
rect -2924 295398 -2688 295634
rect -3244 259718 -3008 259954
rect -2924 259718 -2688 259954
rect -3244 259398 -3008 259634
rect -2924 259398 -2688 259634
rect -3244 223718 -3008 223954
rect -2924 223718 -2688 223954
rect -3244 223398 -3008 223634
rect -2924 223398 -2688 223634
rect -3244 187718 -3008 187954
rect -2924 187718 -2688 187954
rect -3244 187398 -3008 187634
rect -2924 187398 -2688 187634
rect -3244 151718 -3008 151954
rect -2924 151718 -2688 151954
rect -3244 151398 -3008 151634
rect -2924 151398 -2688 151634
rect -3244 115718 -3008 115954
rect -2924 115718 -2688 115954
rect -3244 115398 -3008 115634
rect -2924 115398 -2688 115634
rect -3244 79718 -3008 79954
rect -2924 79718 -2688 79954
rect -3244 79398 -3008 79634
rect -2924 79398 -2688 79634
rect -3244 43718 -3008 43954
rect -2924 43718 -2688 43954
rect -3244 43398 -3008 43634
rect -2924 43398 -2688 43634
rect -3244 7718 -3008 7954
rect -2924 7718 -2688 7954
rect -3244 7398 -3008 7634
rect -2924 7398 -2688 7634
rect -2284 704912 -2048 705148
rect -1964 704912 -1728 705148
rect -2284 704592 -2048 704828
rect -1964 704592 -1728 704828
rect -2284 687218 -2048 687454
rect -1964 687218 -1728 687454
rect -2284 686898 -2048 687134
rect -1964 686898 -1728 687134
rect -2284 651218 -2048 651454
rect -1964 651218 -1728 651454
rect -2284 650898 -2048 651134
rect -1964 650898 -1728 651134
rect -2284 615218 -2048 615454
rect -1964 615218 -1728 615454
rect -2284 614898 -2048 615134
rect -1964 614898 -1728 615134
rect -2284 579218 -2048 579454
rect -1964 579218 -1728 579454
rect -2284 578898 -2048 579134
rect -1964 578898 -1728 579134
rect -2284 543218 -2048 543454
rect -1964 543218 -1728 543454
rect -2284 542898 -2048 543134
rect -1964 542898 -1728 543134
rect -2284 507218 -2048 507454
rect -1964 507218 -1728 507454
rect -2284 506898 -2048 507134
rect -1964 506898 -1728 507134
rect -2284 471218 -2048 471454
rect -1964 471218 -1728 471454
rect -2284 470898 -2048 471134
rect -1964 470898 -1728 471134
rect -2284 435218 -2048 435454
rect -1964 435218 -1728 435454
rect -2284 434898 -2048 435134
rect -1964 434898 -1728 435134
rect -2284 399218 -2048 399454
rect -1964 399218 -1728 399454
rect -2284 398898 -2048 399134
rect -1964 398898 -1728 399134
rect -2284 363218 -2048 363454
rect -1964 363218 -1728 363454
rect -2284 362898 -2048 363134
rect -1964 362898 -1728 363134
rect -2284 327218 -2048 327454
rect -1964 327218 -1728 327454
rect -2284 326898 -2048 327134
rect -1964 326898 -1728 327134
rect -2284 291218 -2048 291454
rect -1964 291218 -1728 291454
rect -2284 290898 -2048 291134
rect -1964 290898 -1728 291134
rect -2284 255218 -2048 255454
rect -1964 255218 -1728 255454
rect -2284 254898 -2048 255134
rect -1964 254898 -1728 255134
rect -2284 219218 -2048 219454
rect -1964 219218 -1728 219454
rect -2284 218898 -2048 219134
rect -1964 218898 -1728 219134
rect -2284 183218 -2048 183454
rect -1964 183218 -1728 183454
rect -2284 182898 -2048 183134
rect -1964 182898 -1728 183134
rect -2284 147218 -2048 147454
rect -1964 147218 -1728 147454
rect -2284 146898 -2048 147134
rect -1964 146898 -1728 147134
rect -2284 111218 -2048 111454
rect -1964 111218 -1728 111454
rect -2284 110898 -2048 111134
rect -1964 110898 -1728 111134
rect -2284 75218 -2048 75454
rect -1964 75218 -1728 75454
rect -2284 74898 -2048 75134
rect -1964 74898 -1728 75134
rect -2284 39218 -2048 39454
rect -1964 39218 -1728 39454
rect -2284 38898 -2048 39134
rect -1964 38898 -1728 39134
rect -2284 3218 -2048 3454
rect -1964 3218 -1728 3454
rect -2284 2898 -2048 3134
rect -1964 2898 -1728 3134
rect -2284 -892 -2048 -656
rect -1964 -892 -1728 -656
rect -2284 -1212 -2048 -976
rect -1964 -1212 -1728 -976
rect 1826 704912 2062 705148
rect 2146 704912 2382 705148
rect 1826 704592 2062 704828
rect 2146 704592 2382 704828
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -892 2062 -656
rect 2146 -892 2382 -656
rect 1826 -1212 2062 -976
rect 2146 -1212 2382 -976
rect -3244 -1852 -3008 -1616
rect -2924 -1852 -2688 -1616
rect -3244 -2172 -3008 -1936
rect -2924 -2172 -2688 -1936
rect -4204 -2812 -3968 -2576
rect -3884 -2812 -3648 -2576
rect -4204 -3132 -3968 -2896
rect -3884 -3132 -3648 -2896
rect -5164 -3772 -4928 -3536
rect -4844 -3772 -4608 -3536
rect -5164 -4092 -4928 -3856
rect -4844 -4092 -4608 -3856
rect -6124 -4732 -5888 -4496
rect -5804 -4732 -5568 -4496
rect -6124 -5052 -5888 -4816
rect -5804 -5052 -5568 -4816
rect -7084 -5692 -6848 -5456
rect -6764 -5692 -6528 -5456
rect -7084 -6012 -6848 -5776
rect -6764 -6012 -6528 -5776
rect -8044 -6652 -7808 -6416
rect -7724 -6652 -7488 -6416
rect -8044 -6972 -7808 -6736
rect -7724 -6972 -7488 -6736
rect -9004 -7612 -8768 -7376
rect -8684 -7612 -8448 -7376
rect -9004 -7932 -8768 -7696
rect -8684 -7932 -8448 -7696
rect 6326 705872 6562 706108
rect 6646 705872 6882 706108
rect 6326 705552 6562 705788
rect 6646 705552 6882 705788
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1852 6562 -1616
rect 6646 -1852 6882 -1616
rect 6326 -2172 6562 -1936
rect 6646 -2172 6882 -1936
rect 10826 706832 11062 707068
rect 11146 706832 11382 707068
rect 10826 706512 11062 706748
rect 11146 706512 11382 706748
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2812 11062 -2576
rect 11146 -2812 11382 -2576
rect 10826 -3132 11062 -2896
rect 11146 -3132 11382 -2896
rect 15326 707792 15562 708028
rect 15646 707792 15882 708028
rect 15326 707472 15562 707708
rect 15646 707472 15882 707708
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3772 15562 -3536
rect 15646 -3772 15882 -3536
rect 15326 -4092 15562 -3856
rect 15646 -4092 15882 -3856
rect 19826 708752 20062 708988
rect 20146 708752 20382 708988
rect 19826 708432 20062 708668
rect 20146 708432 20382 708668
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4732 20062 -4496
rect 20146 -4732 20382 -4496
rect 19826 -5052 20062 -4816
rect 20146 -5052 20382 -4816
rect 24326 709712 24562 709948
rect 24646 709712 24882 709948
rect 24326 709392 24562 709628
rect 24646 709392 24882 709628
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5692 24562 -5456
rect 24646 -5692 24882 -5456
rect 24326 -6012 24562 -5776
rect 24646 -6012 24882 -5776
rect 28826 710672 29062 710908
rect 29146 710672 29382 710908
rect 28826 710352 29062 710588
rect 29146 710352 29382 710588
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6652 29062 -6416
rect 29146 -6652 29382 -6416
rect 28826 -6972 29062 -6736
rect 29146 -6972 29382 -6736
rect 33326 711632 33562 711868
rect 33646 711632 33882 711868
rect 33326 711312 33562 711548
rect 33646 711312 33882 711548
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7612 33562 -7376
rect 33646 -7612 33882 -7376
rect 33326 -7932 33562 -7696
rect 33646 -7932 33882 -7696
rect 37826 704912 38062 705148
rect 38146 704912 38382 705148
rect 37826 704592 38062 704828
rect 38146 704592 38382 704828
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -892 38062 -656
rect 38146 -892 38382 -656
rect 37826 -1212 38062 -976
rect 38146 -1212 38382 -976
rect 42326 705872 42562 706108
rect 42646 705872 42882 706108
rect 42326 705552 42562 705788
rect 42646 705552 42882 705788
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1852 42562 -1616
rect 42646 -1852 42882 -1616
rect 42326 -2172 42562 -1936
rect 42646 -2172 42882 -1936
rect 46826 706832 47062 707068
rect 47146 706832 47382 707068
rect 46826 706512 47062 706748
rect 47146 706512 47382 706748
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2812 47062 -2576
rect 47146 -2812 47382 -2576
rect 46826 -3132 47062 -2896
rect 47146 -3132 47382 -2896
rect 51326 707792 51562 708028
rect 51646 707792 51882 708028
rect 51326 707472 51562 707708
rect 51646 707472 51882 707708
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3772 51562 -3536
rect 51646 -3772 51882 -3536
rect 51326 -4092 51562 -3856
rect 51646 -4092 51882 -3856
rect 55826 708752 56062 708988
rect 56146 708752 56382 708988
rect 55826 708432 56062 708668
rect 56146 708432 56382 708668
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4732 56062 -4496
rect 56146 -4732 56382 -4496
rect 55826 -5052 56062 -4816
rect 56146 -5052 56382 -4816
rect 60326 709712 60562 709948
rect 60646 709712 60882 709948
rect 60326 709392 60562 709628
rect 60646 709392 60882 709628
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5692 60562 -5456
rect 60646 -5692 60882 -5456
rect 60326 -6012 60562 -5776
rect 60646 -6012 60882 -5776
rect 64826 710672 65062 710908
rect 65146 710672 65382 710908
rect 64826 710352 65062 710588
rect 65146 710352 65382 710588
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6652 65062 -6416
rect 65146 -6652 65382 -6416
rect 64826 -6972 65062 -6736
rect 65146 -6972 65382 -6736
rect 69326 711632 69562 711868
rect 69646 711632 69882 711868
rect 69326 711312 69562 711548
rect 69646 711312 69882 711548
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7612 69562 -7376
rect 69646 -7612 69882 -7376
rect 69326 -7932 69562 -7696
rect 69646 -7932 69882 -7696
rect 73826 704912 74062 705148
rect 74146 704912 74382 705148
rect 73826 704592 74062 704828
rect 74146 704592 74382 704828
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -892 74062 -656
rect 74146 -892 74382 -656
rect 73826 -1212 74062 -976
rect 74146 -1212 74382 -976
rect 78326 705872 78562 706108
rect 78646 705872 78882 706108
rect 78326 705552 78562 705788
rect 78646 705552 78882 705788
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1852 78562 -1616
rect 78646 -1852 78882 -1616
rect 78326 -2172 78562 -1936
rect 78646 -2172 78882 -1936
rect 82826 706832 83062 707068
rect 83146 706832 83382 707068
rect 82826 706512 83062 706748
rect 83146 706512 83382 706748
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2812 83062 -2576
rect 83146 -2812 83382 -2576
rect 82826 -3132 83062 -2896
rect 83146 -3132 83382 -2896
rect 87326 707792 87562 708028
rect 87646 707792 87882 708028
rect 87326 707472 87562 707708
rect 87646 707472 87882 707708
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3772 87562 -3536
rect 87646 -3772 87882 -3536
rect 87326 -4092 87562 -3856
rect 87646 -4092 87882 -3856
rect 91826 708752 92062 708988
rect 92146 708752 92382 708988
rect 91826 708432 92062 708668
rect 92146 708432 92382 708668
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4732 92062 -4496
rect 92146 -4732 92382 -4496
rect 91826 -5052 92062 -4816
rect 92146 -5052 92382 -4816
rect 96326 709712 96562 709948
rect 96646 709712 96882 709948
rect 96326 709392 96562 709628
rect 96646 709392 96882 709628
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 100826 710672 101062 710908
rect 101146 710672 101382 710908
rect 100826 710352 101062 710588
rect 101146 710352 101382 710588
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 105326 711632 105562 711868
rect 105646 711632 105882 711868
rect 105326 711312 105562 711548
rect 105646 711312 105882 711548
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 109826 704912 110062 705148
rect 110146 704912 110382 705148
rect 109826 704592 110062 704828
rect 110146 704592 110382 704828
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 114326 705872 114562 706108
rect 114646 705872 114882 706108
rect 114326 705552 114562 705788
rect 114646 705552 114882 705788
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 118826 706832 119062 707068
rect 119146 706832 119382 707068
rect 118826 706512 119062 706748
rect 119146 706512 119382 706748
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 123326 707792 123562 708028
rect 123646 707792 123882 708028
rect 123326 707472 123562 707708
rect 123646 707472 123882 707708
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 127826 708752 128062 708988
rect 128146 708752 128382 708988
rect 127826 708432 128062 708668
rect 128146 708432 128382 708668
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 132326 709712 132562 709948
rect 132646 709712 132882 709948
rect 132326 709392 132562 709628
rect 132646 709392 132882 709628
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 136826 710672 137062 710908
rect 137146 710672 137382 710908
rect 136826 710352 137062 710588
rect 137146 710352 137382 710588
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 141326 711632 141562 711868
rect 141646 711632 141882 711868
rect 141326 711312 141562 711548
rect 141646 711312 141882 711548
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 145826 704912 146062 705148
rect 146146 704912 146382 705148
rect 145826 704592 146062 704828
rect 146146 704592 146382 704828
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 150326 705872 150562 706108
rect 150646 705872 150882 706108
rect 150326 705552 150562 705788
rect 150646 705552 150882 705788
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 154826 706832 155062 707068
rect 155146 706832 155382 707068
rect 154826 706512 155062 706748
rect 155146 706512 155382 706748
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 159326 707792 159562 708028
rect 159646 707792 159882 708028
rect 159326 707472 159562 707708
rect 159646 707472 159882 707708
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 163826 708752 164062 708988
rect 164146 708752 164382 708988
rect 163826 708432 164062 708668
rect 164146 708432 164382 708668
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 168326 709712 168562 709948
rect 168646 709712 168882 709948
rect 168326 709392 168562 709628
rect 168646 709392 168882 709628
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 172826 710672 173062 710908
rect 173146 710672 173382 710908
rect 172826 710352 173062 710588
rect 173146 710352 173382 710588
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 119610 367718 119846 367954
rect 119610 367398 119846 367634
rect 150330 367718 150566 367954
rect 150330 367398 150566 367634
rect 104250 363218 104486 363454
rect 104250 362898 104486 363134
rect 134970 363218 135206 363454
rect 134970 362898 135206 363134
rect 165690 363218 165926 363454
rect 165690 362898 165926 363134
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 119610 331718 119846 331954
rect 119610 331398 119846 331634
rect 150330 331718 150566 331954
rect 150330 331398 150566 331634
rect 104250 327218 104486 327454
rect 104250 326898 104486 327134
rect 134970 327218 135206 327454
rect 134970 326898 135206 327134
rect 165690 327218 165926 327454
rect 165690 326898 165926 327134
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 96326 241718 96562 241954
rect 96646 241718 96882 241954
rect 96326 241398 96562 241634
rect 96646 241398 96882 241634
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5692 96562 -5456
rect 96646 -5692 96882 -5456
rect 96326 -6012 96562 -5776
rect 96646 -6012 96882 -5776
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 100826 246218 101062 246454
rect 101146 246218 101382 246454
rect 100826 245898 101062 246134
rect 101146 245898 101382 246134
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6652 101062 -6416
rect 101146 -6652 101382 -6416
rect 100826 -6972 101062 -6736
rect 101146 -6972 101382 -6736
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7612 105562 -7376
rect 105646 -7612 105882 -7376
rect 105326 -7932 105562 -7696
rect 105646 -7932 105882 -7696
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -892 110062 -656
rect 110146 -892 110382 -656
rect 109826 -1212 110062 -976
rect 110146 -1212 110382 -976
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1852 114562 -1616
rect 114646 -1852 114882 -1616
rect 114326 -2172 114562 -1936
rect 114646 -2172 114882 -1936
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 118826 228218 119062 228454
rect 119146 228218 119382 228454
rect 118826 227898 119062 228134
rect 119146 227898 119382 228134
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 118826 120218 119062 120454
rect 119146 120218 119382 120454
rect 118826 119898 119062 120134
rect 119146 119898 119382 120134
rect 118826 84218 119062 84454
rect 119146 84218 119382 84454
rect 118826 83898 119062 84134
rect 119146 83898 119382 84134
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2812 119062 -2576
rect 119146 -2812 119382 -2576
rect 118826 -3132 119062 -2896
rect 119146 -3132 119382 -2896
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 123326 232718 123562 232954
rect 123646 232718 123882 232954
rect 123326 232398 123562 232634
rect 123646 232398 123882 232634
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 123326 124718 123562 124954
rect 123646 124718 123882 124954
rect 123326 124398 123562 124634
rect 123646 124398 123882 124634
rect 123326 88718 123562 88954
rect 123646 88718 123882 88954
rect 123326 88398 123562 88634
rect 123646 88398 123882 88634
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3772 123562 -3536
rect 123646 -3772 123882 -3536
rect 123326 -4092 123562 -3856
rect 123646 -4092 123882 -3856
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4732 128062 -4496
rect 128146 -4732 128382 -4496
rect 127826 -5052 128062 -4816
rect 128146 -5052 128382 -4816
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 132326 241718 132562 241954
rect 132646 241718 132882 241954
rect 132326 241398 132562 241634
rect 132646 241398 132882 241634
rect 132326 205718 132562 205954
rect 132646 205718 132882 205954
rect 132326 205398 132562 205634
rect 132646 205398 132882 205634
rect 132326 169718 132562 169954
rect 132646 169718 132882 169954
rect 132326 169398 132562 169634
rect 132646 169398 132882 169634
rect 132326 133718 132562 133954
rect 132646 133718 132882 133954
rect 132326 133398 132562 133634
rect 132646 133398 132882 133634
rect 132326 97718 132562 97954
rect 132646 97718 132882 97954
rect 132326 97398 132562 97634
rect 132646 97398 132882 97634
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5692 132562 -5456
rect 132646 -5692 132882 -5456
rect 132326 -6012 132562 -5776
rect 132646 -6012 132882 -5776
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 136826 246218 137062 246454
rect 137146 246218 137382 246454
rect 136826 245898 137062 246134
rect 137146 245898 137382 246134
rect 136826 210218 137062 210454
rect 137146 210218 137382 210454
rect 136826 209898 137062 210134
rect 137146 209898 137382 210134
rect 136826 174218 137062 174454
rect 137146 174218 137382 174454
rect 136826 173898 137062 174134
rect 137146 173898 137382 174134
rect 136826 138218 137062 138454
rect 137146 138218 137382 138454
rect 136826 137898 137062 138134
rect 137146 137898 137382 138134
rect 136826 102218 137062 102454
rect 137146 102218 137382 102454
rect 136826 101898 137062 102134
rect 137146 101898 137382 102134
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6652 137062 -6416
rect 137146 -6652 137382 -6416
rect 136826 -6972 137062 -6736
rect 137146 -6972 137382 -6736
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 141326 214718 141562 214954
rect 141646 214718 141882 214954
rect 141326 214398 141562 214634
rect 141646 214398 141882 214634
rect 141326 178718 141562 178954
rect 141646 178718 141882 178954
rect 141326 178398 141562 178634
rect 141646 178398 141882 178634
rect 141326 142718 141562 142954
rect 141646 142718 141882 142954
rect 141326 142398 141562 142634
rect 141646 142398 141882 142634
rect 141326 106718 141562 106954
rect 141646 106718 141882 106954
rect 141326 106398 141562 106634
rect 141646 106398 141882 106634
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 141326 -7612 141562 -7376
rect 141646 -7612 141882 -7376
rect 141326 -7932 141562 -7696
rect 141646 -7932 141882 -7696
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -892 146062 -656
rect 146146 -892 146382 -656
rect 145826 -1212 146062 -976
rect 146146 -1212 146382 -976
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 150326 223718 150562 223954
rect 150646 223718 150882 223954
rect 150326 223398 150562 223634
rect 150646 223398 150882 223634
rect 150326 187718 150562 187954
rect 150646 187718 150882 187954
rect 150326 187398 150562 187634
rect 150646 187398 150882 187634
rect 150326 151718 150562 151954
rect 150646 151718 150882 151954
rect 150326 151398 150562 151634
rect 150646 151398 150882 151634
rect 150326 115718 150562 115954
rect 150646 115718 150882 115954
rect 150326 115398 150562 115634
rect 150646 115398 150882 115634
rect 150326 79718 150562 79954
rect 150646 79718 150882 79954
rect 150326 79398 150562 79634
rect 150646 79398 150882 79634
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1852 150562 -1616
rect 150646 -1852 150882 -1616
rect 150326 -2172 150562 -1936
rect 150646 -2172 150882 -1936
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 154826 228218 155062 228454
rect 155146 228218 155382 228454
rect 154826 227898 155062 228134
rect 155146 227898 155382 228134
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 154826 156218 155062 156454
rect 155146 156218 155382 156454
rect 154826 155898 155062 156134
rect 155146 155898 155382 156134
rect 154826 120218 155062 120454
rect 155146 120218 155382 120454
rect 154826 119898 155062 120134
rect 155146 119898 155382 120134
rect 154826 84218 155062 84454
rect 155146 84218 155382 84454
rect 154826 83898 155062 84134
rect 155146 83898 155382 84134
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2812 155062 -2576
rect 155146 -2812 155382 -2576
rect 154826 -3132 155062 -2896
rect 155146 -3132 155382 -2896
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 159326 232718 159562 232954
rect 159646 232718 159882 232954
rect 159326 232398 159562 232634
rect 159646 232398 159882 232634
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 159326 160718 159562 160954
rect 159646 160718 159882 160954
rect 159326 160398 159562 160634
rect 159646 160398 159882 160634
rect 159326 124718 159562 124954
rect 159646 124718 159882 124954
rect 159326 124398 159562 124634
rect 159646 124398 159882 124634
rect 159326 88718 159562 88954
rect 159646 88718 159882 88954
rect 159326 88398 159562 88634
rect 159646 88398 159882 88634
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3772 159562 -3536
rect 159646 -3772 159882 -3536
rect 159326 -4092 159562 -3856
rect 159646 -4092 159882 -3856
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4732 164062 -4496
rect 164146 -4732 164382 -4496
rect 163826 -5052 164062 -4816
rect 164146 -5052 164382 -4816
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 168326 241718 168562 241954
rect 168646 241718 168882 241954
rect 168326 241398 168562 241634
rect 168646 241398 168882 241634
rect 168326 205718 168562 205954
rect 168646 205718 168882 205954
rect 168326 205398 168562 205634
rect 168646 205398 168882 205634
rect 168326 169718 168562 169954
rect 168646 169718 168882 169954
rect 168326 169398 168562 169634
rect 168646 169398 168882 169634
rect 168326 133718 168562 133954
rect 168646 133718 168882 133954
rect 168326 133398 168562 133634
rect 168646 133398 168882 133634
rect 168326 97718 168562 97954
rect 168646 97718 168882 97954
rect 168326 97398 168562 97634
rect 168646 97398 168882 97634
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5692 168562 -5456
rect 168646 -5692 168882 -5456
rect 168326 -6012 168562 -5776
rect 168646 -6012 168882 -5776
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 172826 246218 173062 246454
rect 173146 246218 173382 246454
rect 172826 245898 173062 246134
rect 173146 245898 173382 246134
rect 172826 210218 173062 210454
rect 173146 210218 173382 210454
rect 172826 209898 173062 210134
rect 173146 209898 173382 210134
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 172826 138218 173062 138454
rect 173146 138218 173382 138454
rect 172826 137898 173062 138134
rect 173146 137898 173382 138134
rect 172826 102218 173062 102454
rect 173146 102218 173382 102454
rect 172826 101898 173062 102134
rect 173146 101898 173382 102134
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6652 173062 -6416
rect 173146 -6652 173382 -6416
rect 172826 -6972 173062 -6736
rect 173146 -6972 173382 -6736
rect 177326 711632 177562 711868
rect 177646 711632 177882 711868
rect 177326 711312 177562 711548
rect 177646 711312 177882 711548
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 177326 214718 177562 214954
rect 177646 214718 177882 214954
rect 177326 214398 177562 214634
rect 177646 214398 177882 214634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 177326 106718 177562 106954
rect 177646 106718 177882 106954
rect 177326 106398 177562 106634
rect 177646 106398 177882 106634
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7612 177562 -7376
rect 177646 -7612 177882 -7376
rect 177326 -7932 177562 -7696
rect 177646 -7932 177882 -7696
rect 181826 704912 182062 705148
rect 182146 704912 182382 705148
rect 181826 704592 182062 704828
rect 182146 704592 182382 704828
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -892 182062 -656
rect 182146 -892 182382 -656
rect 181826 -1212 182062 -976
rect 182146 -1212 182382 -976
rect 186326 705872 186562 706108
rect 186646 705872 186882 706108
rect 186326 705552 186562 705788
rect 186646 705552 186882 705788
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1852 186562 -1616
rect 186646 -1852 186882 -1616
rect 186326 -2172 186562 -1936
rect 186646 -2172 186882 -1936
rect 190826 706832 191062 707068
rect 191146 706832 191382 707068
rect 190826 706512 191062 706748
rect 191146 706512 191382 706748
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 190826 228218 191062 228454
rect 191146 228218 191382 228454
rect 190826 227898 191062 228134
rect 191146 227898 191382 228134
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2812 191062 -2576
rect 191146 -2812 191382 -2576
rect 190826 -3132 191062 -2896
rect 191146 -3132 191382 -2896
rect 195326 707792 195562 708028
rect 195646 707792 195882 708028
rect 195326 707472 195562 707708
rect 195646 707472 195882 707708
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3772 195562 -3536
rect 195646 -3772 195882 -3536
rect 195326 -4092 195562 -3856
rect 195646 -4092 195882 -3856
rect 199826 708752 200062 708988
rect 200146 708752 200382 708988
rect 199826 708432 200062 708668
rect 200146 708432 200382 708668
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4732 200062 -4496
rect 200146 -4732 200382 -4496
rect 199826 -5052 200062 -4816
rect 200146 -5052 200382 -4816
rect 204326 709712 204562 709948
rect 204646 709712 204882 709948
rect 204326 709392 204562 709628
rect 204646 709392 204882 709628
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 204326 241718 204562 241954
rect 204646 241718 204882 241954
rect 204326 241398 204562 241634
rect 204646 241398 204882 241634
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5692 204562 -5456
rect 204646 -5692 204882 -5456
rect 204326 -6012 204562 -5776
rect 204646 -6012 204882 -5776
rect 208826 710672 209062 710908
rect 209146 710672 209382 710908
rect 208826 710352 209062 710588
rect 209146 710352 209382 710588
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 208826 246218 209062 246454
rect 209146 246218 209382 246454
rect 208826 245898 209062 246134
rect 209146 245898 209382 246134
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6652 209062 -6416
rect 209146 -6652 209382 -6416
rect 208826 -6972 209062 -6736
rect 209146 -6972 209382 -6736
rect 213326 711632 213562 711868
rect 213646 711632 213882 711868
rect 213326 711312 213562 711548
rect 213646 711312 213882 711548
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 217826 704912 218062 705148
rect 218146 704912 218382 705148
rect 217826 704592 218062 704828
rect 218146 704592 218382 704828
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 222326 705872 222562 706108
rect 222646 705872 222882 706108
rect 222326 705552 222562 705788
rect 222646 705552 222882 705788
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 226826 706832 227062 707068
rect 227146 706832 227382 707068
rect 226826 706512 227062 706748
rect 227146 706512 227382 706748
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 231326 707792 231562 708028
rect 231646 707792 231882 708028
rect 231326 707472 231562 707708
rect 231646 707472 231882 707708
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 235826 708752 236062 708988
rect 236146 708752 236382 708988
rect 235826 708432 236062 708668
rect 236146 708432 236382 708668
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 240326 709712 240562 709948
rect 240646 709712 240882 709948
rect 240326 709392 240562 709628
rect 240646 709392 240882 709628
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 244826 710672 245062 710908
rect 245146 710672 245382 710908
rect 244826 710352 245062 710588
rect 245146 710352 245382 710588
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 249326 711632 249562 711868
rect 249646 711632 249882 711868
rect 249326 711312 249562 711548
rect 249646 711312 249882 711548
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 253826 704912 254062 705148
rect 254146 704912 254382 705148
rect 253826 704592 254062 704828
rect 254146 704592 254382 704828
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 258326 705872 258562 706108
rect 258646 705872 258882 706108
rect 258326 705552 258562 705788
rect 258646 705552 258882 705788
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 262826 706832 263062 707068
rect 263146 706832 263382 707068
rect 262826 706512 263062 706748
rect 263146 706512 263382 706748
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 267326 707792 267562 708028
rect 267646 707792 267882 708028
rect 267326 707472 267562 707708
rect 267646 707472 267882 707708
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 271826 708752 272062 708988
rect 272146 708752 272382 708988
rect 271826 708432 272062 708668
rect 272146 708432 272382 708668
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 276326 709712 276562 709948
rect 276646 709712 276882 709948
rect 276326 709392 276562 709628
rect 276646 709392 276882 709628
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 280826 710672 281062 710908
rect 281146 710672 281382 710908
rect 280826 710352 281062 710588
rect 281146 710352 281382 710588
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 285326 711632 285562 711868
rect 285646 711632 285882 711868
rect 285326 711312 285562 711548
rect 285646 711312 285882 711548
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 289826 704912 290062 705148
rect 290146 704912 290382 705148
rect 289826 704592 290062 704828
rect 290146 704592 290382 704828
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 294326 705872 294562 706108
rect 294646 705872 294882 706108
rect 294326 705552 294562 705788
rect 294646 705552 294882 705788
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 298826 706832 299062 707068
rect 299146 706832 299382 707068
rect 298826 706512 299062 706748
rect 299146 706512 299382 706748
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 303326 707792 303562 708028
rect 303646 707792 303882 708028
rect 303326 707472 303562 707708
rect 303646 707472 303882 707708
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 307826 708752 308062 708988
rect 308146 708752 308382 708988
rect 307826 708432 308062 708668
rect 308146 708432 308382 708668
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 312326 709712 312562 709948
rect 312646 709712 312882 709948
rect 312326 709392 312562 709628
rect 312646 709392 312882 709628
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 316826 710672 317062 710908
rect 317146 710672 317382 710908
rect 316826 710352 317062 710588
rect 317146 710352 317382 710588
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 321326 711632 321562 711868
rect 321646 711632 321882 711868
rect 321326 711312 321562 711548
rect 321646 711312 321882 711548
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 325826 704912 326062 705148
rect 326146 704912 326382 705148
rect 325826 704592 326062 704828
rect 326146 704592 326382 704828
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 330326 705872 330562 706108
rect 330646 705872 330882 706108
rect 330326 705552 330562 705788
rect 330646 705552 330882 705788
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 334826 706832 335062 707068
rect 335146 706832 335382 707068
rect 334826 706512 335062 706748
rect 335146 706512 335382 706748
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 339326 707792 339562 708028
rect 339646 707792 339882 708028
rect 339326 707472 339562 707708
rect 339646 707472 339882 707708
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 343826 708752 344062 708988
rect 344146 708752 344382 708988
rect 343826 708432 344062 708668
rect 344146 708432 344382 708668
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 348326 709712 348562 709948
rect 348646 709712 348882 709948
rect 348326 709392 348562 709628
rect 348646 709392 348882 709628
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 352826 710672 353062 710908
rect 353146 710672 353382 710908
rect 352826 710352 353062 710588
rect 353146 710352 353382 710588
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 357326 711632 357562 711868
rect 357646 711632 357882 711868
rect 357326 711312 357562 711548
rect 357646 711312 357882 711548
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 361826 704912 362062 705148
rect 362146 704912 362382 705148
rect 361826 704592 362062 704828
rect 362146 704592 362382 704828
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 220328 547718 220564 547954
rect 220328 547398 220564 547634
rect 356056 547718 356292 547954
rect 356056 547398 356292 547634
rect 221008 543218 221244 543454
rect 221008 542898 221244 543134
rect 355376 543218 355612 543454
rect 355376 542898 355612 543134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 220328 511718 220564 511954
rect 220328 511398 220564 511634
rect 356056 511718 356292 511954
rect 356056 511398 356292 511634
rect 221008 507218 221244 507454
rect 221008 506898 221244 507134
rect 355376 507218 355612 507454
rect 355376 506898 355612 507134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 366326 705872 366562 706108
rect 366646 705872 366882 706108
rect 366326 705552 366562 705788
rect 366646 705552 366882 705788
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 236650 435218 236886 435454
rect 236650 434898 236886 435134
rect 267370 435218 267606 435454
rect 267370 434898 267606 435134
rect 298090 435218 298326 435454
rect 298090 434898 298326 435134
rect 328810 435218 329046 435454
rect 328810 434898 329046 435134
rect 359530 435218 359766 435454
rect 359530 434898 359766 435134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 252010 403718 252246 403954
rect 252010 403398 252246 403634
rect 282730 403718 282966 403954
rect 282730 403398 282966 403634
rect 313450 403718 313686 403954
rect 313450 403398 313686 403634
rect 344170 403718 344406 403954
rect 344170 403398 344406 403634
rect 236650 399218 236886 399454
rect 236650 398898 236886 399134
rect 267370 399218 267606 399454
rect 267370 398898 267606 399134
rect 298090 399218 298326 399454
rect 298090 398898 298326 399134
rect 328810 399218 329046 399454
rect 328810 398898 329046 399134
rect 359530 399218 359766 399454
rect 359530 398898 359766 399134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 252010 367718 252246 367954
rect 252010 367398 252246 367634
rect 282730 367718 282966 367954
rect 282730 367398 282966 367634
rect 313450 367718 313686 367954
rect 313450 367398 313686 367634
rect 344170 367718 344406 367954
rect 344170 367398 344406 367634
rect 236650 363218 236886 363454
rect 236650 362898 236886 363134
rect 267370 363218 267606 363454
rect 267370 362898 267606 363134
rect 298090 363218 298326 363454
rect 298090 362898 298326 363134
rect 328810 363218 329046 363454
rect 328810 362898 329046 363134
rect 359530 363218 359766 363454
rect 359530 362898 359766 363134
rect 252010 331718 252246 331954
rect 252010 331398 252246 331634
rect 282730 331718 282966 331954
rect 282730 331398 282966 331634
rect 313450 331718 313686 331954
rect 313450 331398 313686 331634
rect 344170 331718 344406 331954
rect 344170 331398 344406 331634
rect 236650 327218 236886 327454
rect 236650 326898 236886 327134
rect 267370 327218 267606 327454
rect 267370 326898 267606 327134
rect 298090 327218 298326 327454
rect 298090 326898 298326 327134
rect 328810 327218 329046 327454
rect 328810 326898 329046 327134
rect 359530 327218 359766 327454
rect 359530 326898 359766 327134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 244826 246218 245062 246454
rect 245146 246218 245382 246454
rect 244826 245898 245062 246134
rect 245146 245898 245382 246134
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 280826 246218 281062 246454
rect 281146 246218 281382 246454
rect 280826 245898 281062 246134
rect 281146 245898 281382 246134
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 316826 246218 317062 246454
rect 317146 246218 317382 246454
rect 316826 245898 317062 246134
rect 317146 245898 317382 246134
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 220328 223718 220564 223954
rect 220328 223398 220564 223634
rect 356056 223718 356292 223954
rect 356056 223398 356292 223634
rect 221008 219218 221244 219454
rect 221008 218898 221244 219134
rect 355376 219218 355612 219454
rect 355376 218898 355612 219134
rect 220328 187718 220564 187954
rect 220328 187398 220564 187634
rect 356056 187718 356292 187954
rect 356056 187398 356292 187634
rect 221008 183218 221244 183454
rect 221008 182898 221244 183134
rect 355376 183218 355612 183454
rect 355376 182898 355612 183134
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 213326 -7612 213562 -7376
rect 213646 -7612 213882 -7376
rect 213326 -7932 213562 -7696
rect 213646 -7932 213882 -7696
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -892 218062 -656
rect 218146 -892 218382 -656
rect 217826 -1212 218062 -976
rect 218146 -1212 218382 -976
rect 222326 -1852 222562 -1616
rect 222646 -1852 222882 -1616
rect 222326 -2172 222562 -1936
rect 222646 -2172 222882 -1936
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2812 227062 -2576
rect 227146 -2812 227382 -2576
rect 226826 -3132 227062 -2896
rect 227146 -3132 227382 -2896
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3772 231562 -3536
rect 231646 -3772 231882 -3536
rect 231326 -4092 231562 -3856
rect 231646 -4092 231882 -3856
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4732 236062 -4496
rect 236146 -4732 236382 -4496
rect 235826 -5052 236062 -4816
rect 236146 -5052 236382 -4816
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5692 240562 -5456
rect 240646 -5692 240882 -5456
rect 240326 -6012 240562 -5776
rect 240646 -6012 240882 -5776
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6652 245062 -6416
rect 245146 -6652 245382 -6416
rect 244826 -6972 245062 -6736
rect 245146 -6972 245382 -6736
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7612 249562 -7376
rect 249646 -7612 249882 -7376
rect 249326 -7932 249562 -7696
rect 249646 -7932 249882 -7696
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -892 254062 -656
rect 254146 -892 254382 -656
rect 253826 -1212 254062 -976
rect 254146 -1212 254382 -976
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1852 258562 -1616
rect 258646 -1852 258882 -1616
rect 258326 -2172 258562 -1936
rect 258646 -2172 258882 -1936
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2812 263062 -2576
rect 263146 -2812 263382 -2576
rect 262826 -3132 263062 -2896
rect 263146 -3132 263382 -2896
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3772 267562 -3536
rect 267646 -3772 267882 -3536
rect 267326 -4092 267562 -3856
rect 267646 -4092 267882 -3856
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4732 272062 -4496
rect 272146 -4732 272382 -4496
rect 271826 -5052 272062 -4816
rect 272146 -5052 272382 -4816
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5692 276562 -5456
rect 276646 -5692 276882 -5456
rect 276326 -6012 276562 -5776
rect 276646 -6012 276882 -5776
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6652 281062 -6416
rect 281146 -6652 281382 -6416
rect 280826 -6972 281062 -6736
rect 281146 -6972 281382 -6736
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7612 285562 -7376
rect 285646 -7612 285882 -7376
rect 285326 -7932 285562 -7696
rect 285646 -7932 285882 -7696
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -892 290062 -656
rect 290146 -892 290382 -656
rect 289826 -1212 290062 -976
rect 290146 -1212 290382 -976
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1852 294562 -1616
rect 294646 -1852 294882 -1616
rect 294326 -2172 294562 -1936
rect 294646 -2172 294882 -1936
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2812 299062 -2576
rect 299146 -2812 299382 -2576
rect 298826 -3132 299062 -2896
rect 299146 -3132 299382 -2896
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3772 303562 -3536
rect 303646 -3772 303882 -3536
rect 303326 -4092 303562 -3856
rect 303646 -4092 303882 -3856
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4732 308062 -4496
rect 308146 -4732 308382 -4496
rect 307826 -5052 308062 -4816
rect 308146 -5052 308382 -4816
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5692 312562 -5456
rect 312646 -5692 312882 -5456
rect 312326 -6012 312562 -5776
rect 312646 -6012 312882 -5776
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6652 317062 -6416
rect 317146 -6652 317382 -6416
rect 316826 -6972 317062 -6736
rect 317146 -6972 317382 -6736
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7612 321562 -7376
rect 321646 -7612 321882 -7376
rect 321326 -7932 321562 -7696
rect 321646 -7932 321882 -7696
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -892 326062 -656
rect 326146 -892 326382 -656
rect 325826 -1212 326062 -976
rect 326146 -1212 326382 -976
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1852 330562 -1616
rect 330646 -1852 330882 -1616
rect 330326 -2172 330562 -1936
rect 330646 -2172 330882 -1936
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2812 335062 -2576
rect 335146 -2812 335382 -2576
rect 334826 -3132 335062 -2896
rect 335146 -3132 335382 -2896
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3772 339562 -3536
rect 339646 -3772 339882 -3536
rect 339326 -4092 339562 -3856
rect 339646 -4092 339882 -3856
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4732 344062 -4496
rect 344146 -4732 344382 -4496
rect 343826 -5052 344062 -4816
rect 344146 -5052 344382 -4816
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5692 348562 -5456
rect 348646 -5692 348882 -5456
rect 348326 -6012 348562 -5776
rect 348646 -6012 348882 -5776
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6652 353062 -6416
rect 353146 -6652 353382 -6416
rect 352826 -6972 353062 -6736
rect 353146 -6972 353382 -6736
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 357326 -7612 357562 -7376
rect 357646 -7612 357882 -7376
rect 357326 -7932 357562 -7696
rect 357646 -7932 357882 -7696
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 370826 706832 371062 707068
rect 371146 706832 371382 707068
rect 370826 706512 371062 706748
rect 371146 706512 371382 706748
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 361826 -892 362062 -656
rect 362146 -892 362382 -656
rect 361826 -1212 362062 -976
rect 362146 -1212 362382 -976
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 366326 -1852 366562 -1616
rect 366646 -1852 366882 -1616
rect 366326 -2172 366562 -1936
rect 366646 -2172 366882 -1936
rect 370826 -2812 371062 -2576
rect 371146 -2812 371382 -2576
rect 370826 -3132 371062 -2896
rect 371146 -3132 371382 -2896
rect 375326 707792 375562 708028
rect 375646 707792 375882 708028
rect 375326 707472 375562 707708
rect 375646 707472 375882 707708
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3772 375562 -3536
rect 375646 -3772 375882 -3536
rect 375326 -4092 375562 -3856
rect 375646 -4092 375882 -3856
rect 379826 708752 380062 708988
rect 380146 708752 380382 708988
rect 379826 708432 380062 708668
rect 380146 708432 380382 708668
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4732 380062 -4496
rect 380146 -4732 380382 -4496
rect 379826 -5052 380062 -4816
rect 380146 -5052 380382 -4816
rect 384326 709712 384562 709948
rect 384646 709712 384882 709948
rect 384326 709392 384562 709628
rect 384646 709392 384882 709628
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5692 384562 -5456
rect 384646 -5692 384882 -5456
rect 384326 -6012 384562 -5776
rect 384646 -6012 384882 -5776
rect 388826 710672 389062 710908
rect 389146 710672 389382 710908
rect 388826 710352 389062 710588
rect 389146 710352 389382 710588
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6652 389062 -6416
rect 389146 -6652 389382 -6416
rect 388826 -6972 389062 -6736
rect 389146 -6972 389382 -6736
rect 393326 711632 393562 711868
rect 393646 711632 393882 711868
rect 393326 711312 393562 711548
rect 393646 711312 393882 711548
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7612 393562 -7376
rect 393646 -7612 393882 -7376
rect 393326 -7932 393562 -7696
rect 393646 -7932 393882 -7696
rect 397826 704912 398062 705148
rect 398146 704912 398382 705148
rect 397826 704592 398062 704828
rect 398146 704592 398382 704828
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -892 398062 -656
rect 398146 -892 398382 -656
rect 397826 -1212 398062 -976
rect 398146 -1212 398382 -976
rect 402326 705872 402562 706108
rect 402646 705872 402882 706108
rect 402326 705552 402562 705788
rect 402646 705552 402882 705788
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1852 402562 -1616
rect 402646 -1852 402882 -1616
rect 402326 -2172 402562 -1936
rect 402646 -2172 402882 -1936
rect 406826 706832 407062 707068
rect 407146 706832 407382 707068
rect 406826 706512 407062 706748
rect 407146 706512 407382 706748
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2812 407062 -2576
rect 407146 -2812 407382 -2576
rect 406826 -3132 407062 -2896
rect 407146 -3132 407382 -2896
rect 411326 707792 411562 708028
rect 411646 707792 411882 708028
rect 411326 707472 411562 707708
rect 411646 707472 411882 707708
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3772 411562 -3536
rect 411646 -3772 411882 -3536
rect 411326 -4092 411562 -3856
rect 411646 -4092 411882 -3856
rect 415826 708752 416062 708988
rect 416146 708752 416382 708988
rect 415826 708432 416062 708668
rect 416146 708432 416382 708668
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4732 416062 -4496
rect 416146 -4732 416382 -4496
rect 415826 -5052 416062 -4816
rect 416146 -5052 416382 -4816
rect 420326 709712 420562 709948
rect 420646 709712 420882 709948
rect 420326 709392 420562 709628
rect 420646 709392 420882 709628
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5692 420562 -5456
rect 420646 -5692 420882 -5456
rect 420326 -6012 420562 -5776
rect 420646 -6012 420882 -5776
rect 424826 710672 425062 710908
rect 425146 710672 425382 710908
rect 424826 710352 425062 710588
rect 425146 710352 425382 710588
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6652 425062 -6416
rect 425146 -6652 425382 -6416
rect 424826 -6972 425062 -6736
rect 425146 -6972 425382 -6736
rect 429326 711632 429562 711868
rect 429646 711632 429882 711868
rect 429326 711312 429562 711548
rect 429646 711312 429882 711548
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7612 429562 -7376
rect 429646 -7612 429882 -7376
rect 429326 -7932 429562 -7696
rect 429646 -7932 429882 -7696
rect 433826 704912 434062 705148
rect 434146 704912 434382 705148
rect 433826 704592 434062 704828
rect 434146 704592 434382 704828
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -892 434062 -656
rect 434146 -892 434382 -656
rect 433826 -1212 434062 -976
rect 434146 -1212 434382 -976
rect 438326 705872 438562 706108
rect 438646 705872 438882 706108
rect 438326 705552 438562 705788
rect 438646 705552 438882 705788
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1852 438562 -1616
rect 438646 -1852 438882 -1616
rect 438326 -2172 438562 -1936
rect 438646 -2172 438882 -1936
rect 442826 706832 443062 707068
rect 443146 706832 443382 707068
rect 442826 706512 443062 706748
rect 443146 706512 443382 706748
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2812 443062 -2576
rect 443146 -2812 443382 -2576
rect 442826 -3132 443062 -2896
rect 443146 -3132 443382 -2896
rect 447326 707792 447562 708028
rect 447646 707792 447882 708028
rect 447326 707472 447562 707708
rect 447646 707472 447882 707708
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3772 447562 -3536
rect 447646 -3772 447882 -3536
rect 447326 -4092 447562 -3856
rect 447646 -4092 447882 -3856
rect 451826 708752 452062 708988
rect 452146 708752 452382 708988
rect 451826 708432 452062 708668
rect 452146 708432 452382 708668
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4732 452062 -4496
rect 452146 -4732 452382 -4496
rect 451826 -5052 452062 -4816
rect 452146 -5052 452382 -4816
rect 456326 709712 456562 709948
rect 456646 709712 456882 709948
rect 456326 709392 456562 709628
rect 456646 709392 456882 709628
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5692 456562 -5456
rect 456646 -5692 456882 -5456
rect 456326 -6012 456562 -5776
rect 456646 -6012 456882 -5776
rect 460826 710672 461062 710908
rect 461146 710672 461382 710908
rect 460826 710352 461062 710588
rect 461146 710352 461382 710588
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6652 461062 -6416
rect 461146 -6652 461382 -6416
rect 460826 -6972 461062 -6736
rect 461146 -6972 461382 -6736
rect 465326 711632 465562 711868
rect 465646 711632 465882 711868
rect 465326 711312 465562 711548
rect 465646 711312 465882 711548
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7612 465562 -7376
rect 465646 -7612 465882 -7376
rect 465326 -7932 465562 -7696
rect 465646 -7932 465882 -7696
rect 469826 704912 470062 705148
rect 470146 704912 470382 705148
rect 469826 704592 470062 704828
rect 470146 704592 470382 704828
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -892 470062 -656
rect 470146 -892 470382 -656
rect 469826 -1212 470062 -976
rect 470146 -1212 470382 -976
rect 474326 705872 474562 706108
rect 474646 705872 474882 706108
rect 474326 705552 474562 705788
rect 474646 705552 474882 705788
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1852 474562 -1616
rect 474646 -1852 474882 -1616
rect 474326 -2172 474562 -1936
rect 474646 -2172 474882 -1936
rect 478826 706832 479062 707068
rect 479146 706832 479382 707068
rect 478826 706512 479062 706748
rect 479146 706512 479382 706748
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2812 479062 -2576
rect 479146 -2812 479382 -2576
rect 478826 -3132 479062 -2896
rect 479146 -3132 479382 -2896
rect 483326 707792 483562 708028
rect 483646 707792 483882 708028
rect 483326 707472 483562 707708
rect 483646 707472 483882 707708
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3772 483562 -3536
rect 483646 -3772 483882 -3536
rect 483326 -4092 483562 -3856
rect 483646 -4092 483882 -3856
rect 487826 708752 488062 708988
rect 488146 708752 488382 708988
rect 487826 708432 488062 708668
rect 488146 708432 488382 708668
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4732 488062 -4496
rect 488146 -4732 488382 -4496
rect 487826 -5052 488062 -4816
rect 488146 -5052 488382 -4816
rect 492326 709712 492562 709948
rect 492646 709712 492882 709948
rect 492326 709392 492562 709628
rect 492646 709392 492882 709628
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5692 492562 -5456
rect 492646 -5692 492882 -5456
rect 492326 -6012 492562 -5776
rect 492646 -6012 492882 -5776
rect 496826 710672 497062 710908
rect 497146 710672 497382 710908
rect 496826 710352 497062 710588
rect 497146 710352 497382 710588
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6652 497062 -6416
rect 497146 -6652 497382 -6416
rect 496826 -6972 497062 -6736
rect 497146 -6972 497382 -6736
rect 501326 711632 501562 711868
rect 501646 711632 501882 711868
rect 501326 711312 501562 711548
rect 501646 711312 501882 711548
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7612 501562 -7376
rect 501646 -7612 501882 -7376
rect 501326 -7932 501562 -7696
rect 501646 -7932 501882 -7696
rect 505826 704912 506062 705148
rect 506146 704912 506382 705148
rect 505826 704592 506062 704828
rect 506146 704592 506382 704828
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -892 506062 -656
rect 506146 -892 506382 -656
rect 505826 -1212 506062 -976
rect 506146 -1212 506382 -976
rect 510326 705872 510562 706108
rect 510646 705872 510882 706108
rect 510326 705552 510562 705788
rect 510646 705552 510882 705788
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1852 510562 -1616
rect 510646 -1852 510882 -1616
rect 510326 -2172 510562 -1936
rect 510646 -2172 510882 -1936
rect 514826 706832 515062 707068
rect 515146 706832 515382 707068
rect 514826 706512 515062 706748
rect 515146 706512 515382 706748
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2812 515062 -2576
rect 515146 -2812 515382 -2576
rect 514826 -3132 515062 -2896
rect 515146 -3132 515382 -2896
rect 519326 707792 519562 708028
rect 519646 707792 519882 708028
rect 519326 707472 519562 707708
rect 519646 707472 519882 707708
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3772 519562 -3536
rect 519646 -3772 519882 -3536
rect 519326 -4092 519562 -3856
rect 519646 -4092 519882 -3856
rect 523826 708752 524062 708988
rect 524146 708752 524382 708988
rect 523826 708432 524062 708668
rect 524146 708432 524382 708668
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4732 524062 -4496
rect 524146 -4732 524382 -4496
rect 523826 -5052 524062 -4816
rect 524146 -5052 524382 -4816
rect 528326 709712 528562 709948
rect 528646 709712 528882 709948
rect 528326 709392 528562 709628
rect 528646 709392 528882 709628
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5692 528562 -5456
rect 528646 -5692 528882 -5456
rect 528326 -6012 528562 -5776
rect 528646 -6012 528882 -5776
rect 532826 710672 533062 710908
rect 533146 710672 533382 710908
rect 532826 710352 533062 710588
rect 533146 710352 533382 710588
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6652 533062 -6416
rect 533146 -6652 533382 -6416
rect 532826 -6972 533062 -6736
rect 533146 -6972 533382 -6736
rect 537326 711632 537562 711868
rect 537646 711632 537882 711868
rect 537326 711312 537562 711548
rect 537646 711312 537882 711548
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7612 537562 -7376
rect 537646 -7612 537882 -7376
rect 537326 -7932 537562 -7696
rect 537646 -7932 537882 -7696
rect 541826 704912 542062 705148
rect 542146 704912 542382 705148
rect 541826 704592 542062 704828
rect 542146 704592 542382 704828
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -892 542062 -656
rect 542146 -892 542382 -656
rect 541826 -1212 542062 -976
rect 542146 -1212 542382 -976
rect 546326 705872 546562 706108
rect 546646 705872 546882 706108
rect 546326 705552 546562 705788
rect 546646 705552 546882 705788
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1852 546562 -1616
rect 546646 -1852 546882 -1616
rect 546326 -2172 546562 -1936
rect 546646 -2172 546882 -1936
rect 550826 706832 551062 707068
rect 551146 706832 551382 707068
rect 550826 706512 551062 706748
rect 551146 706512 551382 706748
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2812 551062 -2576
rect 551146 -2812 551382 -2576
rect 550826 -3132 551062 -2896
rect 551146 -3132 551382 -2896
rect 555326 707792 555562 708028
rect 555646 707792 555882 708028
rect 555326 707472 555562 707708
rect 555646 707472 555882 707708
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3772 555562 -3536
rect 555646 -3772 555882 -3536
rect 555326 -4092 555562 -3856
rect 555646 -4092 555882 -3856
rect 559826 708752 560062 708988
rect 560146 708752 560382 708988
rect 559826 708432 560062 708668
rect 560146 708432 560382 708668
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4732 560062 -4496
rect 560146 -4732 560382 -4496
rect 559826 -5052 560062 -4816
rect 560146 -5052 560382 -4816
rect 564326 709712 564562 709948
rect 564646 709712 564882 709948
rect 564326 709392 564562 709628
rect 564646 709392 564882 709628
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5692 564562 -5456
rect 564646 -5692 564882 -5456
rect 564326 -6012 564562 -5776
rect 564646 -6012 564882 -5776
rect 568826 710672 569062 710908
rect 569146 710672 569382 710908
rect 568826 710352 569062 710588
rect 569146 710352 569382 710588
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6652 569062 -6416
rect 569146 -6652 569382 -6416
rect 568826 -6972 569062 -6736
rect 569146 -6972 569382 -6736
rect 573326 711632 573562 711868
rect 573646 711632 573882 711868
rect 573326 711312 573562 711548
rect 573646 711312 573882 711548
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7612 573562 -7376
rect 573646 -7612 573882 -7376
rect 573326 -7932 573562 -7696
rect 573646 -7932 573882 -7696
rect 577826 704912 578062 705148
rect 578146 704912 578382 705148
rect 577826 704592 578062 704828
rect 578146 704592 578382 704828
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -892 578062 -656
rect 578146 -892 578382 -656
rect 577826 -1212 578062 -976
rect 578146 -1212 578382 -976
rect 592372 711632 592608 711868
rect 592692 711632 592928 711868
rect 592372 711312 592608 711548
rect 592692 711312 592928 711548
rect 591412 710672 591648 710908
rect 591732 710672 591968 710908
rect 591412 710352 591648 710588
rect 591732 710352 591968 710588
rect 590452 709712 590688 709948
rect 590772 709712 591008 709948
rect 590452 709392 590688 709628
rect 590772 709392 591008 709628
rect 589492 708752 589728 708988
rect 589812 708752 590048 708988
rect 589492 708432 589728 708668
rect 589812 708432 590048 708668
rect 588532 707792 588768 708028
rect 588852 707792 589088 708028
rect 588532 707472 588768 707708
rect 588852 707472 589088 707708
rect 587572 706832 587808 707068
rect 587892 706832 588128 707068
rect 587572 706512 587808 706748
rect 587892 706512 588128 706748
rect 582326 705872 582562 706108
rect 582646 705872 582882 706108
rect 582326 705552 582562 705788
rect 582646 705552 582882 705788
rect 586612 705872 586848 706108
rect 586932 705872 587168 706108
rect 586612 705552 586848 705788
rect 586932 705552 587168 705788
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585652 704912 585888 705148
rect 585972 704912 586208 705148
rect 585652 704592 585888 704828
rect 585972 704592 586208 704828
rect 585652 687218 585888 687454
rect 585972 687218 586208 687454
rect 585652 686898 585888 687134
rect 585972 686898 586208 687134
rect 585652 651218 585888 651454
rect 585972 651218 586208 651454
rect 585652 650898 585888 651134
rect 585972 650898 586208 651134
rect 585652 615218 585888 615454
rect 585972 615218 586208 615454
rect 585652 614898 585888 615134
rect 585972 614898 586208 615134
rect 585652 579218 585888 579454
rect 585972 579218 586208 579454
rect 585652 578898 585888 579134
rect 585972 578898 586208 579134
rect 585652 543218 585888 543454
rect 585972 543218 586208 543454
rect 585652 542898 585888 543134
rect 585972 542898 586208 543134
rect 585652 507218 585888 507454
rect 585972 507218 586208 507454
rect 585652 506898 585888 507134
rect 585972 506898 586208 507134
rect 585652 471218 585888 471454
rect 585972 471218 586208 471454
rect 585652 470898 585888 471134
rect 585972 470898 586208 471134
rect 585652 435218 585888 435454
rect 585972 435218 586208 435454
rect 585652 434898 585888 435134
rect 585972 434898 586208 435134
rect 585652 399218 585888 399454
rect 585972 399218 586208 399454
rect 585652 398898 585888 399134
rect 585972 398898 586208 399134
rect 585652 363218 585888 363454
rect 585972 363218 586208 363454
rect 585652 362898 585888 363134
rect 585972 362898 586208 363134
rect 585652 327218 585888 327454
rect 585972 327218 586208 327454
rect 585652 326898 585888 327134
rect 585972 326898 586208 327134
rect 585652 291218 585888 291454
rect 585972 291218 586208 291454
rect 585652 290898 585888 291134
rect 585972 290898 586208 291134
rect 585652 255218 585888 255454
rect 585972 255218 586208 255454
rect 585652 254898 585888 255134
rect 585972 254898 586208 255134
rect 585652 219218 585888 219454
rect 585972 219218 586208 219454
rect 585652 218898 585888 219134
rect 585972 218898 586208 219134
rect 585652 183218 585888 183454
rect 585972 183218 586208 183454
rect 585652 182898 585888 183134
rect 585972 182898 586208 183134
rect 585652 147218 585888 147454
rect 585972 147218 586208 147454
rect 585652 146898 585888 147134
rect 585972 146898 586208 147134
rect 585652 111218 585888 111454
rect 585972 111218 586208 111454
rect 585652 110898 585888 111134
rect 585972 110898 586208 111134
rect 585652 75218 585888 75454
rect 585972 75218 586208 75454
rect 585652 74898 585888 75134
rect 585972 74898 586208 75134
rect 585652 39218 585888 39454
rect 585972 39218 586208 39454
rect 585652 38898 585888 39134
rect 585972 38898 586208 39134
rect 585652 3218 585888 3454
rect 585972 3218 586208 3454
rect 585652 2898 585888 3134
rect 585972 2898 586208 3134
rect 585652 -892 585888 -656
rect 585972 -892 586208 -656
rect 585652 -1212 585888 -976
rect 585972 -1212 586208 -976
rect 586612 691718 586848 691954
rect 586932 691718 587168 691954
rect 586612 691398 586848 691634
rect 586932 691398 587168 691634
rect 586612 655718 586848 655954
rect 586932 655718 587168 655954
rect 586612 655398 586848 655634
rect 586932 655398 587168 655634
rect 586612 619718 586848 619954
rect 586932 619718 587168 619954
rect 586612 619398 586848 619634
rect 586932 619398 587168 619634
rect 586612 583718 586848 583954
rect 586932 583718 587168 583954
rect 586612 583398 586848 583634
rect 586932 583398 587168 583634
rect 586612 547718 586848 547954
rect 586932 547718 587168 547954
rect 586612 547398 586848 547634
rect 586932 547398 587168 547634
rect 586612 511718 586848 511954
rect 586932 511718 587168 511954
rect 586612 511398 586848 511634
rect 586932 511398 587168 511634
rect 586612 475718 586848 475954
rect 586932 475718 587168 475954
rect 586612 475398 586848 475634
rect 586932 475398 587168 475634
rect 586612 439718 586848 439954
rect 586932 439718 587168 439954
rect 586612 439398 586848 439634
rect 586932 439398 587168 439634
rect 586612 403718 586848 403954
rect 586932 403718 587168 403954
rect 586612 403398 586848 403634
rect 586932 403398 587168 403634
rect 586612 367718 586848 367954
rect 586932 367718 587168 367954
rect 586612 367398 586848 367634
rect 586932 367398 587168 367634
rect 586612 331718 586848 331954
rect 586932 331718 587168 331954
rect 586612 331398 586848 331634
rect 586932 331398 587168 331634
rect 586612 295718 586848 295954
rect 586932 295718 587168 295954
rect 586612 295398 586848 295634
rect 586932 295398 587168 295634
rect 586612 259718 586848 259954
rect 586932 259718 587168 259954
rect 586612 259398 586848 259634
rect 586932 259398 587168 259634
rect 586612 223718 586848 223954
rect 586932 223718 587168 223954
rect 586612 223398 586848 223634
rect 586932 223398 587168 223634
rect 586612 187718 586848 187954
rect 586932 187718 587168 187954
rect 586612 187398 586848 187634
rect 586932 187398 587168 187634
rect 586612 151718 586848 151954
rect 586932 151718 587168 151954
rect 586612 151398 586848 151634
rect 586932 151398 587168 151634
rect 586612 115718 586848 115954
rect 586932 115718 587168 115954
rect 586612 115398 586848 115634
rect 586932 115398 587168 115634
rect 586612 79718 586848 79954
rect 586932 79718 587168 79954
rect 586612 79398 586848 79634
rect 586932 79398 587168 79634
rect 586612 43718 586848 43954
rect 586932 43718 587168 43954
rect 586612 43398 586848 43634
rect 586932 43398 587168 43634
rect 586612 7718 586848 7954
rect 586932 7718 587168 7954
rect 586612 7398 586848 7634
rect 586932 7398 587168 7634
rect 582326 -1852 582562 -1616
rect 582646 -1852 582882 -1616
rect 582326 -2172 582562 -1936
rect 582646 -2172 582882 -1936
rect 586612 -1852 586848 -1616
rect 586932 -1852 587168 -1616
rect 586612 -2172 586848 -1936
rect 586932 -2172 587168 -1936
rect 587572 696218 587808 696454
rect 587892 696218 588128 696454
rect 587572 695898 587808 696134
rect 587892 695898 588128 696134
rect 587572 660218 587808 660454
rect 587892 660218 588128 660454
rect 587572 659898 587808 660134
rect 587892 659898 588128 660134
rect 587572 624218 587808 624454
rect 587892 624218 588128 624454
rect 587572 623898 587808 624134
rect 587892 623898 588128 624134
rect 587572 588218 587808 588454
rect 587892 588218 588128 588454
rect 587572 587898 587808 588134
rect 587892 587898 588128 588134
rect 587572 552218 587808 552454
rect 587892 552218 588128 552454
rect 587572 551898 587808 552134
rect 587892 551898 588128 552134
rect 587572 516218 587808 516454
rect 587892 516218 588128 516454
rect 587572 515898 587808 516134
rect 587892 515898 588128 516134
rect 587572 480218 587808 480454
rect 587892 480218 588128 480454
rect 587572 479898 587808 480134
rect 587892 479898 588128 480134
rect 587572 444218 587808 444454
rect 587892 444218 588128 444454
rect 587572 443898 587808 444134
rect 587892 443898 588128 444134
rect 587572 408218 587808 408454
rect 587892 408218 588128 408454
rect 587572 407898 587808 408134
rect 587892 407898 588128 408134
rect 587572 372218 587808 372454
rect 587892 372218 588128 372454
rect 587572 371898 587808 372134
rect 587892 371898 588128 372134
rect 587572 336218 587808 336454
rect 587892 336218 588128 336454
rect 587572 335898 587808 336134
rect 587892 335898 588128 336134
rect 587572 300218 587808 300454
rect 587892 300218 588128 300454
rect 587572 299898 587808 300134
rect 587892 299898 588128 300134
rect 587572 264218 587808 264454
rect 587892 264218 588128 264454
rect 587572 263898 587808 264134
rect 587892 263898 588128 264134
rect 587572 228218 587808 228454
rect 587892 228218 588128 228454
rect 587572 227898 587808 228134
rect 587892 227898 588128 228134
rect 587572 192218 587808 192454
rect 587892 192218 588128 192454
rect 587572 191898 587808 192134
rect 587892 191898 588128 192134
rect 587572 156218 587808 156454
rect 587892 156218 588128 156454
rect 587572 155898 587808 156134
rect 587892 155898 588128 156134
rect 587572 120218 587808 120454
rect 587892 120218 588128 120454
rect 587572 119898 587808 120134
rect 587892 119898 588128 120134
rect 587572 84218 587808 84454
rect 587892 84218 588128 84454
rect 587572 83898 587808 84134
rect 587892 83898 588128 84134
rect 587572 48218 587808 48454
rect 587892 48218 588128 48454
rect 587572 47898 587808 48134
rect 587892 47898 588128 48134
rect 587572 12218 587808 12454
rect 587892 12218 588128 12454
rect 587572 11898 587808 12134
rect 587892 11898 588128 12134
rect 587572 -2812 587808 -2576
rect 587892 -2812 588128 -2576
rect 587572 -3132 587808 -2896
rect 587892 -3132 588128 -2896
rect 588532 700718 588768 700954
rect 588852 700718 589088 700954
rect 588532 700398 588768 700634
rect 588852 700398 589088 700634
rect 588532 664718 588768 664954
rect 588852 664718 589088 664954
rect 588532 664398 588768 664634
rect 588852 664398 589088 664634
rect 588532 628718 588768 628954
rect 588852 628718 589088 628954
rect 588532 628398 588768 628634
rect 588852 628398 589088 628634
rect 588532 592718 588768 592954
rect 588852 592718 589088 592954
rect 588532 592398 588768 592634
rect 588852 592398 589088 592634
rect 588532 556718 588768 556954
rect 588852 556718 589088 556954
rect 588532 556398 588768 556634
rect 588852 556398 589088 556634
rect 588532 520718 588768 520954
rect 588852 520718 589088 520954
rect 588532 520398 588768 520634
rect 588852 520398 589088 520634
rect 588532 484718 588768 484954
rect 588852 484718 589088 484954
rect 588532 484398 588768 484634
rect 588852 484398 589088 484634
rect 588532 448718 588768 448954
rect 588852 448718 589088 448954
rect 588532 448398 588768 448634
rect 588852 448398 589088 448634
rect 588532 412718 588768 412954
rect 588852 412718 589088 412954
rect 588532 412398 588768 412634
rect 588852 412398 589088 412634
rect 588532 376718 588768 376954
rect 588852 376718 589088 376954
rect 588532 376398 588768 376634
rect 588852 376398 589088 376634
rect 588532 340718 588768 340954
rect 588852 340718 589088 340954
rect 588532 340398 588768 340634
rect 588852 340398 589088 340634
rect 588532 304718 588768 304954
rect 588852 304718 589088 304954
rect 588532 304398 588768 304634
rect 588852 304398 589088 304634
rect 588532 268718 588768 268954
rect 588852 268718 589088 268954
rect 588532 268398 588768 268634
rect 588852 268398 589088 268634
rect 588532 232718 588768 232954
rect 588852 232718 589088 232954
rect 588532 232398 588768 232634
rect 588852 232398 589088 232634
rect 588532 196718 588768 196954
rect 588852 196718 589088 196954
rect 588532 196398 588768 196634
rect 588852 196398 589088 196634
rect 588532 160718 588768 160954
rect 588852 160718 589088 160954
rect 588532 160398 588768 160634
rect 588852 160398 589088 160634
rect 588532 124718 588768 124954
rect 588852 124718 589088 124954
rect 588532 124398 588768 124634
rect 588852 124398 589088 124634
rect 588532 88718 588768 88954
rect 588852 88718 589088 88954
rect 588532 88398 588768 88634
rect 588852 88398 589088 88634
rect 588532 52718 588768 52954
rect 588852 52718 589088 52954
rect 588532 52398 588768 52634
rect 588852 52398 589088 52634
rect 588532 16718 588768 16954
rect 588852 16718 589088 16954
rect 588532 16398 588768 16634
rect 588852 16398 589088 16634
rect 588532 -3772 588768 -3536
rect 588852 -3772 589088 -3536
rect 588532 -4092 588768 -3856
rect 588852 -4092 589088 -3856
rect 589492 669218 589728 669454
rect 589812 669218 590048 669454
rect 589492 668898 589728 669134
rect 589812 668898 590048 669134
rect 589492 633218 589728 633454
rect 589812 633218 590048 633454
rect 589492 632898 589728 633134
rect 589812 632898 590048 633134
rect 589492 597218 589728 597454
rect 589812 597218 590048 597454
rect 589492 596898 589728 597134
rect 589812 596898 590048 597134
rect 589492 561218 589728 561454
rect 589812 561218 590048 561454
rect 589492 560898 589728 561134
rect 589812 560898 590048 561134
rect 589492 525218 589728 525454
rect 589812 525218 590048 525454
rect 589492 524898 589728 525134
rect 589812 524898 590048 525134
rect 589492 489218 589728 489454
rect 589812 489218 590048 489454
rect 589492 488898 589728 489134
rect 589812 488898 590048 489134
rect 589492 453218 589728 453454
rect 589812 453218 590048 453454
rect 589492 452898 589728 453134
rect 589812 452898 590048 453134
rect 589492 417218 589728 417454
rect 589812 417218 590048 417454
rect 589492 416898 589728 417134
rect 589812 416898 590048 417134
rect 589492 381218 589728 381454
rect 589812 381218 590048 381454
rect 589492 380898 589728 381134
rect 589812 380898 590048 381134
rect 589492 345218 589728 345454
rect 589812 345218 590048 345454
rect 589492 344898 589728 345134
rect 589812 344898 590048 345134
rect 589492 309218 589728 309454
rect 589812 309218 590048 309454
rect 589492 308898 589728 309134
rect 589812 308898 590048 309134
rect 589492 273218 589728 273454
rect 589812 273218 590048 273454
rect 589492 272898 589728 273134
rect 589812 272898 590048 273134
rect 589492 237218 589728 237454
rect 589812 237218 590048 237454
rect 589492 236898 589728 237134
rect 589812 236898 590048 237134
rect 589492 201218 589728 201454
rect 589812 201218 590048 201454
rect 589492 200898 589728 201134
rect 589812 200898 590048 201134
rect 589492 165218 589728 165454
rect 589812 165218 590048 165454
rect 589492 164898 589728 165134
rect 589812 164898 590048 165134
rect 589492 129218 589728 129454
rect 589812 129218 590048 129454
rect 589492 128898 589728 129134
rect 589812 128898 590048 129134
rect 589492 93218 589728 93454
rect 589812 93218 590048 93454
rect 589492 92898 589728 93134
rect 589812 92898 590048 93134
rect 589492 57218 589728 57454
rect 589812 57218 590048 57454
rect 589492 56898 589728 57134
rect 589812 56898 590048 57134
rect 589492 21218 589728 21454
rect 589812 21218 590048 21454
rect 589492 20898 589728 21134
rect 589812 20898 590048 21134
rect 589492 -4732 589728 -4496
rect 589812 -4732 590048 -4496
rect 589492 -5052 589728 -4816
rect 589812 -5052 590048 -4816
rect 590452 673718 590688 673954
rect 590772 673718 591008 673954
rect 590452 673398 590688 673634
rect 590772 673398 591008 673634
rect 590452 637718 590688 637954
rect 590772 637718 591008 637954
rect 590452 637398 590688 637634
rect 590772 637398 591008 637634
rect 590452 601718 590688 601954
rect 590772 601718 591008 601954
rect 590452 601398 590688 601634
rect 590772 601398 591008 601634
rect 590452 565718 590688 565954
rect 590772 565718 591008 565954
rect 590452 565398 590688 565634
rect 590772 565398 591008 565634
rect 590452 529718 590688 529954
rect 590772 529718 591008 529954
rect 590452 529398 590688 529634
rect 590772 529398 591008 529634
rect 590452 493718 590688 493954
rect 590772 493718 591008 493954
rect 590452 493398 590688 493634
rect 590772 493398 591008 493634
rect 590452 457718 590688 457954
rect 590772 457718 591008 457954
rect 590452 457398 590688 457634
rect 590772 457398 591008 457634
rect 590452 421718 590688 421954
rect 590772 421718 591008 421954
rect 590452 421398 590688 421634
rect 590772 421398 591008 421634
rect 590452 385718 590688 385954
rect 590772 385718 591008 385954
rect 590452 385398 590688 385634
rect 590772 385398 591008 385634
rect 590452 349718 590688 349954
rect 590772 349718 591008 349954
rect 590452 349398 590688 349634
rect 590772 349398 591008 349634
rect 590452 313718 590688 313954
rect 590772 313718 591008 313954
rect 590452 313398 590688 313634
rect 590772 313398 591008 313634
rect 590452 277718 590688 277954
rect 590772 277718 591008 277954
rect 590452 277398 590688 277634
rect 590772 277398 591008 277634
rect 590452 241718 590688 241954
rect 590772 241718 591008 241954
rect 590452 241398 590688 241634
rect 590772 241398 591008 241634
rect 590452 205718 590688 205954
rect 590772 205718 591008 205954
rect 590452 205398 590688 205634
rect 590772 205398 591008 205634
rect 590452 169718 590688 169954
rect 590772 169718 591008 169954
rect 590452 169398 590688 169634
rect 590772 169398 591008 169634
rect 590452 133718 590688 133954
rect 590772 133718 591008 133954
rect 590452 133398 590688 133634
rect 590772 133398 591008 133634
rect 590452 97718 590688 97954
rect 590772 97718 591008 97954
rect 590452 97398 590688 97634
rect 590772 97398 591008 97634
rect 590452 61718 590688 61954
rect 590772 61718 591008 61954
rect 590452 61398 590688 61634
rect 590772 61398 591008 61634
rect 590452 25718 590688 25954
rect 590772 25718 591008 25954
rect 590452 25398 590688 25634
rect 590772 25398 591008 25634
rect 590452 -5692 590688 -5456
rect 590772 -5692 591008 -5456
rect 590452 -6012 590688 -5776
rect 590772 -6012 591008 -5776
rect 591412 678218 591648 678454
rect 591732 678218 591968 678454
rect 591412 677898 591648 678134
rect 591732 677898 591968 678134
rect 591412 642218 591648 642454
rect 591732 642218 591968 642454
rect 591412 641898 591648 642134
rect 591732 641898 591968 642134
rect 591412 606218 591648 606454
rect 591732 606218 591968 606454
rect 591412 605898 591648 606134
rect 591732 605898 591968 606134
rect 591412 570218 591648 570454
rect 591732 570218 591968 570454
rect 591412 569898 591648 570134
rect 591732 569898 591968 570134
rect 591412 534218 591648 534454
rect 591732 534218 591968 534454
rect 591412 533898 591648 534134
rect 591732 533898 591968 534134
rect 591412 498218 591648 498454
rect 591732 498218 591968 498454
rect 591412 497898 591648 498134
rect 591732 497898 591968 498134
rect 591412 462218 591648 462454
rect 591732 462218 591968 462454
rect 591412 461898 591648 462134
rect 591732 461898 591968 462134
rect 591412 426218 591648 426454
rect 591732 426218 591968 426454
rect 591412 425898 591648 426134
rect 591732 425898 591968 426134
rect 591412 390218 591648 390454
rect 591732 390218 591968 390454
rect 591412 389898 591648 390134
rect 591732 389898 591968 390134
rect 591412 354218 591648 354454
rect 591732 354218 591968 354454
rect 591412 353898 591648 354134
rect 591732 353898 591968 354134
rect 591412 318218 591648 318454
rect 591732 318218 591968 318454
rect 591412 317898 591648 318134
rect 591732 317898 591968 318134
rect 591412 282218 591648 282454
rect 591732 282218 591968 282454
rect 591412 281898 591648 282134
rect 591732 281898 591968 282134
rect 591412 246218 591648 246454
rect 591732 246218 591968 246454
rect 591412 245898 591648 246134
rect 591732 245898 591968 246134
rect 591412 210218 591648 210454
rect 591732 210218 591968 210454
rect 591412 209898 591648 210134
rect 591732 209898 591968 210134
rect 591412 174218 591648 174454
rect 591732 174218 591968 174454
rect 591412 173898 591648 174134
rect 591732 173898 591968 174134
rect 591412 138218 591648 138454
rect 591732 138218 591968 138454
rect 591412 137898 591648 138134
rect 591732 137898 591968 138134
rect 591412 102218 591648 102454
rect 591732 102218 591968 102454
rect 591412 101898 591648 102134
rect 591732 101898 591968 102134
rect 591412 66218 591648 66454
rect 591732 66218 591968 66454
rect 591412 65898 591648 66134
rect 591732 65898 591968 66134
rect 591412 30218 591648 30454
rect 591732 30218 591968 30454
rect 591412 29898 591648 30134
rect 591732 29898 591968 30134
rect 591412 -6652 591648 -6416
rect 591732 -6652 591968 -6416
rect 591412 -6972 591648 -6736
rect 591732 -6972 591968 -6736
rect 592372 682718 592608 682954
rect 592692 682718 592928 682954
rect 592372 682398 592608 682634
rect 592692 682398 592928 682634
rect 592372 646718 592608 646954
rect 592692 646718 592928 646954
rect 592372 646398 592608 646634
rect 592692 646398 592928 646634
rect 592372 610718 592608 610954
rect 592692 610718 592928 610954
rect 592372 610398 592608 610634
rect 592692 610398 592928 610634
rect 592372 574718 592608 574954
rect 592692 574718 592928 574954
rect 592372 574398 592608 574634
rect 592692 574398 592928 574634
rect 592372 538718 592608 538954
rect 592692 538718 592928 538954
rect 592372 538398 592608 538634
rect 592692 538398 592928 538634
rect 592372 502718 592608 502954
rect 592692 502718 592928 502954
rect 592372 502398 592608 502634
rect 592692 502398 592928 502634
rect 592372 466718 592608 466954
rect 592692 466718 592928 466954
rect 592372 466398 592608 466634
rect 592692 466398 592928 466634
rect 592372 430718 592608 430954
rect 592692 430718 592928 430954
rect 592372 430398 592608 430634
rect 592692 430398 592928 430634
rect 592372 394718 592608 394954
rect 592692 394718 592928 394954
rect 592372 394398 592608 394634
rect 592692 394398 592928 394634
rect 592372 358718 592608 358954
rect 592692 358718 592928 358954
rect 592372 358398 592608 358634
rect 592692 358398 592928 358634
rect 592372 322718 592608 322954
rect 592692 322718 592928 322954
rect 592372 322398 592608 322634
rect 592692 322398 592928 322634
rect 592372 286718 592608 286954
rect 592692 286718 592928 286954
rect 592372 286398 592608 286634
rect 592692 286398 592928 286634
rect 592372 250718 592608 250954
rect 592692 250718 592928 250954
rect 592372 250398 592608 250634
rect 592692 250398 592928 250634
rect 592372 214718 592608 214954
rect 592692 214718 592928 214954
rect 592372 214398 592608 214634
rect 592692 214398 592928 214634
rect 592372 178718 592608 178954
rect 592692 178718 592928 178954
rect 592372 178398 592608 178634
rect 592692 178398 592928 178634
rect 592372 142718 592608 142954
rect 592692 142718 592928 142954
rect 592372 142398 592608 142634
rect 592692 142398 592928 142634
rect 592372 106718 592608 106954
rect 592692 106718 592928 106954
rect 592372 106398 592608 106634
rect 592692 106398 592928 106634
rect 592372 70718 592608 70954
rect 592692 70718 592928 70954
rect 592372 70398 592608 70634
rect 592692 70398 592928 70634
rect 592372 34718 592608 34954
rect 592692 34718 592928 34954
rect 592372 34398 592608 34634
rect 592692 34398 592928 34634
rect 592372 -7612 592608 -7376
rect 592692 -7612 592928 -7376
rect 592372 -7932 592608 -7696
rect 592692 -7932 592928 -7696
<< metal5 >>
rect -9036 711868 592960 711900
rect -9036 711632 -9004 711868
rect -8768 711632 -8684 711868
rect -8448 711632 33326 711868
rect 33562 711632 33646 711868
rect 33882 711632 69326 711868
rect 69562 711632 69646 711868
rect 69882 711632 105326 711868
rect 105562 711632 105646 711868
rect 105882 711632 141326 711868
rect 141562 711632 141646 711868
rect 141882 711632 177326 711868
rect 177562 711632 177646 711868
rect 177882 711632 213326 711868
rect 213562 711632 213646 711868
rect 213882 711632 249326 711868
rect 249562 711632 249646 711868
rect 249882 711632 285326 711868
rect 285562 711632 285646 711868
rect 285882 711632 321326 711868
rect 321562 711632 321646 711868
rect 321882 711632 357326 711868
rect 357562 711632 357646 711868
rect 357882 711632 393326 711868
rect 393562 711632 393646 711868
rect 393882 711632 429326 711868
rect 429562 711632 429646 711868
rect 429882 711632 465326 711868
rect 465562 711632 465646 711868
rect 465882 711632 501326 711868
rect 501562 711632 501646 711868
rect 501882 711632 537326 711868
rect 537562 711632 537646 711868
rect 537882 711632 573326 711868
rect 573562 711632 573646 711868
rect 573882 711632 592372 711868
rect 592608 711632 592692 711868
rect 592928 711632 592960 711868
rect -9036 711548 592960 711632
rect -9036 711312 -9004 711548
rect -8768 711312 -8684 711548
rect -8448 711312 33326 711548
rect 33562 711312 33646 711548
rect 33882 711312 69326 711548
rect 69562 711312 69646 711548
rect 69882 711312 105326 711548
rect 105562 711312 105646 711548
rect 105882 711312 141326 711548
rect 141562 711312 141646 711548
rect 141882 711312 177326 711548
rect 177562 711312 177646 711548
rect 177882 711312 213326 711548
rect 213562 711312 213646 711548
rect 213882 711312 249326 711548
rect 249562 711312 249646 711548
rect 249882 711312 285326 711548
rect 285562 711312 285646 711548
rect 285882 711312 321326 711548
rect 321562 711312 321646 711548
rect 321882 711312 357326 711548
rect 357562 711312 357646 711548
rect 357882 711312 393326 711548
rect 393562 711312 393646 711548
rect 393882 711312 429326 711548
rect 429562 711312 429646 711548
rect 429882 711312 465326 711548
rect 465562 711312 465646 711548
rect 465882 711312 501326 711548
rect 501562 711312 501646 711548
rect 501882 711312 537326 711548
rect 537562 711312 537646 711548
rect 537882 711312 573326 711548
rect 573562 711312 573646 711548
rect 573882 711312 592372 711548
rect 592608 711312 592692 711548
rect 592928 711312 592960 711548
rect -9036 711280 592960 711312
rect -8076 710908 592000 710940
rect -8076 710672 -8044 710908
rect -7808 710672 -7724 710908
rect -7488 710672 28826 710908
rect 29062 710672 29146 710908
rect 29382 710672 64826 710908
rect 65062 710672 65146 710908
rect 65382 710672 100826 710908
rect 101062 710672 101146 710908
rect 101382 710672 136826 710908
rect 137062 710672 137146 710908
rect 137382 710672 172826 710908
rect 173062 710672 173146 710908
rect 173382 710672 208826 710908
rect 209062 710672 209146 710908
rect 209382 710672 244826 710908
rect 245062 710672 245146 710908
rect 245382 710672 280826 710908
rect 281062 710672 281146 710908
rect 281382 710672 316826 710908
rect 317062 710672 317146 710908
rect 317382 710672 352826 710908
rect 353062 710672 353146 710908
rect 353382 710672 388826 710908
rect 389062 710672 389146 710908
rect 389382 710672 424826 710908
rect 425062 710672 425146 710908
rect 425382 710672 460826 710908
rect 461062 710672 461146 710908
rect 461382 710672 496826 710908
rect 497062 710672 497146 710908
rect 497382 710672 532826 710908
rect 533062 710672 533146 710908
rect 533382 710672 568826 710908
rect 569062 710672 569146 710908
rect 569382 710672 591412 710908
rect 591648 710672 591732 710908
rect 591968 710672 592000 710908
rect -8076 710588 592000 710672
rect -8076 710352 -8044 710588
rect -7808 710352 -7724 710588
rect -7488 710352 28826 710588
rect 29062 710352 29146 710588
rect 29382 710352 64826 710588
rect 65062 710352 65146 710588
rect 65382 710352 100826 710588
rect 101062 710352 101146 710588
rect 101382 710352 136826 710588
rect 137062 710352 137146 710588
rect 137382 710352 172826 710588
rect 173062 710352 173146 710588
rect 173382 710352 208826 710588
rect 209062 710352 209146 710588
rect 209382 710352 244826 710588
rect 245062 710352 245146 710588
rect 245382 710352 280826 710588
rect 281062 710352 281146 710588
rect 281382 710352 316826 710588
rect 317062 710352 317146 710588
rect 317382 710352 352826 710588
rect 353062 710352 353146 710588
rect 353382 710352 388826 710588
rect 389062 710352 389146 710588
rect 389382 710352 424826 710588
rect 425062 710352 425146 710588
rect 425382 710352 460826 710588
rect 461062 710352 461146 710588
rect 461382 710352 496826 710588
rect 497062 710352 497146 710588
rect 497382 710352 532826 710588
rect 533062 710352 533146 710588
rect 533382 710352 568826 710588
rect 569062 710352 569146 710588
rect 569382 710352 591412 710588
rect 591648 710352 591732 710588
rect 591968 710352 592000 710588
rect -8076 710320 592000 710352
rect -7116 709948 591040 709980
rect -7116 709712 -7084 709948
rect -6848 709712 -6764 709948
rect -6528 709712 24326 709948
rect 24562 709712 24646 709948
rect 24882 709712 60326 709948
rect 60562 709712 60646 709948
rect 60882 709712 96326 709948
rect 96562 709712 96646 709948
rect 96882 709712 132326 709948
rect 132562 709712 132646 709948
rect 132882 709712 168326 709948
rect 168562 709712 168646 709948
rect 168882 709712 204326 709948
rect 204562 709712 204646 709948
rect 204882 709712 240326 709948
rect 240562 709712 240646 709948
rect 240882 709712 276326 709948
rect 276562 709712 276646 709948
rect 276882 709712 312326 709948
rect 312562 709712 312646 709948
rect 312882 709712 348326 709948
rect 348562 709712 348646 709948
rect 348882 709712 384326 709948
rect 384562 709712 384646 709948
rect 384882 709712 420326 709948
rect 420562 709712 420646 709948
rect 420882 709712 456326 709948
rect 456562 709712 456646 709948
rect 456882 709712 492326 709948
rect 492562 709712 492646 709948
rect 492882 709712 528326 709948
rect 528562 709712 528646 709948
rect 528882 709712 564326 709948
rect 564562 709712 564646 709948
rect 564882 709712 590452 709948
rect 590688 709712 590772 709948
rect 591008 709712 591040 709948
rect -7116 709628 591040 709712
rect -7116 709392 -7084 709628
rect -6848 709392 -6764 709628
rect -6528 709392 24326 709628
rect 24562 709392 24646 709628
rect 24882 709392 60326 709628
rect 60562 709392 60646 709628
rect 60882 709392 96326 709628
rect 96562 709392 96646 709628
rect 96882 709392 132326 709628
rect 132562 709392 132646 709628
rect 132882 709392 168326 709628
rect 168562 709392 168646 709628
rect 168882 709392 204326 709628
rect 204562 709392 204646 709628
rect 204882 709392 240326 709628
rect 240562 709392 240646 709628
rect 240882 709392 276326 709628
rect 276562 709392 276646 709628
rect 276882 709392 312326 709628
rect 312562 709392 312646 709628
rect 312882 709392 348326 709628
rect 348562 709392 348646 709628
rect 348882 709392 384326 709628
rect 384562 709392 384646 709628
rect 384882 709392 420326 709628
rect 420562 709392 420646 709628
rect 420882 709392 456326 709628
rect 456562 709392 456646 709628
rect 456882 709392 492326 709628
rect 492562 709392 492646 709628
rect 492882 709392 528326 709628
rect 528562 709392 528646 709628
rect 528882 709392 564326 709628
rect 564562 709392 564646 709628
rect 564882 709392 590452 709628
rect 590688 709392 590772 709628
rect 591008 709392 591040 709628
rect -7116 709360 591040 709392
rect -6156 708988 590080 709020
rect -6156 708752 -6124 708988
rect -5888 708752 -5804 708988
rect -5568 708752 19826 708988
rect 20062 708752 20146 708988
rect 20382 708752 55826 708988
rect 56062 708752 56146 708988
rect 56382 708752 91826 708988
rect 92062 708752 92146 708988
rect 92382 708752 127826 708988
rect 128062 708752 128146 708988
rect 128382 708752 163826 708988
rect 164062 708752 164146 708988
rect 164382 708752 199826 708988
rect 200062 708752 200146 708988
rect 200382 708752 235826 708988
rect 236062 708752 236146 708988
rect 236382 708752 271826 708988
rect 272062 708752 272146 708988
rect 272382 708752 307826 708988
rect 308062 708752 308146 708988
rect 308382 708752 343826 708988
rect 344062 708752 344146 708988
rect 344382 708752 379826 708988
rect 380062 708752 380146 708988
rect 380382 708752 415826 708988
rect 416062 708752 416146 708988
rect 416382 708752 451826 708988
rect 452062 708752 452146 708988
rect 452382 708752 487826 708988
rect 488062 708752 488146 708988
rect 488382 708752 523826 708988
rect 524062 708752 524146 708988
rect 524382 708752 559826 708988
rect 560062 708752 560146 708988
rect 560382 708752 589492 708988
rect 589728 708752 589812 708988
rect 590048 708752 590080 708988
rect -6156 708668 590080 708752
rect -6156 708432 -6124 708668
rect -5888 708432 -5804 708668
rect -5568 708432 19826 708668
rect 20062 708432 20146 708668
rect 20382 708432 55826 708668
rect 56062 708432 56146 708668
rect 56382 708432 91826 708668
rect 92062 708432 92146 708668
rect 92382 708432 127826 708668
rect 128062 708432 128146 708668
rect 128382 708432 163826 708668
rect 164062 708432 164146 708668
rect 164382 708432 199826 708668
rect 200062 708432 200146 708668
rect 200382 708432 235826 708668
rect 236062 708432 236146 708668
rect 236382 708432 271826 708668
rect 272062 708432 272146 708668
rect 272382 708432 307826 708668
rect 308062 708432 308146 708668
rect 308382 708432 343826 708668
rect 344062 708432 344146 708668
rect 344382 708432 379826 708668
rect 380062 708432 380146 708668
rect 380382 708432 415826 708668
rect 416062 708432 416146 708668
rect 416382 708432 451826 708668
rect 452062 708432 452146 708668
rect 452382 708432 487826 708668
rect 488062 708432 488146 708668
rect 488382 708432 523826 708668
rect 524062 708432 524146 708668
rect 524382 708432 559826 708668
rect 560062 708432 560146 708668
rect 560382 708432 589492 708668
rect 589728 708432 589812 708668
rect 590048 708432 590080 708668
rect -6156 708400 590080 708432
rect -5196 708028 589120 708060
rect -5196 707792 -5164 708028
rect -4928 707792 -4844 708028
rect -4608 707792 15326 708028
rect 15562 707792 15646 708028
rect 15882 707792 51326 708028
rect 51562 707792 51646 708028
rect 51882 707792 87326 708028
rect 87562 707792 87646 708028
rect 87882 707792 123326 708028
rect 123562 707792 123646 708028
rect 123882 707792 159326 708028
rect 159562 707792 159646 708028
rect 159882 707792 195326 708028
rect 195562 707792 195646 708028
rect 195882 707792 231326 708028
rect 231562 707792 231646 708028
rect 231882 707792 267326 708028
rect 267562 707792 267646 708028
rect 267882 707792 303326 708028
rect 303562 707792 303646 708028
rect 303882 707792 339326 708028
rect 339562 707792 339646 708028
rect 339882 707792 375326 708028
rect 375562 707792 375646 708028
rect 375882 707792 411326 708028
rect 411562 707792 411646 708028
rect 411882 707792 447326 708028
rect 447562 707792 447646 708028
rect 447882 707792 483326 708028
rect 483562 707792 483646 708028
rect 483882 707792 519326 708028
rect 519562 707792 519646 708028
rect 519882 707792 555326 708028
rect 555562 707792 555646 708028
rect 555882 707792 588532 708028
rect 588768 707792 588852 708028
rect 589088 707792 589120 708028
rect -5196 707708 589120 707792
rect -5196 707472 -5164 707708
rect -4928 707472 -4844 707708
rect -4608 707472 15326 707708
rect 15562 707472 15646 707708
rect 15882 707472 51326 707708
rect 51562 707472 51646 707708
rect 51882 707472 87326 707708
rect 87562 707472 87646 707708
rect 87882 707472 123326 707708
rect 123562 707472 123646 707708
rect 123882 707472 159326 707708
rect 159562 707472 159646 707708
rect 159882 707472 195326 707708
rect 195562 707472 195646 707708
rect 195882 707472 231326 707708
rect 231562 707472 231646 707708
rect 231882 707472 267326 707708
rect 267562 707472 267646 707708
rect 267882 707472 303326 707708
rect 303562 707472 303646 707708
rect 303882 707472 339326 707708
rect 339562 707472 339646 707708
rect 339882 707472 375326 707708
rect 375562 707472 375646 707708
rect 375882 707472 411326 707708
rect 411562 707472 411646 707708
rect 411882 707472 447326 707708
rect 447562 707472 447646 707708
rect 447882 707472 483326 707708
rect 483562 707472 483646 707708
rect 483882 707472 519326 707708
rect 519562 707472 519646 707708
rect 519882 707472 555326 707708
rect 555562 707472 555646 707708
rect 555882 707472 588532 707708
rect 588768 707472 588852 707708
rect 589088 707472 589120 707708
rect -5196 707440 589120 707472
rect -4236 707068 588160 707100
rect -4236 706832 -4204 707068
rect -3968 706832 -3884 707068
rect -3648 706832 10826 707068
rect 11062 706832 11146 707068
rect 11382 706832 46826 707068
rect 47062 706832 47146 707068
rect 47382 706832 82826 707068
rect 83062 706832 83146 707068
rect 83382 706832 118826 707068
rect 119062 706832 119146 707068
rect 119382 706832 154826 707068
rect 155062 706832 155146 707068
rect 155382 706832 190826 707068
rect 191062 706832 191146 707068
rect 191382 706832 226826 707068
rect 227062 706832 227146 707068
rect 227382 706832 262826 707068
rect 263062 706832 263146 707068
rect 263382 706832 298826 707068
rect 299062 706832 299146 707068
rect 299382 706832 334826 707068
rect 335062 706832 335146 707068
rect 335382 706832 370826 707068
rect 371062 706832 371146 707068
rect 371382 706832 406826 707068
rect 407062 706832 407146 707068
rect 407382 706832 442826 707068
rect 443062 706832 443146 707068
rect 443382 706832 478826 707068
rect 479062 706832 479146 707068
rect 479382 706832 514826 707068
rect 515062 706832 515146 707068
rect 515382 706832 550826 707068
rect 551062 706832 551146 707068
rect 551382 706832 587572 707068
rect 587808 706832 587892 707068
rect 588128 706832 588160 707068
rect -4236 706748 588160 706832
rect -4236 706512 -4204 706748
rect -3968 706512 -3884 706748
rect -3648 706512 10826 706748
rect 11062 706512 11146 706748
rect 11382 706512 46826 706748
rect 47062 706512 47146 706748
rect 47382 706512 82826 706748
rect 83062 706512 83146 706748
rect 83382 706512 118826 706748
rect 119062 706512 119146 706748
rect 119382 706512 154826 706748
rect 155062 706512 155146 706748
rect 155382 706512 190826 706748
rect 191062 706512 191146 706748
rect 191382 706512 226826 706748
rect 227062 706512 227146 706748
rect 227382 706512 262826 706748
rect 263062 706512 263146 706748
rect 263382 706512 298826 706748
rect 299062 706512 299146 706748
rect 299382 706512 334826 706748
rect 335062 706512 335146 706748
rect 335382 706512 370826 706748
rect 371062 706512 371146 706748
rect 371382 706512 406826 706748
rect 407062 706512 407146 706748
rect 407382 706512 442826 706748
rect 443062 706512 443146 706748
rect 443382 706512 478826 706748
rect 479062 706512 479146 706748
rect 479382 706512 514826 706748
rect 515062 706512 515146 706748
rect 515382 706512 550826 706748
rect 551062 706512 551146 706748
rect 551382 706512 587572 706748
rect 587808 706512 587892 706748
rect 588128 706512 588160 706748
rect -4236 706480 588160 706512
rect -3276 706108 587200 706140
rect -3276 705872 -3244 706108
rect -3008 705872 -2924 706108
rect -2688 705872 6326 706108
rect 6562 705872 6646 706108
rect 6882 705872 42326 706108
rect 42562 705872 42646 706108
rect 42882 705872 78326 706108
rect 78562 705872 78646 706108
rect 78882 705872 114326 706108
rect 114562 705872 114646 706108
rect 114882 705872 150326 706108
rect 150562 705872 150646 706108
rect 150882 705872 186326 706108
rect 186562 705872 186646 706108
rect 186882 705872 222326 706108
rect 222562 705872 222646 706108
rect 222882 705872 258326 706108
rect 258562 705872 258646 706108
rect 258882 705872 294326 706108
rect 294562 705872 294646 706108
rect 294882 705872 330326 706108
rect 330562 705872 330646 706108
rect 330882 705872 366326 706108
rect 366562 705872 366646 706108
rect 366882 705872 402326 706108
rect 402562 705872 402646 706108
rect 402882 705872 438326 706108
rect 438562 705872 438646 706108
rect 438882 705872 474326 706108
rect 474562 705872 474646 706108
rect 474882 705872 510326 706108
rect 510562 705872 510646 706108
rect 510882 705872 546326 706108
rect 546562 705872 546646 706108
rect 546882 705872 582326 706108
rect 582562 705872 582646 706108
rect 582882 705872 586612 706108
rect 586848 705872 586932 706108
rect 587168 705872 587200 706108
rect -3276 705788 587200 705872
rect -3276 705552 -3244 705788
rect -3008 705552 -2924 705788
rect -2688 705552 6326 705788
rect 6562 705552 6646 705788
rect 6882 705552 42326 705788
rect 42562 705552 42646 705788
rect 42882 705552 78326 705788
rect 78562 705552 78646 705788
rect 78882 705552 114326 705788
rect 114562 705552 114646 705788
rect 114882 705552 150326 705788
rect 150562 705552 150646 705788
rect 150882 705552 186326 705788
rect 186562 705552 186646 705788
rect 186882 705552 222326 705788
rect 222562 705552 222646 705788
rect 222882 705552 258326 705788
rect 258562 705552 258646 705788
rect 258882 705552 294326 705788
rect 294562 705552 294646 705788
rect 294882 705552 330326 705788
rect 330562 705552 330646 705788
rect 330882 705552 366326 705788
rect 366562 705552 366646 705788
rect 366882 705552 402326 705788
rect 402562 705552 402646 705788
rect 402882 705552 438326 705788
rect 438562 705552 438646 705788
rect 438882 705552 474326 705788
rect 474562 705552 474646 705788
rect 474882 705552 510326 705788
rect 510562 705552 510646 705788
rect 510882 705552 546326 705788
rect 546562 705552 546646 705788
rect 546882 705552 582326 705788
rect 582562 705552 582646 705788
rect 582882 705552 586612 705788
rect 586848 705552 586932 705788
rect 587168 705552 587200 705788
rect -3276 705520 587200 705552
rect -2316 705148 586240 705180
rect -2316 704912 -2284 705148
rect -2048 704912 -1964 705148
rect -1728 704912 1826 705148
rect 2062 704912 2146 705148
rect 2382 704912 37826 705148
rect 38062 704912 38146 705148
rect 38382 704912 73826 705148
rect 74062 704912 74146 705148
rect 74382 704912 109826 705148
rect 110062 704912 110146 705148
rect 110382 704912 145826 705148
rect 146062 704912 146146 705148
rect 146382 704912 181826 705148
rect 182062 704912 182146 705148
rect 182382 704912 217826 705148
rect 218062 704912 218146 705148
rect 218382 704912 253826 705148
rect 254062 704912 254146 705148
rect 254382 704912 289826 705148
rect 290062 704912 290146 705148
rect 290382 704912 325826 705148
rect 326062 704912 326146 705148
rect 326382 704912 361826 705148
rect 362062 704912 362146 705148
rect 362382 704912 397826 705148
rect 398062 704912 398146 705148
rect 398382 704912 433826 705148
rect 434062 704912 434146 705148
rect 434382 704912 469826 705148
rect 470062 704912 470146 705148
rect 470382 704912 505826 705148
rect 506062 704912 506146 705148
rect 506382 704912 541826 705148
rect 542062 704912 542146 705148
rect 542382 704912 577826 705148
rect 578062 704912 578146 705148
rect 578382 704912 585652 705148
rect 585888 704912 585972 705148
rect 586208 704912 586240 705148
rect -2316 704828 586240 704912
rect -2316 704592 -2284 704828
rect -2048 704592 -1964 704828
rect -1728 704592 1826 704828
rect 2062 704592 2146 704828
rect 2382 704592 37826 704828
rect 38062 704592 38146 704828
rect 38382 704592 73826 704828
rect 74062 704592 74146 704828
rect 74382 704592 109826 704828
rect 110062 704592 110146 704828
rect 110382 704592 145826 704828
rect 146062 704592 146146 704828
rect 146382 704592 181826 704828
rect 182062 704592 182146 704828
rect 182382 704592 217826 704828
rect 218062 704592 218146 704828
rect 218382 704592 253826 704828
rect 254062 704592 254146 704828
rect 254382 704592 289826 704828
rect 290062 704592 290146 704828
rect 290382 704592 325826 704828
rect 326062 704592 326146 704828
rect 326382 704592 361826 704828
rect 362062 704592 362146 704828
rect 362382 704592 397826 704828
rect 398062 704592 398146 704828
rect 398382 704592 433826 704828
rect 434062 704592 434146 704828
rect 434382 704592 469826 704828
rect 470062 704592 470146 704828
rect 470382 704592 505826 704828
rect 506062 704592 506146 704828
rect 506382 704592 541826 704828
rect 542062 704592 542146 704828
rect 542382 704592 577826 704828
rect 578062 704592 578146 704828
rect 578382 704592 585652 704828
rect 585888 704592 585972 704828
rect 586208 704592 586240 704828
rect -2316 704560 586240 704592
rect -9036 700954 592960 700986
rect -9036 700718 -5164 700954
rect -4928 700718 -4844 700954
rect -4608 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588532 700954
rect 588768 700718 588852 700954
rect 589088 700718 592960 700954
rect -9036 700634 592960 700718
rect -9036 700398 -5164 700634
rect -4928 700398 -4844 700634
rect -4608 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588532 700634
rect 588768 700398 588852 700634
rect 589088 700398 592960 700634
rect -9036 700366 592960 700398
rect -9036 696454 592960 696486
rect -9036 696218 -4204 696454
rect -3968 696218 -3884 696454
rect -3648 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587572 696454
rect 587808 696218 587892 696454
rect 588128 696218 592960 696454
rect -9036 696134 592960 696218
rect -9036 695898 -4204 696134
rect -3968 695898 -3884 696134
rect -3648 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587572 696134
rect 587808 695898 587892 696134
rect 588128 695898 592960 696134
rect -9036 695866 592960 695898
rect -9036 691954 592960 691986
rect -9036 691718 -3244 691954
rect -3008 691718 -2924 691954
rect -2688 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586612 691954
rect 586848 691718 586932 691954
rect 587168 691718 592960 691954
rect -9036 691634 592960 691718
rect -9036 691398 -3244 691634
rect -3008 691398 -2924 691634
rect -2688 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586612 691634
rect 586848 691398 586932 691634
rect 587168 691398 592960 691634
rect -9036 691366 592960 691398
rect -9036 687454 592960 687486
rect -9036 687218 -2284 687454
rect -2048 687218 -1964 687454
rect -1728 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585652 687454
rect 585888 687218 585972 687454
rect 586208 687218 592960 687454
rect -9036 687134 592960 687218
rect -9036 686898 -2284 687134
rect -2048 686898 -1964 687134
rect -1728 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585652 687134
rect 585888 686898 585972 687134
rect 586208 686898 592960 687134
rect -9036 686866 592960 686898
rect -9036 682954 592960 682986
rect -9036 682718 -9004 682954
rect -8768 682718 -8684 682954
rect -8448 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592372 682954
rect 592608 682718 592692 682954
rect 592928 682718 592960 682954
rect -9036 682634 592960 682718
rect -9036 682398 -9004 682634
rect -8768 682398 -8684 682634
rect -8448 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592372 682634
rect 592608 682398 592692 682634
rect 592928 682398 592960 682634
rect -9036 682366 592960 682398
rect -9036 678454 592960 678486
rect -9036 678218 -8044 678454
rect -7808 678218 -7724 678454
rect -7488 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591412 678454
rect 591648 678218 591732 678454
rect 591968 678218 592960 678454
rect -9036 678134 592960 678218
rect -9036 677898 -8044 678134
rect -7808 677898 -7724 678134
rect -7488 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591412 678134
rect 591648 677898 591732 678134
rect 591968 677898 592960 678134
rect -9036 677866 592960 677898
rect -9036 673954 592960 673986
rect -9036 673718 -7084 673954
rect -6848 673718 -6764 673954
rect -6528 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590452 673954
rect 590688 673718 590772 673954
rect 591008 673718 592960 673954
rect -9036 673634 592960 673718
rect -9036 673398 -7084 673634
rect -6848 673398 -6764 673634
rect -6528 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590452 673634
rect 590688 673398 590772 673634
rect 591008 673398 592960 673634
rect -9036 673366 592960 673398
rect -9036 669454 592960 669486
rect -9036 669218 -6124 669454
rect -5888 669218 -5804 669454
rect -5568 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589492 669454
rect 589728 669218 589812 669454
rect 590048 669218 592960 669454
rect -9036 669134 592960 669218
rect -9036 668898 -6124 669134
rect -5888 668898 -5804 669134
rect -5568 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589492 669134
rect 589728 668898 589812 669134
rect 590048 668898 592960 669134
rect -9036 668866 592960 668898
rect -9036 664954 592960 664986
rect -9036 664718 -5164 664954
rect -4928 664718 -4844 664954
rect -4608 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588532 664954
rect 588768 664718 588852 664954
rect 589088 664718 592960 664954
rect -9036 664634 592960 664718
rect -9036 664398 -5164 664634
rect -4928 664398 -4844 664634
rect -4608 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588532 664634
rect 588768 664398 588852 664634
rect 589088 664398 592960 664634
rect -9036 664366 592960 664398
rect -9036 660454 592960 660486
rect -9036 660218 -4204 660454
rect -3968 660218 -3884 660454
rect -3648 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587572 660454
rect 587808 660218 587892 660454
rect 588128 660218 592960 660454
rect -9036 660134 592960 660218
rect -9036 659898 -4204 660134
rect -3968 659898 -3884 660134
rect -3648 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587572 660134
rect 587808 659898 587892 660134
rect 588128 659898 592960 660134
rect -9036 659866 592960 659898
rect -9036 655954 592960 655986
rect -9036 655718 -3244 655954
rect -3008 655718 -2924 655954
rect -2688 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586612 655954
rect 586848 655718 586932 655954
rect 587168 655718 592960 655954
rect -9036 655634 592960 655718
rect -9036 655398 -3244 655634
rect -3008 655398 -2924 655634
rect -2688 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586612 655634
rect 586848 655398 586932 655634
rect 587168 655398 592960 655634
rect -9036 655366 592960 655398
rect -9036 651454 592960 651486
rect -9036 651218 -2284 651454
rect -2048 651218 -1964 651454
rect -1728 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585652 651454
rect 585888 651218 585972 651454
rect 586208 651218 592960 651454
rect -9036 651134 592960 651218
rect -9036 650898 -2284 651134
rect -2048 650898 -1964 651134
rect -1728 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585652 651134
rect 585888 650898 585972 651134
rect 586208 650898 592960 651134
rect -9036 650866 592960 650898
rect -9036 646954 592960 646986
rect -9036 646718 -9004 646954
rect -8768 646718 -8684 646954
rect -8448 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592372 646954
rect 592608 646718 592692 646954
rect 592928 646718 592960 646954
rect -9036 646634 592960 646718
rect -9036 646398 -9004 646634
rect -8768 646398 -8684 646634
rect -8448 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592372 646634
rect 592608 646398 592692 646634
rect 592928 646398 592960 646634
rect -9036 646366 592960 646398
rect -9036 642454 592960 642486
rect -9036 642218 -8044 642454
rect -7808 642218 -7724 642454
rect -7488 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591412 642454
rect 591648 642218 591732 642454
rect 591968 642218 592960 642454
rect -9036 642134 592960 642218
rect -9036 641898 -8044 642134
rect -7808 641898 -7724 642134
rect -7488 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591412 642134
rect 591648 641898 591732 642134
rect 591968 641898 592960 642134
rect -9036 641866 592960 641898
rect -9036 637954 592960 637986
rect -9036 637718 -7084 637954
rect -6848 637718 -6764 637954
rect -6528 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590452 637954
rect 590688 637718 590772 637954
rect 591008 637718 592960 637954
rect -9036 637634 592960 637718
rect -9036 637398 -7084 637634
rect -6848 637398 -6764 637634
rect -6528 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590452 637634
rect 590688 637398 590772 637634
rect 591008 637398 592960 637634
rect -9036 637366 592960 637398
rect -9036 633454 592960 633486
rect -9036 633218 -6124 633454
rect -5888 633218 -5804 633454
rect -5568 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589492 633454
rect 589728 633218 589812 633454
rect 590048 633218 592960 633454
rect -9036 633134 592960 633218
rect -9036 632898 -6124 633134
rect -5888 632898 -5804 633134
rect -5568 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589492 633134
rect 589728 632898 589812 633134
rect 590048 632898 592960 633134
rect -9036 632866 592960 632898
rect -9036 628954 592960 628986
rect -9036 628718 -5164 628954
rect -4928 628718 -4844 628954
rect -4608 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588532 628954
rect 588768 628718 588852 628954
rect 589088 628718 592960 628954
rect -9036 628634 592960 628718
rect -9036 628398 -5164 628634
rect -4928 628398 -4844 628634
rect -4608 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588532 628634
rect 588768 628398 588852 628634
rect 589088 628398 592960 628634
rect -9036 628366 592960 628398
rect -9036 624454 592960 624486
rect -9036 624218 -4204 624454
rect -3968 624218 -3884 624454
rect -3648 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587572 624454
rect 587808 624218 587892 624454
rect 588128 624218 592960 624454
rect -9036 624134 592960 624218
rect -9036 623898 -4204 624134
rect -3968 623898 -3884 624134
rect -3648 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587572 624134
rect 587808 623898 587892 624134
rect 588128 623898 592960 624134
rect -9036 623866 592960 623898
rect -9036 619954 592960 619986
rect -9036 619718 -3244 619954
rect -3008 619718 -2924 619954
rect -2688 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586612 619954
rect 586848 619718 586932 619954
rect 587168 619718 592960 619954
rect -9036 619634 592960 619718
rect -9036 619398 -3244 619634
rect -3008 619398 -2924 619634
rect -2688 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586612 619634
rect 586848 619398 586932 619634
rect 587168 619398 592960 619634
rect -9036 619366 592960 619398
rect -9036 615454 592960 615486
rect -9036 615218 -2284 615454
rect -2048 615218 -1964 615454
rect -1728 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585652 615454
rect 585888 615218 585972 615454
rect 586208 615218 592960 615454
rect -9036 615134 592960 615218
rect -9036 614898 -2284 615134
rect -2048 614898 -1964 615134
rect -1728 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585652 615134
rect 585888 614898 585972 615134
rect 586208 614898 592960 615134
rect -9036 614866 592960 614898
rect -9036 610954 592960 610986
rect -9036 610718 -9004 610954
rect -8768 610718 -8684 610954
rect -8448 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592372 610954
rect 592608 610718 592692 610954
rect 592928 610718 592960 610954
rect -9036 610634 592960 610718
rect -9036 610398 -9004 610634
rect -8768 610398 -8684 610634
rect -8448 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592372 610634
rect 592608 610398 592692 610634
rect 592928 610398 592960 610634
rect -9036 610366 592960 610398
rect -9036 606454 592960 606486
rect -9036 606218 -8044 606454
rect -7808 606218 -7724 606454
rect -7488 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591412 606454
rect 591648 606218 591732 606454
rect 591968 606218 592960 606454
rect -9036 606134 592960 606218
rect -9036 605898 -8044 606134
rect -7808 605898 -7724 606134
rect -7488 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591412 606134
rect 591648 605898 591732 606134
rect 591968 605898 592960 606134
rect -9036 605866 592960 605898
rect -9036 601954 592960 601986
rect -9036 601718 -7084 601954
rect -6848 601718 -6764 601954
rect -6528 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590452 601954
rect 590688 601718 590772 601954
rect 591008 601718 592960 601954
rect -9036 601634 592960 601718
rect -9036 601398 -7084 601634
rect -6848 601398 -6764 601634
rect -6528 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590452 601634
rect 590688 601398 590772 601634
rect 591008 601398 592960 601634
rect -9036 601366 592960 601398
rect -9036 597454 592960 597486
rect -9036 597218 -6124 597454
rect -5888 597218 -5804 597454
rect -5568 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589492 597454
rect 589728 597218 589812 597454
rect 590048 597218 592960 597454
rect -9036 597134 592960 597218
rect -9036 596898 -6124 597134
rect -5888 596898 -5804 597134
rect -5568 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589492 597134
rect 589728 596898 589812 597134
rect 590048 596898 592960 597134
rect -9036 596866 592960 596898
rect -9036 592954 592960 592986
rect -9036 592718 -5164 592954
rect -4928 592718 -4844 592954
rect -4608 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588532 592954
rect 588768 592718 588852 592954
rect 589088 592718 592960 592954
rect -9036 592634 592960 592718
rect -9036 592398 -5164 592634
rect -4928 592398 -4844 592634
rect -4608 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588532 592634
rect 588768 592398 588852 592634
rect 589088 592398 592960 592634
rect -9036 592366 592960 592398
rect -9036 588454 592960 588486
rect -9036 588218 -4204 588454
rect -3968 588218 -3884 588454
rect -3648 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587572 588454
rect 587808 588218 587892 588454
rect 588128 588218 592960 588454
rect -9036 588134 592960 588218
rect -9036 587898 -4204 588134
rect -3968 587898 -3884 588134
rect -3648 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587572 588134
rect 587808 587898 587892 588134
rect 588128 587898 592960 588134
rect -9036 587866 592960 587898
rect -9036 583954 592960 583986
rect -9036 583718 -3244 583954
rect -3008 583718 -2924 583954
rect -2688 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586612 583954
rect 586848 583718 586932 583954
rect 587168 583718 592960 583954
rect -9036 583634 592960 583718
rect -9036 583398 -3244 583634
rect -3008 583398 -2924 583634
rect -2688 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586612 583634
rect 586848 583398 586932 583634
rect 587168 583398 592960 583634
rect -9036 583366 592960 583398
rect -9036 579454 592960 579486
rect -9036 579218 -2284 579454
rect -2048 579218 -1964 579454
rect -1728 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585652 579454
rect 585888 579218 585972 579454
rect 586208 579218 592960 579454
rect -9036 579134 592960 579218
rect -9036 578898 -2284 579134
rect -2048 578898 -1964 579134
rect -1728 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585652 579134
rect 585888 578898 585972 579134
rect 586208 578898 592960 579134
rect -9036 578866 592960 578898
rect -9036 574954 592960 574986
rect -9036 574718 -9004 574954
rect -8768 574718 -8684 574954
rect -8448 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592372 574954
rect 592608 574718 592692 574954
rect 592928 574718 592960 574954
rect -9036 574634 592960 574718
rect -9036 574398 -9004 574634
rect -8768 574398 -8684 574634
rect -8448 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592372 574634
rect 592608 574398 592692 574634
rect 592928 574398 592960 574634
rect -9036 574366 592960 574398
rect -9036 570454 592960 570486
rect -9036 570218 -8044 570454
rect -7808 570218 -7724 570454
rect -7488 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591412 570454
rect 591648 570218 591732 570454
rect 591968 570218 592960 570454
rect -9036 570134 592960 570218
rect -9036 569898 -8044 570134
rect -7808 569898 -7724 570134
rect -7488 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591412 570134
rect 591648 569898 591732 570134
rect 591968 569898 592960 570134
rect -9036 569866 592960 569898
rect -9036 565954 592960 565986
rect -9036 565718 -7084 565954
rect -6848 565718 -6764 565954
rect -6528 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590452 565954
rect 590688 565718 590772 565954
rect 591008 565718 592960 565954
rect -9036 565634 592960 565718
rect -9036 565398 -7084 565634
rect -6848 565398 -6764 565634
rect -6528 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590452 565634
rect 590688 565398 590772 565634
rect 591008 565398 592960 565634
rect -9036 565366 592960 565398
rect -9036 561454 592960 561486
rect -9036 561218 -6124 561454
rect -5888 561218 -5804 561454
rect -5568 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589492 561454
rect 589728 561218 589812 561454
rect 590048 561218 592960 561454
rect -9036 561134 592960 561218
rect -9036 560898 -6124 561134
rect -5888 560898 -5804 561134
rect -5568 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589492 561134
rect 589728 560898 589812 561134
rect 590048 560898 592960 561134
rect -9036 560866 592960 560898
rect -9036 556954 592960 556986
rect -9036 556718 -5164 556954
rect -4928 556718 -4844 556954
rect -4608 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588532 556954
rect 588768 556718 588852 556954
rect 589088 556718 592960 556954
rect -9036 556634 592960 556718
rect -9036 556398 -5164 556634
rect -4928 556398 -4844 556634
rect -4608 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588532 556634
rect 588768 556398 588852 556634
rect 589088 556398 592960 556634
rect -9036 556366 592960 556398
rect -9036 552454 592960 552486
rect -9036 552218 -4204 552454
rect -3968 552218 -3884 552454
rect -3648 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587572 552454
rect 587808 552218 587892 552454
rect 588128 552218 592960 552454
rect -9036 552134 592960 552218
rect -9036 551898 -4204 552134
rect -3968 551898 -3884 552134
rect -3648 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587572 552134
rect 587808 551898 587892 552134
rect 588128 551898 592960 552134
rect -9036 551866 592960 551898
rect -9036 547954 592960 547986
rect -9036 547718 -3244 547954
rect -3008 547718 -2924 547954
rect -2688 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 220328 547954
rect 220564 547718 356056 547954
rect 356292 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586612 547954
rect 586848 547718 586932 547954
rect 587168 547718 592960 547954
rect -9036 547634 592960 547718
rect -9036 547398 -3244 547634
rect -3008 547398 -2924 547634
rect -2688 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 220328 547634
rect 220564 547398 356056 547634
rect 356292 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586612 547634
rect 586848 547398 586932 547634
rect 587168 547398 592960 547634
rect -9036 547366 592960 547398
rect -9036 543454 592960 543486
rect -9036 543218 -2284 543454
rect -2048 543218 -1964 543454
rect -1728 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 221008 543454
rect 221244 543218 355376 543454
rect 355612 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585652 543454
rect 585888 543218 585972 543454
rect 586208 543218 592960 543454
rect -9036 543134 592960 543218
rect -9036 542898 -2284 543134
rect -2048 542898 -1964 543134
rect -1728 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 221008 543134
rect 221244 542898 355376 543134
rect 355612 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585652 543134
rect 585888 542898 585972 543134
rect 586208 542898 592960 543134
rect -9036 542866 592960 542898
rect -9036 538954 592960 538986
rect -9036 538718 -9004 538954
rect -8768 538718 -8684 538954
rect -8448 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592372 538954
rect 592608 538718 592692 538954
rect 592928 538718 592960 538954
rect -9036 538634 592960 538718
rect -9036 538398 -9004 538634
rect -8768 538398 -8684 538634
rect -8448 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592372 538634
rect 592608 538398 592692 538634
rect 592928 538398 592960 538634
rect -9036 538366 592960 538398
rect -9036 534454 592960 534486
rect -9036 534218 -8044 534454
rect -7808 534218 -7724 534454
rect -7488 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591412 534454
rect 591648 534218 591732 534454
rect 591968 534218 592960 534454
rect -9036 534134 592960 534218
rect -9036 533898 -8044 534134
rect -7808 533898 -7724 534134
rect -7488 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591412 534134
rect 591648 533898 591732 534134
rect 591968 533898 592960 534134
rect -9036 533866 592960 533898
rect -9036 529954 592960 529986
rect -9036 529718 -7084 529954
rect -6848 529718 -6764 529954
rect -6528 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590452 529954
rect 590688 529718 590772 529954
rect 591008 529718 592960 529954
rect -9036 529634 592960 529718
rect -9036 529398 -7084 529634
rect -6848 529398 -6764 529634
rect -6528 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590452 529634
rect 590688 529398 590772 529634
rect 591008 529398 592960 529634
rect -9036 529366 592960 529398
rect -9036 525454 592960 525486
rect -9036 525218 -6124 525454
rect -5888 525218 -5804 525454
rect -5568 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589492 525454
rect 589728 525218 589812 525454
rect 590048 525218 592960 525454
rect -9036 525134 592960 525218
rect -9036 524898 -6124 525134
rect -5888 524898 -5804 525134
rect -5568 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589492 525134
rect 589728 524898 589812 525134
rect 590048 524898 592960 525134
rect -9036 524866 592960 524898
rect -9036 520954 592960 520986
rect -9036 520718 -5164 520954
rect -4928 520718 -4844 520954
rect -4608 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588532 520954
rect 588768 520718 588852 520954
rect 589088 520718 592960 520954
rect -9036 520634 592960 520718
rect -9036 520398 -5164 520634
rect -4928 520398 -4844 520634
rect -4608 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588532 520634
rect 588768 520398 588852 520634
rect 589088 520398 592960 520634
rect -9036 520366 592960 520398
rect -9036 516454 592960 516486
rect -9036 516218 -4204 516454
rect -3968 516218 -3884 516454
rect -3648 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587572 516454
rect 587808 516218 587892 516454
rect 588128 516218 592960 516454
rect -9036 516134 592960 516218
rect -9036 515898 -4204 516134
rect -3968 515898 -3884 516134
rect -3648 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587572 516134
rect 587808 515898 587892 516134
rect 588128 515898 592960 516134
rect -9036 515866 592960 515898
rect -9036 511954 592960 511986
rect -9036 511718 -3244 511954
rect -3008 511718 -2924 511954
rect -2688 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 220328 511954
rect 220564 511718 356056 511954
rect 356292 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586612 511954
rect 586848 511718 586932 511954
rect 587168 511718 592960 511954
rect -9036 511634 592960 511718
rect -9036 511398 -3244 511634
rect -3008 511398 -2924 511634
rect -2688 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 220328 511634
rect 220564 511398 356056 511634
rect 356292 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586612 511634
rect 586848 511398 586932 511634
rect 587168 511398 592960 511634
rect -9036 511366 592960 511398
rect -9036 507454 592960 507486
rect -9036 507218 -2284 507454
rect -2048 507218 -1964 507454
rect -1728 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 221008 507454
rect 221244 507218 355376 507454
rect 355612 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585652 507454
rect 585888 507218 585972 507454
rect 586208 507218 592960 507454
rect -9036 507134 592960 507218
rect -9036 506898 -2284 507134
rect -2048 506898 -1964 507134
rect -1728 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 221008 507134
rect 221244 506898 355376 507134
rect 355612 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585652 507134
rect 585888 506898 585972 507134
rect 586208 506898 592960 507134
rect -9036 506866 592960 506898
rect -9036 502954 592960 502986
rect -9036 502718 -9004 502954
rect -8768 502718 -8684 502954
rect -8448 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592372 502954
rect 592608 502718 592692 502954
rect 592928 502718 592960 502954
rect -9036 502634 592960 502718
rect -9036 502398 -9004 502634
rect -8768 502398 -8684 502634
rect -8448 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592372 502634
rect 592608 502398 592692 502634
rect 592928 502398 592960 502634
rect -9036 502366 592960 502398
rect -9036 498454 592960 498486
rect -9036 498218 -8044 498454
rect -7808 498218 -7724 498454
rect -7488 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591412 498454
rect 591648 498218 591732 498454
rect 591968 498218 592960 498454
rect -9036 498134 592960 498218
rect -9036 497898 -8044 498134
rect -7808 497898 -7724 498134
rect -7488 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591412 498134
rect 591648 497898 591732 498134
rect 591968 497898 592960 498134
rect -9036 497866 592960 497898
rect -9036 493954 592960 493986
rect -9036 493718 -7084 493954
rect -6848 493718 -6764 493954
rect -6528 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590452 493954
rect 590688 493718 590772 493954
rect 591008 493718 592960 493954
rect -9036 493634 592960 493718
rect -9036 493398 -7084 493634
rect -6848 493398 -6764 493634
rect -6528 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590452 493634
rect 590688 493398 590772 493634
rect 591008 493398 592960 493634
rect -9036 493366 592960 493398
rect -9036 489454 592960 489486
rect -9036 489218 -6124 489454
rect -5888 489218 -5804 489454
rect -5568 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589492 489454
rect 589728 489218 589812 489454
rect 590048 489218 592960 489454
rect -9036 489134 592960 489218
rect -9036 488898 -6124 489134
rect -5888 488898 -5804 489134
rect -5568 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589492 489134
rect 589728 488898 589812 489134
rect 590048 488898 592960 489134
rect -9036 488866 592960 488898
rect -9036 484954 592960 484986
rect -9036 484718 -5164 484954
rect -4928 484718 -4844 484954
rect -4608 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588532 484954
rect 588768 484718 588852 484954
rect 589088 484718 592960 484954
rect -9036 484634 592960 484718
rect -9036 484398 -5164 484634
rect -4928 484398 -4844 484634
rect -4608 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588532 484634
rect 588768 484398 588852 484634
rect 589088 484398 592960 484634
rect -9036 484366 592960 484398
rect -9036 480454 592960 480486
rect -9036 480218 -4204 480454
rect -3968 480218 -3884 480454
rect -3648 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587572 480454
rect 587808 480218 587892 480454
rect 588128 480218 592960 480454
rect -9036 480134 592960 480218
rect -9036 479898 -4204 480134
rect -3968 479898 -3884 480134
rect -3648 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587572 480134
rect 587808 479898 587892 480134
rect 588128 479898 592960 480134
rect -9036 479866 592960 479898
rect -9036 475954 592960 475986
rect -9036 475718 -3244 475954
rect -3008 475718 -2924 475954
rect -2688 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586612 475954
rect 586848 475718 586932 475954
rect 587168 475718 592960 475954
rect -9036 475634 592960 475718
rect -9036 475398 -3244 475634
rect -3008 475398 -2924 475634
rect -2688 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586612 475634
rect 586848 475398 586932 475634
rect 587168 475398 592960 475634
rect -9036 475366 592960 475398
rect -9036 471454 592960 471486
rect -9036 471218 -2284 471454
rect -2048 471218 -1964 471454
rect -1728 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585652 471454
rect 585888 471218 585972 471454
rect 586208 471218 592960 471454
rect -9036 471134 592960 471218
rect -9036 470898 -2284 471134
rect -2048 470898 -1964 471134
rect -1728 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585652 471134
rect 585888 470898 585972 471134
rect 586208 470898 592960 471134
rect -9036 470866 592960 470898
rect -9036 466954 592960 466986
rect -9036 466718 -9004 466954
rect -8768 466718 -8684 466954
rect -8448 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592372 466954
rect 592608 466718 592692 466954
rect 592928 466718 592960 466954
rect -9036 466634 592960 466718
rect -9036 466398 -9004 466634
rect -8768 466398 -8684 466634
rect -8448 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592372 466634
rect 592608 466398 592692 466634
rect 592928 466398 592960 466634
rect -9036 466366 592960 466398
rect -9036 462454 592960 462486
rect -9036 462218 -8044 462454
rect -7808 462218 -7724 462454
rect -7488 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591412 462454
rect 591648 462218 591732 462454
rect 591968 462218 592960 462454
rect -9036 462134 592960 462218
rect -9036 461898 -8044 462134
rect -7808 461898 -7724 462134
rect -7488 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591412 462134
rect 591648 461898 591732 462134
rect 591968 461898 592960 462134
rect -9036 461866 592960 461898
rect -9036 457954 592960 457986
rect -9036 457718 -7084 457954
rect -6848 457718 -6764 457954
rect -6528 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590452 457954
rect 590688 457718 590772 457954
rect 591008 457718 592960 457954
rect -9036 457634 592960 457718
rect -9036 457398 -7084 457634
rect -6848 457398 -6764 457634
rect -6528 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590452 457634
rect 590688 457398 590772 457634
rect 591008 457398 592960 457634
rect -9036 457366 592960 457398
rect -9036 453454 592960 453486
rect -9036 453218 -6124 453454
rect -5888 453218 -5804 453454
rect -5568 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589492 453454
rect 589728 453218 589812 453454
rect 590048 453218 592960 453454
rect -9036 453134 592960 453218
rect -9036 452898 -6124 453134
rect -5888 452898 -5804 453134
rect -5568 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589492 453134
rect 589728 452898 589812 453134
rect 590048 452898 592960 453134
rect -9036 452866 592960 452898
rect -9036 448954 592960 448986
rect -9036 448718 -5164 448954
rect -4928 448718 -4844 448954
rect -4608 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588532 448954
rect 588768 448718 588852 448954
rect 589088 448718 592960 448954
rect -9036 448634 592960 448718
rect -9036 448398 -5164 448634
rect -4928 448398 -4844 448634
rect -4608 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588532 448634
rect 588768 448398 588852 448634
rect 589088 448398 592960 448634
rect -9036 448366 592960 448398
rect -9036 444454 592960 444486
rect -9036 444218 -4204 444454
rect -3968 444218 -3884 444454
rect -3648 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587572 444454
rect 587808 444218 587892 444454
rect 588128 444218 592960 444454
rect -9036 444134 592960 444218
rect -9036 443898 -4204 444134
rect -3968 443898 -3884 444134
rect -3648 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587572 444134
rect 587808 443898 587892 444134
rect 588128 443898 592960 444134
rect -9036 443866 592960 443898
rect -9036 439954 592960 439986
rect -9036 439718 -3244 439954
rect -3008 439718 -2924 439954
rect -2688 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586612 439954
rect 586848 439718 586932 439954
rect 587168 439718 592960 439954
rect -9036 439634 592960 439718
rect -9036 439398 -3244 439634
rect -3008 439398 -2924 439634
rect -2688 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586612 439634
rect 586848 439398 586932 439634
rect 587168 439398 592960 439634
rect -9036 439366 592960 439398
rect -9036 435454 592960 435486
rect -9036 435218 -2284 435454
rect -2048 435218 -1964 435454
rect -1728 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 236650 435454
rect 236886 435218 267370 435454
rect 267606 435218 298090 435454
rect 298326 435218 328810 435454
rect 329046 435218 359530 435454
rect 359766 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585652 435454
rect 585888 435218 585972 435454
rect 586208 435218 592960 435454
rect -9036 435134 592960 435218
rect -9036 434898 -2284 435134
rect -2048 434898 -1964 435134
rect -1728 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 236650 435134
rect 236886 434898 267370 435134
rect 267606 434898 298090 435134
rect 298326 434898 328810 435134
rect 329046 434898 359530 435134
rect 359766 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585652 435134
rect 585888 434898 585972 435134
rect 586208 434898 592960 435134
rect -9036 434866 592960 434898
rect -9036 430954 592960 430986
rect -9036 430718 -9004 430954
rect -8768 430718 -8684 430954
rect -8448 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592372 430954
rect 592608 430718 592692 430954
rect 592928 430718 592960 430954
rect -9036 430634 592960 430718
rect -9036 430398 -9004 430634
rect -8768 430398 -8684 430634
rect -8448 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592372 430634
rect 592608 430398 592692 430634
rect 592928 430398 592960 430634
rect -9036 430366 592960 430398
rect -9036 426454 592960 426486
rect -9036 426218 -8044 426454
rect -7808 426218 -7724 426454
rect -7488 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591412 426454
rect 591648 426218 591732 426454
rect 591968 426218 592960 426454
rect -9036 426134 592960 426218
rect -9036 425898 -8044 426134
rect -7808 425898 -7724 426134
rect -7488 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591412 426134
rect 591648 425898 591732 426134
rect 591968 425898 592960 426134
rect -9036 425866 592960 425898
rect -9036 421954 592960 421986
rect -9036 421718 -7084 421954
rect -6848 421718 -6764 421954
rect -6528 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590452 421954
rect 590688 421718 590772 421954
rect 591008 421718 592960 421954
rect -9036 421634 592960 421718
rect -9036 421398 -7084 421634
rect -6848 421398 -6764 421634
rect -6528 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590452 421634
rect 590688 421398 590772 421634
rect 591008 421398 592960 421634
rect -9036 421366 592960 421398
rect -9036 417454 592960 417486
rect -9036 417218 -6124 417454
rect -5888 417218 -5804 417454
rect -5568 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589492 417454
rect 589728 417218 589812 417454
rect 590048 417218 592960 417454
rect -9036 417134 592960 417218
rect -9036 416898 -6124 417134
rect -5888 416898 -5804 417134
rect -5568 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589492 417134
rect 589728 416898 589812 417134
rect 590048 416898 592960 417134
rect -9036 416866 592960 416898
rect -9036 412954 592960 412986
rect -9036 412718 -5164 412954
rect -4928 412718 -4844 412954
rect -4608 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588532 412954
rect 588768 412718 588852 412954
rect 589088 412718 592960 412954
rect -9036 412634 592960 412718
rect -9036 412398 -5164 412634
rect -4928 412398 -4844 412634
rect -4608 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588532 412634
rect 588768 412398 588852 412634
rect 589088 412398 592960 412634
rect -9036 412366 592960 412398
rect -9036 408454 592960 408486
rect -9036 408218 -4204 408454
rect -3968 408218 -3884 408454
rect -3648 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587572 408454
rect 587808 408218 587892 408454
rect 588128 408218 592960 408454
rect -9036 408134 592960 408218
rect -9036 407898 -4204 408134
rect -3968 407898 -3884 408134
rect -3648 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587572 408134
rect 587808 407898 587892 408134
rect 588128 407898 592960 408134
rect -9036 407866 592960 407898
rect -9036 403954 592960 403986
rect -9036 403718 -3244 403954
rect -3008 403718 -2924 403954
rect -2688 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 252010 403954
rect 252246 403718 282730 403954
rect 282966 403718 313450 403954
rect 313686 403718 344170 403954
rect 344406 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586612 403954
rect 586848 403718 586932 403954
rect 587168 403718 592960 403954
rect -9036 403634 592960 403718
rect -9036 403398 -3244 403634
rect -3008 403398 -2924 403634
rect -2688 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 252010 403634
rect 252246 403398 282730 403634
rect 282966 403398 313450 403634
rect 313686 403398 344170 403634
rect 344406 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586612 403634
rect 586848 403398 586932 403634
rect 587168 403398 592960 403634
rect -9036 403366 592960 403398
rect -9036 399454 592960 399486
rect -9036 399218 -2284 399454
rect -2048 399218 -1964 399454
rect -1728 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 236650 399454
rect 236886 399218 267370 399454
rect 267606 399218 298090 399454
rect 298326 399218 328810 399454
rect 329046 399218 359530 399454
rect 359766 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585652 399454
rect 585888 399218 585972 399454
rect 586208 399218 592960 399454
rect -9036 399134 592960 399218
rect -9036 398898 -2284 399134
rect -2048 398898 -1964 399134
rect -1728 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 236650 399134
rect 236886 398898 267370 399134
rect 267606 398898 298090 399134
rect 298326 398898 328810 399134
rect 329046 398898 359530 399134
rect 359766 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585652 399134
rect 585888 398898 585972 399134
rect 586208 398898 592960 399134
rect -9036 398866 592960 398898
rect -9036 394954 592960 394986
rect -9036 394718 -9004 394954
rect -8768 394718 -8684 394954
rect -8448 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592372 394954
rect 592608 394718 592692 394954
rect 592928 394718 592960 394954
rect -9036 394634 592960 394718
rect -9036 394398 -9004 394634
rect -8768 394398 -8684 394634
rect -8448 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592372 394634
rect 592608 394398 592692 394634
rect 592928 394398 592960 394634
rect -9036 394366 592960 394398
rect -9036 390454 592960 390486
rect -9036 390218 -8044 390454
rect -7808 390218 -7724 390454
rect -7488 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591412 390454
rect 591648 390218 591732 390454
rect 591968 390218 592960 390454
rect -9036 390134 592960 390218
rect -9036 389898 -8044 390134
rect -7808 389898 -7724 390134
rect -7488 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591412 390134
rect 591648 389898 591732 390134
rect 591968 389898 592960 390134
rect -9036 389866 592960 389898
rect -9036 385954 592960 385986
rect -9036 385718 -7084 385954
rect -6848 385718 -6764 385954
rect -6528 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590452 385954
rect 590688 385718 590772 385954
rect 591008 385718 592960 385954
rect -9036 385634 592960 385718
rect -9036 385398 -7084 385634
rect -6848 385398 -6764 385634
rect -6528 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590452 385634
rect 590688 385398 590772 385634
rect 591008 385398 592960 385634
rect -9036 385366 592960 385398
rect -9036 381454 592960 381486
rect -9036 381218 -6124 381454
rect -5888 381218 -5804 381454
rect -5568 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589492 381454
rect 589728 381218 589812 381454
rect 590048 381218 592960 381454
rect -9036 381134 592960 381218
rect -9036 380898 -6124 381134
rect -5888 380898 -5804 381134
rect -5568 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589492 381134
rect 589728 380898 589812 381134
rect 590048 380898 592960 381134
rect -9036 380866 592960 380898
rect -9036 376954 592960 376986
rect -9036 376718 -5164 376954
rect -4928 376718 -4844 376954
rect -4608 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588532 376954
rect 588768 376718 588852 376954
rect 589088 376718 592960 376954
rect -9036 376634 592960 376718
rect -9036 376398 -5164 376634
rect -4928 376398 -4844 376634
rect -4608 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588532 376634
rect 588768 376398 588852 376634
rect 589088 376398 592960 376634
rect -9036 376366 592960 376398
rect -9036 372454 592960 372486
rect -9036 372218 -4204 372454
rect -3968 372218 -3884 372454
rect -3648 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587572 372454
rect 587808 372218 587892 372454
rect 588128 372218 592960 372454
rect -9036 372134 592960 372218
rect -9036 371898 -4204 372134
rect -3968 371898 -3884 372134
rect -3648 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587572 372134
rect 587808 371898 587892 372134
rect 588128 371898 592960 372134
rect -9036 371866 592960 371898
rect -9036 367954 592960 367986
rect -9036 367718 -3244 367954
rect -3008 367718 -2924 367954
rect -2688 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 119610 367954
rect 119846 367718 150330 367954
rect 150566 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 252010 367954
rect 252246 367718 282730 367954
rect 282966 367718 313450 367954
rect 313686 367718 344170 367954
rect 344406 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586612 367954
rect 586848 367718 586932 367954
rect 587168 367718 592960 367954
rect -9036 367634 592960 367718
rect -9036 367398 -3244 367634
rect -3008 367398 -2924 367634
rect -2688 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 119610 367634
rect 119846 367398 150330 367634
rect 150566 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 252010 367634
rect 252246 367398 282730 367634
rect 282966 367398 313450 367634
rect 313686 367398 344170 367634
rect 344406 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586612 367634
rect 586848 367398 586932 367634
rect 587168 367398 592960 367634
rect -9036 367366 592960 367398
rect -9036 363454 592960 363486
rect -9036 363218 -2284 363454
rect -2048 363218 -1964 363454
rect -1728 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 104250 363454
rect 104486 363218 134970 363454
rect 135206 363218 165690 363454
rect 165926 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 236650 363454
rect 236886 363218 267370 363454
rect 267606 363218 298090 363454
rect 298326 363218 328810 363454
rect 329046 363218 359530 363454
rect 359766 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585652 363454
rect 585888 363218 585972 363454
rect 586208 363218 592960 363454
rect -9036 363134 592960 363218
rect -9036 362898 -2284 363134
rect -2048 362898 -1964 363134
rect -1728 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 104250 363134
rect 104486 362898 134970 363134
rect 135206 362898 165690 363134
rect 165926 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 236650 363134
rect 236886 362898 267370 363134
rect 267606 362898 298090 363134
rect 298326 362898 328810 363134
rect 329046 362898 359530 363134
rect 359766 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585652 363134
rect 585888 362898 585972 363134
rect 586208 362898 592960 363134
rect -9036 362866 592960 362898
rect -9036 358954 592960 358986
rect -9036 358718 -9004 358954
rect -8768 358718 -8684 358954
rect -8448 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592372 358954
rect 592608 358718 592692 358954
rect 592928 358718 592960 358954
rect -9036 358634 592960 358718
rect -9036 358398 -9004 358634
rect -8768 358398 -8684 358634
rect -8448 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592372 358634
rect 592608 358398 592692 358634
rect 592928 358398 592960 358634
rect -9036 358366 592960 358398
rect -9036 354454 592960 354486
rect -9036 354218 -8044 354454
rect -7808 354218 -7724 354454
rect -7488 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591412 354454
rect 591648 354218 591732 354454
rect 591968 354218 592960 354454
rect -9036 354134 592960 354218
rect -9036 353898 -8044 354134
rect -7808 353898 -7724 354134
rect -7488 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591412 354134
rect 591648 353898 591732 354134
rect 591968 353898 592960 354134
rect -9036 353866 592960 353898
rect -9036 349954 592960 349986
rect -9036 349718 -7084 349954
rect -6848 349718 -6764 349954
rect -6528 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590452 349954
rect 590688 349718 590772 349954
rect 591008 349718 592960 349954
rect -9036 349634 592960 349718
rect -9036 349398 -7084 349634
rect -6848 349398 -6764 349634
rect -6528 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590452 349634
rect 590688 349398 590772 349634
rect 591008 349398 592960 349634
rect -9036 349366 592960 349398
rect -9036 345454 592960 345486
rect -9036 345218 -6124 345454
rect -5888 345218 -5804 345454
rect -5568 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589492 345454
rect 589728 345218 589812 345454
rect 590048 345218 592960 345454
rect -9036 345134 592960 345218
rect -9036 344898 -6124 345134
rect -5888 344898 -5804 345134
rect -5568 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589492 345134
rect 589728 344898 589812 345134
rect 590048 344898 592960 345134
rect -9036 344866 592960 344898
rect -9036 340954 592960 340986
rect -9036 340718 -5164 340954
rect -4928 340718 -4844 340954
rect -4608 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588532 340954
rect 588768 340718 588852 340954
rect 589088 340718 592960 340954
rect -9036 340634 592960 340718
rect -9036 340398 -5164 340634
rect -4928 340398 -4844 340634
rect -4608 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588532 340634
rect 588768 340398 588852 340634
rect 589088 340398 592960 340634
rect -9036 340366 592960 340398
rect -9036 336454 592960 336486
rect -9036 336218 -4204 336454
rect -3968 336218 -3884 336454
rect -3648 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587572 336454
rect 587808 336218 587892 336454
rect 588128 336218 592960 336454
rect -9036 336134 592960 336218
rect -9036 335898 -4204 336134
rect -3968 335898 -3884 336134
rect -3648 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587572 336134
rect 587808 335898 587892 336134
rect 588128 335898 592960 336134
rect -9036 335866 592960 335898
rect -9036 331954 592960 331986
rect -9036 331718 -3244 331954
rect -3008 331718 -2924 331954
rect -2688 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 119610 331954
rect 119846 331718 150330 331954
rect 150566 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 252010 331954
rect 252246 331718 282730 331954
rect 282966 331718 313450 331954
rect 313686 331718 344170 331954
rect 344406 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586612 331954
rect 586848 331718 586932 331954
rect 587168 331718 592960 331954
rect -9036 331634 592960 331718
rect -9036 331398 -3244 331634
rect -3008 331398 -2924 331634
rect -2688 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 119610 331634
rect 119846 331398 150330 331634
rect 150566 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 252010 331634
rect 252246 331398 282730 331634
rect 282966 331398 313450 331634
rect 313686 331398 344170 331634
rect 344406 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586612 331634
rect 586848 331398 586932 331634
rect 587168 331398 592960 331634
rect -9036 331366 592960 331398
rect -9036 327454 592960 327486
rect -9036 327218 -2284 327454
rect -2048 327218 -1964 327454
rect -1728 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 104250 327454
rect 104486 327218 134970 327454
rect 135206 327218 165690 327454
rect 165926 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 236650 327454
rect 236886 327218 267370 327454
rect 267606 327218 298090 327454
rect 298326 327218 328810 327454
rect 329046 327218 359530 327454
rect 359766 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585652 327454
rect 585888 327218 585972 327454
rect 586208 327218 592960 327454
rect -9036 327134 592960 327218
rect -9036 326898 -2284 327134
rect -2048 326898 -1964 327134
rect -1728 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 104250 327134
rect 104486 326898 134970 327134
rect 135206 326898 165690 327134
rect 165926 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 236650 327134
rect 236886 326898 267370 327134
rect 267606 326898 298090 327134
rect 298326 326898 328810 327134
rect 329046 326898 359530 327134
rect 359766 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585652 327134
rect 585888 326898 585972 327134
rect 586208 326898 592960 327134
rect -9036 326866 592960 326898
rect -9036 322954 592960 322986
rect -9036 322718 -9004 322954
rect -8768 322718 -8684 322954
rect -8448 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592372 322954
rect 592608 322718 592692 322954
rect 592928 322718 592960 322954
rect -9036 322634 592960 322718
rect -9036 322398 -9004 322634
rect -8768 322398 -8684 322634
rect -8448 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592372 322634
rect 592608 322398 592692 322634
rect 592928 322398 592960 322634
rect -9036 322366 592960 322398
rect -9036 318454 592960 318486
rect -9036 318218 -8044 318454
rect -7808 318218 -7724 318454
rect -7488 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591412 318454
rect 591648 318218 591732 318454
rect 591968 318218 592960 318454
rect -9036 318134 592960 318218
rect -9036 317898 -8044 318134
rect -7808 317898 -7724 318134
rect -7488 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591412 318134
rect 591648 317898 591732 318134
rect 591968 317898 592960 318134
rect -9036 317866 592960 317898
rect -9036 313954 592960 313986
rect -9036 313718 -7084 313954
rect -6848 313718 -6764 313954
rect -6528 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590452 313954
rect 590688 313718 590772 313954
rect 591008 313718 592960 313954
rect -9036 313634 592960 313718
rect -9036 313398 -7084 313634
rect -6848 313398 -6764 313634
rect -6528 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590452 313634
rect 590688 313398 590772 313634
rect 591008 313398 592960 313634
rect -9036 313366 592960 313398
rect -9036 309454 592960 309486
rect -9036 309218 -6124 309454
rect -5888 309218 -5804 309454
rect -5568 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589492 309454
rect 589728 309218 589812 309454
rect 590048 309218 592960 309454
rect -9036 309134 592960 309218
rect -9036 308898 -6124 309134
rect -5888 308898 -5804 309134
rect -5568 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589492 309134
rect 589728 308898 589812 309134
rect 590048 308898 592960 309134
rect -9036 308866 592960 308898
rect -9036 304954 592960 304986
rect -9036 304718 -5164 304954
rect -4928 304718 -4844 304954
rect -4608 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588532 304954
rect 588768 304718 588852 304954
rect 589088 304718 592960 304954
rect -9036 304634 592960 304718
rect -9036 304398 -5164 304634
rect -4928 304398 -4844 304634
rect -4608 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588532 304634
rect 588768 304398 588852 304634
rect 589088 304398 592960 304634
rect -9036 304366 592960 304398
rect -9036 300454 592960 300486
rect -9036 300218 -4204 300454
rect -3968 300218 -3884 300454
rect -3648 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587572 300454
rect 587808 300218 587892 300454
rect 588128 300218 592960 300454
rect -9036 300134 592960 300218
rect -9036 299898 -4204 300134
rect -3968 299898 -3884 300134
rect -3648 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587572 300134
rect 587808 299898 587892 300134
rect 588128 299898 592960 300134
rect -9036 299866 592960 299898
rect -9036 295954 592960 295986
rect -9036 295718 -3244 295954
rect -3008 295718 -2924 295954
rect -2688 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586612 295954
rect 586848 295718 586932 295954
rect 587168 295718 592960 295954
rect -9036 295634 592960 295718
rect -9036 295398 -3244 295634
rect -3008 295398 -2924 295634
rect -2688 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586612 295634
rect 586848 295398 586932 295634
rect 587168 295398 592960 295634
rect -9036 295366 592960 295398
rect -9036 291454 592960 291486
rect -9036 291218 -2284 291454
rect -2048 291218 -1964 291454
rect -1728 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585652 291454
rect 585888 291218 585972 291454
rect 586208 291218 592960 291454
rect -9036 291134 592960 291218
rect -9036 290898 -2284 291134
rect -2048 290898 -1964 291134
rect -1728 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585652 291134
rect 585888 290898 585972 291134
rect 586208 290898 592960 291134
rect -9036 290866 592960 290898
rect -9036 286954 592960 286986
rect -9036 286718 -9004 286954
rect -8768 286718 -8684 286954
rect -8448 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592372 286954
rect 592608 286718 592692 286954
rect 592928 286718 592960 286954
rect -9036 286634 592960 286718
rect -9036 286398 -9004 286634
rect -8768 286398 -8684 286634
rect -8448 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592372 286634
rect 592608 286398 592692 286634
rect 592928 286398 592960 286634
rect -9036 286366 592960 286398
rect -9036 282454 592960 282486
rect -9036 282218 -8044 282454
rect -7808 282218 -7724 282454
rect -7488 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591412 282454
rect 591648 282218 591732 282454
rect 591968 282218 592960 282454
rect -9036 282134 592960 282218
rect -9036 281898 -8044 282134
rect -7808 281898 -7724 282134
rect -7488 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591412 282134
rect 591648 281898 591732 282134
rect 591968 281898 592960 282134
rect -9036 281866 592960 281898
rect -9036 277954 592960 277986
rect -9036 277718 -7084 277954
rect -6848 277718 -6764 277954
rect -6528 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590452 277954
rect 590688 277718 590772 277954
rect 591008 277718 592960 277954
rect -9036 277634 592960 277718
rect -9036 277398 -7084 277634
rect -6848 277398 -6764 277634
rect -6528 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590452 277634
rect 590688 277398 590772 277634
rect 591008 277398 592960 277634
rect -9036 277366 592960 277398
rect -9036 273454 592960 273486
rect -9036 273218 -6124 273454
rect -5888 273218 -5804 273454
rect -5568 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589492 273454
rect 589728 273218 589812 273454
rect 590048 273218 592960 273454
rect -9036 273134 592960 273218
rect -9036 272898 -6124 273134
rect -5888 272898 -5804 273134
rect -5568 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589492 273134
rect 589728 272898 589812 273134
rect 590048 272898 592960 273134
rect -9036 272866 592960 272898
rect -9036 268954 592960 268986
rect -9036 268718 -5164 268954
rect -4928 268718 -4844 268954
rect -4608 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588532 268954
rect 588768 268718 588852 268954
rect 589088 268718 592960 268954
rect -9036 268634 592960 268718
rect -9036 268398 -5164 268634
rect -4928 268398 -4844 268634
rect -4608 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588532 268634
rect 588768 268398 588852 268634
rect 589088 268398 592960 268634
rect -9036 268366 592960 268398
rect -9036 264454 592960 264486
rect -9036 264218 -4204 264454
rect -3968 264218 -3884 264454
rect -3648 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587572 264454
rect 587808 264218 587892 264454
rect 588128 264218 592960 264454
rect -9036 264134 592960 264218
rect -9036 263898 -4204 264134
rect -3968 263898 -3884 264134
rect -3648 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587572 264134
rect 587808 263898 587892 264134
rect 588128 263898 592960 264134
rect -9036 263866 592960 263898
rect -9036 259954 592960 259986
rect -9036 259718 -3244 259954
rect -3008 259718 -2924 259954
rect -2688 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586612 259954
rect 586848 259718 586932 259954
rect 587168 259718 592960 259954
rect -9036 259634 592960 259718
rect -9036 259398 -3244 259634
rect -3008 259398 -2924 259634
rect -2688 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586612 259634
rect 586848 259398 586932 259634
rect 587168 259398 592960 259634
rect -9036 259366 592960 259398
rect -9036 255454 592960 255486
rect -9036 255218 -2284 255454
rect -2048 255218 -1964 255454
rect -1728 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585652 255454
rect 585888 255218 585972 255454
rect 586208 255218 592960 255454
rect -9036 255134 592960 255218
rect -9036 254898 -2284 255134
rect -2048 254898 -1964 255134
rect -1728 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585652 255134
rect 585888 254898 585972 255134
rect 586208 254898 592960 255134
rect -9036 254866 592960 254898
rect -9036 250954 592960 250986
rect -9036 250718 -9004 250954
rect -8768 250718 -8684 250954
rect -8448 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592372 250954
rect 592608 250718 592692 250954
rect 592928 250718 592960 250954
rect -9036 250634 592960 250718
rect -9036 250398 -9004 250634
rect -8768 250398 -8684 250634
rect -8448 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592372 250634
rect 592608 250398 592692 250634
rect 592928 250398 592960 250634
rect -9036 250366 592960 250398
rect -9036 246454 592960 246486
rect -9036 246218 -8044 246454
rect -7808 246218 -7724 246454
rect -7488 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591412 246454
rect 591648 246218 591732 246454
rect 591968 246218 592960 246454
rect -9036 246134 592960 246218
rect -9036 245898 -8044 246134
rect -7808 245898 -7724 246134
rect -7488 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591412 246134
rect 591648 245898 591732 246134
rect 591968 245898 592960 246134
rect -9036 245866 592960 245898
rect -9036 241954 592960 241986
rect -9036 241718 -7084 241954
rect -6848 241718 -6764 241954
rect -6528 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590452 241954
rect 590688 241718 590772 241954
rect 591008 241718 592960 241954
rect -9036 241634 592960 241718
rect -9036 241398 -7084 241634
rect -6848 241398 -6764 241634
rect -6528 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590452 241634
rect 590688 241398 590772 241634
rect 591008 241398 592960 241634
rect -9036 241366 592960 241398
rect -9036 237454 592960 237486
rect -9036 237218 -6124 237454
rect -5888 237218 -5804 237454
rect -5568 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589492 237454
rect 589728 237218 589812 237454
rect 590048 237218 592960 237454
rect -9036 237134 592960 237218
rect -9036 236898 -6124 237134
rect -5888 236898 -5804 237134
rect -5568 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589492 237134
rect 589728 236898 589812 237134
rect 590048 236898 592960 237134
rect -9036 236866 592960 236898
rect -9036 232954 592960 232986
rect -9036 232718 -5164 232954
rect -4928 232718 -4844 232954
rect -4608 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588532 232954
rect 588768 232718 588852 232954
rect 589088 232718 592960 232954
rect -9036 232634 592960 232718
rect -9036 232398 -5164 232634
rect -4928 232398 -4844 232634
rect -4608 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588532 232634
rect 588768 232398 588852 232634
rect 589088 232398 592960 232634
rect -9036 232366 592960 232398
rect -9036 228454 592960 228486
rect -9036 228218 -4204 228454
rect -3968 228218 -3884 228454
rect -3648 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587572 228454
rect 587808 228218 587892 228454
rect 588128 228218 592960 228454
rect -9036 228134 592960 228218
rect -9036 227898 -4204 228134
rect -3968 227898 -3884 228134
rect -3648 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587572 228134
rect 587808 227898 587892 228134
rect 588128 227898 592960 228134
rect -9036 227866 592960 227898
rect -9036 223954 592960 223986
rect -9036 223718 -3244 223954
rect -3008 223718 -2924 223954
rect -2688 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 220328 223954
rect 220564 223718 356056 223954
rect 356292 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586612 223954
rect 586848 223718 586932 223954
rect 587168 223718 592960 223954
rect -9036 223634 592960 223718
rect -9036 223398 -3244 223634
rect -3008 223398 -2924 223634
rect -2688 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 220328 223634
rect 220564 223398 356056 223634
rect 356292 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586612 223634
rect 586848 223398 586932 223634
rect 587168 223398 592960 223634
rect -9036 223366 592960 223398
rect -9036 219454 592960 219486
rect -9036 219218 -2284 219454
rect -2048 219218 -1964 219454
rect -1728 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 221008 219454
rect 221244 219218 355376 219454
rect 355612 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585652 219454
rect 585888 219218 585972 219454
rect 586208 219218 592960 219454
rect -9036 219134 592960 219218
rect -9036 218898 -2284 219134
rect -2048 218898 -1964 219134
rect -1728 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 221008 219134
rect 221244 218898 355376 219134
rect 355612 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585652 219134
rect 585888 218898 585972 219134
rect 586208 218898 592960 219134
rect -9036 218866 592960 218898
rect -9036 214954 592960 214986
rect -9036 214718 -9004 214954
rect -8768 214718 -8684 214954
rect -8448 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592372 214954
rect 592608 214718 592692 214954
rect 592928 214718 592960 214954
rect -9036 214634 592960 214718
rect -9036 214398 -9004 214634
rect -8768 214398 -8684 214634
rect -8448 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592372 214634
rect 592608 214398 592692 214634
rect 592928 214398 592960 214634
rect -9036 214366 592960 214398
rect -9036 210454 592960 210486
rect -9036 210218 -8044 210454
rect -7808 210218 -7724 210454
rect -7488 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591412 210454
rect 591648 210218 591732 210454
rect 591968 210218 592960 210454
rect -9036 210134 592960 210218
rect -9036 209898 -8044 210134
rect -7808 209898 -7724 210134
rect -7488 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591412 210134
rect 591648 209898 591732 210134
rect 591968 209898 592960 210134
rect -9036 209866 592960 209898
rect -9036 205954 592960 205986
rect -9036 205718 -7084 205954
rect -6848 205718 -6764 205954
rect -6528 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590452 205954
rect 590688 205718 590772 205954
rect 591008 205718 592960 205954
rect -9036 205634 592960 205718
rect -9036 205398 -7084 205634
rect -6848 205398 -6764 205634
rect -6528 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590452 205634
rect 590688 205398 590772 205634
rect 591008 205398 592960 205634
rect -9036 205366 592960 205398
rect -9036 201454 592960 201486
rect -9036 201218 -6124 201454
rect -5888 201218 -5804 201454
rect -5568 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589492 201454
rect 589728 201218 589812 201454
rect 590048 201218 592960 201454
rect -9036 201134 592960 201218
rect -9036 200898 -6124 201134
rect -5888 200898 -5804 201134
rect -5568 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589492 201134
rect 589728 200898 589812 201134
rect 590048 200898 592960 201134
rect -9036 200866 592960 200898
rect -9036 196954 592960 196986
rect -9036 196718 -5164 196954
rect -4928 196718 -4844 196954
rect -4608 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588532 196954
rect 588768 196718 588852 196954
rect 589088 196718 592960 196954
rect -9036 196634 592960 196718
rect -9036 196398 -5164 196634
rect -4928 196398 -4844 196634
rect -4608 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588532 196634
rect 588768 196398 588852 196634
rect 589088 196398 592960 196634
rect -9036 196366 592960 196398
rect -9036 192454 592960 192486
rect -9036 192218 -4204 192454
rect -3968 192218 -3884 192454
rect -3648 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587572 192454
rect 587808 192218 587892 192454
rect 588128 192218 592960 192454
rect -9036 192134 592960 192218
rect -9036 191898 -4204 192134
rect -3968 191898 -3884 192134
rect -3648 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587572 192134
rect 587808 191898 587892 192134
rect 588128 191898 592960 192134
rect -9036 191866 592960 191898
rect -9036 187954 592960 187986
rect -9036 187718 -3244 187954
rect -3008 187718 -2924 187954
rect -2688 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 220328 187954
rect 220564 187718 356056 187954
rect 356292 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586612 187954
rect 586848 187718 586932 187954
rect 587168 187718 592960 187954
rect -9036 187634 592960 187718
rect -9036 187398 -3244 187634
rect -3008 187398 -2924 187634
rect -2688 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 220328 187634
rect 220564 187398 356056 187634
rect 356292 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586612 187634
rect 586848 187398 586932 187634
rect 587168 187398 592960 187634
rect -9036 187366 592960 187398
rect -9036 183454 592960 183486
rect -9036 183218 -2284 183454
rect -2048 183218 -1964 183454
rect -1728 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 221008 183454
rect 221244 183218 355376 183454
rect 355612 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585652 183454
rect 585888 183218 585972 183454
rect 586208 183218 592960 183454
rect -9036 183134 592960 183218
rect -9036 182898 -2284 183134
rect -2048 182898 -1964 183134
rect -1728 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 221008 183134
rect 221244 182898 355376 183134
rect 355612 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585652 183134
rect 585888 182898 585972 183134
rect 586208 182898 592960 183134
rect -9036 182866 592960 182898
rect -9036 178954 592960 178986
rect -9036 178718 -9004 178954
rect -8768 178718 -8684 178954
rect -8448 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592372 178954
rect 592608 178718 592692 178954
rect 592928 178718 592960 178954
rect -9036 178634 592960 178718
rect -9036 178398 -9004 178634
rect -8768 178398 -8684 178634
rect -8448 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592372 178634
rect 592608 178398 592692 178634
rect 592928 178398 592960 178634
rect -9036 178366 592960 178398
rect -9036 174454 592960 174486
rect -9036 174218 -8044 174454
rect -7808 174218 -7724 174454
rect -7488 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591412 174454
rect 591648 174218 591732 174454
rect 591968 174218 592960 174454
rect -9036 174134 592960 174218
rect -9036 173898 -8044 174134
rect -7808 173898 -7724 174134
rect -7488 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591412 174134
rect 591648 173898 591732 174134
rect 591968 173898 592960 174134
rect -9036 173866 592960 173898
rect -9036 169954 592960 169986
rect -9036 169718 -7084 169954
rect -6848 169718 -6764 169954
rect -6528 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590452 169954
rect 590688 169718 590772 169954
rect 591008 169718 592960 169954
rect -9036 169634 592960 169718
rect -9036 169398 -7084 169634
rect -6848 169398 -6764 169634
rect -6528 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590452 169634
rect 590688 169398 590772 169634
rect 591008 169398 592960 169634
rect -9036 169366 592960 169398
rect -9036 165454 592960 165486
rect -9036 165218 -6124 165454
rect -5888 165218 -5804 165454
rect -5568 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589492 165454
rect 589728 165218 589812 165454
rect 590048 165218 592960 165454
rect -9036 165134 592960 165218
rect -9036 164898 -6124 165134
rect -5888 164898 -5804 165134
rect -5568 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589492 165134
rect 589728 164898 589812 165134
rect 590048 164898 592960 165134
rect -9036 164866 592960 164898
rect -9036 160954 592960 160986
rect -9036 160718 -5164 160954
rect -4928 160718 -4844 160954
rect -4608 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588532 160954
rect 588768 160718 588852 160954
rect 589088 160718 592960 160954
rect -9036 160634 592960 160718
rect -9036 160398 -5164 160634
rect -4928 160398 -4844 160634
rect -4608 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588532 160634
rect 588768 160398 588852 160634
rect 589088 160398 592960 160634
rect -9036 160366 592960 160398
rect -9036 156454 592960 156486
rect -9036 156218 -4204 156454
rect -3968 156218 -3884 156454
rect -3648 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587572 156454
rect 587808 156218 587892 156454
rect 588128 156218 592960 156454
rect -9036 156134 592960 156218
rect -9036 155898 -4204 156134
rect -3968 155898 -3884 156134
rect -3648 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587572 156134
rect 587808 155898 587892 156134
rect 588128 155898 592960 156134
rect -9036 155866 592960 155898
rect -9036 151954 592960 151986
rect -9036 151718 -3244 151954
rect -3008 151718 -2924 151954
rect -2688 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586612 151954
rect 586848 151718 586932 151954
rect 587168 151718 592960 151954
rect -9036 151634 592960 151718
rect -9036 151398 -3244 151634
rect -3008 151398 -2924 151634
rect -2688 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586612 151634
rect 586848 151398 586932 151634
rect 587168 151398 592960 151634
rect -9036 151366 592960 151398
rect -9036 147454 592960 147486
rect -9036 147218 -2284 147454
rect -2048 147218 -1964 147454
rect -1728 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585652 147454
rect 585888 147218 585972 147454
rect 586208 147218 592960 147454
rect -9036 147134 592960 147218
rect -9036 146898 -2284 147134
rect -2048 146898 -1964 147134
rect -1728 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585652 147134
rect 585888 146898 585972 147134
rect 586208 146898 592960 147134
rect -9036 146866 592960 146898
rect -9036 142954 592960 142986
rect -9036 142718 -9004 142954
rect -8768 142718 -8684 142954
rect -8448 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592372 142954
rect 592608 142718 592692 142954
rect 592928 142718 592960 142954
rect -9036 142634 592960 142718
rect -9036 142398 -9004 142634
rect -8768 142398 -8684 142634
rect -8448 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592372 142634
rect 592608 142398 592692 142634
rect 592928 142398 592960 142634
rect -9036 142366 592960 142398
rect -9036 138454 592960 138486
rect -9036 138218 -8044 138454
rect -7808 138218 -7724 138454
rect -7488 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591412 138454
rect 591648 138218 591732 138454
rect 591968 138218 592960 138454
rect -9036 138134 592960 138218
rect -9036 137898 -8044 138134
rect -7808 137898 -7724 138134
rect -7488 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591412 138134
rect 591648 137898 591732 138134
rect 591968 137898 592960 138134
rect -9036 137866 592960 137898
rect -9036 133954 592960 133986
rect -9036 133718 -7084 133954
rect -6848 133718 -6764 133954
rect -6528 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590452 133954
rect 590688 133718 590772 133954
rect 591008 133718 592960 133954
rect -9036 133634 592960 133718
rect -9036 133398 -7084 133634
rect -6848 133398 -6764 133634
rect -6528 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590452 133634
rect 590688 133398 590772 133634
rect 591008 133398 592960 133634
rect -9036 133366 592960 133398
rect -9036 129454 592960 129486
rect -9036 129218 -6124 129454
rect -5888 129218 -5804 129454
rect -5568 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589492 129454
rect 589728 129218 589812 129454
rect 590048 129218 592960 129454
rect -9036 129134 592960 129218
rect -9036 128898 -6124 129134
rect -5888 128898 -5804 129134
rect -5568 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589492 129134
rect 589728 128898 589812 129134
rect 590048 128898 592960 129134
rect -9036 128866 592960 128898
rect -9036 124954 592960 124986
rect -9036 124718 -5164 124954
rect -4928 124718 -4844 124954
rect -4608 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 123326 124954
rect 123562 124718 123646 124954
rect 123882 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588532 124954
rect 588768 124718 588852 124954
rect 589088 124718 592960 124954
rect -9036 124634 592960 124718
rect -9036 124398 -5164 124634
rect -4928 124398 -4844 124634
rect -4608 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 123326 124634
rect 123562 124398 123646 124634
rect 123882 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588532 124634
rect 588768 124398 588852 124634
rect 589088 124398 592960 124634
rect -9036 124366 592960 124398
rect -9036 120454 592960 120486
rect -9036 120218 -4204 120454
rect -3968 120218 -3884 120454
rect -3648 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587572 120454
rect 587808 120218 587892 120454
rect 588128 120218 592960 120454
rect -9036 120134 592960 120218
rect -9036 119898 -4204 120134
rect -3968 119898 -3884 120134
rect -3648 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587572 120134
rect 587808 119898 587892 120134
rect 588128 119898 592960 120134
rect -9036 119866 592960 119898
rect -9036 115954 592960 115986
rect -9036 115718 -3244 115954
rect -3008 115718 -2924 115954
rect -2688 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586612 115954
rect 586848 115718 586932 115954
rect 587168 115718 592960 115954
rect -9036 115634 592960 115718
rect -9036 115398 -3244 115634
rect -3008 115398 -2924 115634
rect -2688 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586612 115634
rect 586848 115398 586932 115634
rect 587168 115398 592960 115634
rect -9036 115366 592960 115398
rect -9036 111454 592960 111486
rect -9036 111218 -2284 111454
rect -2048 111218 -1964 111454
rect -1728 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585652 111454
rect 585888 111218 585972 111454
rect 586208 111218 592960 111454
rect -9036 111134 592960 111218
rect -9036 110898 -2284 111134
rect -2048 110898 -1964 111134
rect -1728 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585652 111134
rect 585888 110898 585972 111134
rect 586208 110898 592960 111134
rect -9036 110866 592960 110898
rect -9036 106954 592960 106986
rect -9036 106718 -9004 106954
rect -8768 106718 -8684 106954
rect -8448 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592372 106954
rect 592608 106718 592692 106954
rect 592928 106718 592960 106954
rect -9036 106634 592960 106718
rect -9036 106398 -9004 106634
rect -8768 106398 -8684 106634
rect -8448 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592372 106634
rect 592608 106398 592692 106634
rect 592928 106398 592960 106634
rect -9036 106366 592960 106398
rect -9036 102454 592960 102486
rect -9036 102218 -8044 102454
rect -7808 102218 -7724 102454
rect -7488 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591412 102454
rect 591648 102218 591732 102454
rect 591968 102218 592960 102454
rect -9036 102134 592960 102218
rect -9036 101898 -8044 102134
rect -7808 101898 -7724 102134
rect -7488 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591412 102134
rect 591648 101898 591732 102134
rect 591968 101898 592960 102134
rect -9036 101866 592960 101898
rect -9036 97954 592960 97986
rect -9036 97718 -7084 97954
rect -6848 97718 -6764 97954
rect -6528 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590452 97954
rect 590688 97718 590772 97954
rect 591008 97718 592960 97954
rect -9036 97634 592960 97718
rect -9036 97398 -7084 97634
rect -6848 97398 -6764 97634
rect -6528 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590452 97634
rect 590688 97398 590772 97634
rect 591008 97398 592960 97634
rect -9036 97366 592960 97398
rect -9036 93454 592960 93486
rect -9036 93218 -6124 93454
rect -5888 93218 -5804 93454
rect -5568 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589492 93454
rect 589728 93218 589812 93454
rect 590048 93218 592960 93454
rect -9036 93134 592960 93218
rect -9036 92898 -6124 93134
rect -5888 92898 -5804 93134
rect -5568 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589492 93134
rect 589728 92898 589812 93134
rect 590048 92898 592960 93134
rect -9036 92866 592960 92898
rect -9036 88954 592960 88986
rect -9036 88718 -5164 88954
rect -4928 88718 -4844 88954
rect -4608 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588532 88954
rect 588768 88718 588852 88954
rect 589088 88718 592960 88954
rect -9036 88634 592960 88718
rect -9036 88398 -5164 88634
rect -4928 88398 -4844 88634
rect -4608 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588532 88634
rect 588768 88398 588852 88634
rect 589088 88398 592960 88634
rect -9036 88366 592960 88398
rect -9036 84454 592960 84486
rect -9036 84218 -4204 84454
rect -3968 84218 -3884 84454
rect -3648 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587572 84454
rect 587808 84218 587892 84454
rect 588128 84218 592960 84454
rect -9036 84134 592960 84218
rect -9036 83898 -4204 84134
rect -3968 83898 -3884 84134
rect -3648 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587572 84134
rect 587808 83898 587892 84134
rect 588128 83898 592960 84134
rect -9036 83866 592960 83898
rect -9036 79954 592960 79986
rect -9036 79718 -3244 79954
rect -3008 79718 -2924 79954
rect -2688 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586612 79954
rect 586848 79718 586932 79954
rect 587168 79718 592960 79954
rect -9036 79634 592960 79718
rect -9036 79398 -3244 79634
rect -3008 79398 -2924 79634
rect -2688 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586612 79634
rect 586848 79398 586932 79634
rect 587168 79398 592960 79634
rect -9036 79366 592960 79398
rect -9036 75454 592960 75486
rect -9036 75218 -2284 75454
rect -2048 75218 -1964 75454
rect -1728 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585652 75454
rect 585888 75218 585972 75454
rect 586208 75218 592960 75454
rect -9036 75134 592960 75218
rect -9036 74898 -2284 75134
rect -2048 74898 -1964 75134
rect -1728 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585652 75134
rect 585888 74898 585972 75134
rect 586208 74898 592960 75134
rect -9036 74866 592960 74898
rect -9036 70954 592960 70986
rect -9036 70718 -9004 70954
rect -8768 70718 -8684 70954
rect -8448 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592372 70954
rect 592608 70718 592692 70954
rect 592928 70718 592960 70954
rect -9036 70634 592960 70718
rect -9036 70398 -9004 70634
rect -8768 70398 -8684 70634
rect -8448 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592372 70634
rect 592608 70398 592692 70634
rect 592928 70398 592960 70634
rect -9036 70366 592960 70398
rect -9036 66454 592960 66486
rect -9036 66218 -8044 66454
rect -7808 66218 -7724 66454
rect -7488 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591412 66454
rect 591648 66218 591732 66454
rect 591968 66218 592960 66454
rect -9036 66134 592960 66218
rect -9036 65898 -8044 66134
rect -7808 65898 -7724 66134
rect -7488 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591412 66134
rect 591648 65898 591732 66134
rect 591968 65898 592960 66134
rect -9036 65866 592960 65898
rect -9036 61954 592960 61986
rect -9036 61718 -7084 61954
rect -6848 61718 -6764 61954
rect -6528 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590452 61954
rect 590688 61718 590772 61954
rect 591008 61718 592960 61954
rect -9036 61634 592960 61718
rect -9036 61398 -7084 61634
rect -6848 61398 -6764 61634
rect -6528 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590452 61634
rect 590688 61398 590772 61634
rect 591008 61398 592960 61634
rect -9036 61366 592960 61398
rect -9036 57454 592960 57486
rect -9036 57218 -6124 57454
rect -5888 57218 -5804 57454
rect -5568 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589492 57454
rect 589728 57218 589812 57454
rect 590048 57218 592960 57454
rect -9036 57134 592960 57218
rect -9036 56898 -6124 57134
rect -5888 56898 -5804 57134
rect -5568 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589492 57134
rect 589728 56898 589812 57134
rect 590048 56898 592960 57134
rect -9036 56866 592960 56898
rect -9036 52954 592960 52986
rect -9036 52718 -5164 52954
rect -4928 52718 -4844 52954
rect -4608 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588532 52954
rect 588768 52718 588852 52954
rect 589088 52718 592960 52954
rect -9036 52634 592960 52718
rect -9036 52398 -5164 52634
rect -4928 52398 -4844 52634
rect -4608 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588532 52634
rect 588768 52398 588852 52634
rect 589088 52398 592960 52634
rect -9036 52366 592960 52398
rect -9036 48454 592960 48486
rect -9036 48218 -4204 48454
rect -3968 48218 -3884 48454
rect -3648 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587572 48454
rect 587808 48218 587892 48454
rect 588128 48218 592960 48454
rect -9036 48134 592960 48218
rect -9036 47898 -4204 48134
rect -3968 47898 -3884 48134
rect -3648 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587572 48134
rect 587808 47898 587892 48134
rect 588128 47898 592960 48134
rect -9036 47866 592960 47898
rect -9036 43954 592960 43986
rect -9036 43718 -3244 43954
rect -3008 43718 -2924 43954
rect -2688 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586612 43954
rect 586848 43718 586932 43954
rect 587168 43718 592960 43954
rect -9036 43634 592960 43718
rect -9036 43398 -3244 43634
rect -3008 43398 -2924 43634
rect -2688 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586612 43634
rect 586848 43398 586932 43634
rect 587168 43398 592960 43634
rect -9036 43366 592960 43398
rect -9036 39454 592960 39486
rect -9036 39218 -2284 39454
rect -2048 39218 -1964 39454
rect -1728 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585652 39454
rect 585888 39218 585972 39454
rect 586208 39218 592960 39454
rect -9036 39134 592960 39218
rect -9036 38898 -2284 39134
rect -2048 38898 -1964 39134
rect -1728 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585652 39134
rect 585888 38898 585972 39134
rect 586208 38898 592960 39134
rect -9036 38866 592960 38898
rect -9036 34954 592960 34986
rect -9036 34718 -9004 34954
rect -8768 34718 -8684 34954
rect -8448 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592372 34954
rect 592608 34718 592692 34954
rect 592928 34718 592960 34954
rect -9036 34634 592960 34718
rect -9036 34398 -9004 34634
rect -8768 34398 -8684 34634
rect -8448 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592372 34634
rect 592608 34398 592692 34634
rect 592928 34398 592960 34634
rect -9036 34366 592960 34398
rect -9036 30454 592960 30486
rect -9036 30218 -8044 30454
rect -7808 30218 -7724 30454
rect -7488 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591412 30454
rect 591648 30218 591732 30454
rect 591968 30218 592960 30454
rect -9036 30134 592960 30218
rect -9036 29898 -8044 30134
rect -7808 29898 -7724 30134
rect -7488 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591412 30134
rect 591648 29898 591732 30134
rect 591968 29898 592960 30134
rect -9036 29866 592960 29898
rect -9036 25954 592960 25986
rect -9036 25718 -7084 25954
rect -6848 25718 -6764 25954
rect -6528 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590452 25954
rect 590688 25718 590772 25954
rect 591008 25718 592960 25954
rect -9036 25634 592960 25718
rect -9036 25398 -7084 25634
rect -6848 25398 -6764 25634
rect -6528 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590452 25634
rect 590688 25398 590772 25634
rect 591008 25398 592960 25634
rect -9036 25366 592960 25398
rect -9036 21454 592960 21486
rect -9036 21218 -6124 21454
rect -5888 21218 -5804 21454
rect -5568 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589492 21454
rect 589728 21218 589812 21454
rect 590048 21218 592960 21454
rect -9036 21134 592960 21218
rect -9036 20898 -6124 21134
rect -5888 20898 -5804 21134
rect -5568 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589492 21134
rect 589728 20898 589812 21134
rect 590048 20898 592960 21134
rect -9036 20866 592960 20898
rect -9036 16954 592960 16986
rect -9036 16718 -5164 16954
rect -4928 16718 -4844 16954
rect -4608 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588532 16954
rect 588768 16718 588852 16954
rect 589088 16718 592960 16954
rect -9036 16634 592960 16718
rect -9036 16398 -5164 16634
rect -4928 16398 -4844 16634
rect -4608 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588532 16634
rect 588768 16398 588852 16634
rect 589088 16398 592960 16634
rect -9036 16366 592960 16398
rect -9036 12454 592960 12486
rect -9036 12218 -4204 12454
rect -3968 12218 -3884 12454
rect -3648 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587572 12454
rect 587808 12218 587892 12454
rect 588128 12218 592960 12454
rect -9036 12134 592960 12218
rect -9036 11898 -4204 12134
rect -3968 11898 -3884 12134
rect -3648 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587572 12134
rect 587808 11898 587892 12134
rect 588128 11898 592960 12134
rect -9036 11866 592960 11898
rect -9036 7954 592960 7986
rect -9036 7718 -3244 7954
rect -3008 7718 -2924 7954
rect -2688 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586612 7954
rect 586848 7718 586932 7954
rect 587168 7718 592960 7954
rect -9036 7634 592960 7718
rect -9036 7398 -3244 7634
rect -3008 7398 -2924 7634
rect -2688 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586612 7634
rect 586848 7398 586932 7634
rect 587168 7398 592960 7634
rect -9036 7366 592960 7398
rect -9036 3454 592960 3486
rect -9036 3218 -2284 3454
rect -2048 3218 -1964 3454
rect -1728 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585652 3454
rect 585888 3218 585972 3454
rect 586208 3218 592960 3454
rect -9036 3134 592960 3218
rect -9036 2898 -2284 3134
rect -2048 2898 -1964 3134
rect -1728 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585652 3134
rect 585888 2898 585972 3134
rect 586208 2898 592960 3134
rect -9036 2866 592960 2898
rect -2316 -656 586240 -624
rect -2316 -892 -2284 -656
rect -2048 -892 -1964 -656
rect -1728 -892 1826 -656
rect 2062 -892 2146 -656
rect 2382 -892 37826 -656
rect 38062 -892 38146 -656
rect 38382 -892 73826 -656
rect 74062 -892 74146 -656
rect 74382 -892 109826 -656
rect 110062 -892 110146 -656
rect 110382 -892 145826 -656
rect 146062 -892 146146 -656
rect 146382 -892 181826 -656
rect 182062 -892 182146 -656
rect 182382 -892 217826 -656
rect 218062 -892 218146 -656
rect 218382 -892 253826 -656
rect 254062 -892 254146 -656
rect 254382 -892 289826 -656
rect 290062 -892 290146 -656
rect 290382 -892 325826 -656
rect 326062 -892 326146 -656
rect 326382 -892 361826 -656
rect 362062 -892 362146 -656
rect 362382 -892 397826 -656
rect 398062 -892 398146 -656
rect 398382 -892 433826 -656
rect 434062 -892 434146 -656
rect 434382 -892 469826 -656
rect 470062 -892 470146 -656
rect 470382 -892 505826 -656
rect 506062 -892 506146 -656
rect 506382 -892 541826 -656
rect 542062 -892 542146 -656
rect 542382 -892 577826 -656
rect 578062 -892 578146 -656
rect 578382 -892 585652 -656
rect 585888 -892 585972 -656
rect 586208 -892 586240 -656
rect -2316 -976 586240 -892
rect -2316 -1212 -2284 -976
rect -2048 -1212 -1964 -976
rect -1728 -1212 1826 -976
rect 2062 -1212 2146 -976
rect 2382 -1212 37826 -976
rect 38062 -1212 38146 -976
rect 38382 -1212 73826 -976
rect 74062 -1212 74146 -976
rect 74382 -1212 109826 -976
rect 110062 -1212 110146 -976
rect 110382 -1212 145826 -976
rect 146062 -1212 146146 -976
rect 146382 -1212 181826 -976
rect 182062 -1212 182146 -976
rect 182382 -1212 217826 -976
rect 218062 -1212 218146 -976
rect 218382 -1212 253826 -976
rect 254062 -1212 254146 -976
rect 254382 -1212 289826 -976
rect 290062 -1212 290146 -976
rect 290382 -1212 325826 -976
rect 326062 -1212 326146 -976
rect 326382 -1212 361826 -976
rect 362062 -1212 362146 -976
rect 362382 -1212 397826 -976
rect 398062 -1212 398146 -976
rect 398382 -1212 433826 -976
rect 434062 -1212 434146 -976
rect 434382 -1212 469826 -976
rect 470062 -1212 470146 -976
rect 470382 -1212 505826 -976
rect 506062 -1212 506146 -976
rect 506382 -1212 541826 -976
rect 542062 -1212 542146 -976
rect 542382 -1212 577826 -976
rect 578062 -1212 578146 -976
rect 578382 -1212 585652 -976
rect 585888 -1212 585972 -976
rect 586208 -1212 586240 -976
rect -2316 -1244 586240 -1212
rect -3276 -1616 587200 -1584
rect -3276 -1852 -3244 -1616
rect -3008 -1852 -2924 -1616
rect -2688 -1852 6326 -1616
rect 6562 -1852 6646 -1616
rect 6882 -1852 42326 -1616
rect 42562 -1852 42646 -1616
rect 42882 -1852 78326 -1616
rect 78562 -1852 78646 -1616
rect 78882 -1852 114326 -1616
rect 114562 -1852 114646 -1616
rect 114882 -1852 150326 -1616
rect 150562 -1852 150646 -1616
rect 150882 -1852 186326 -1616
rect 186562 -1852 186646 -1616
rect 186882 -1852 222326 -1616
rect 222562 -1852 222646 -1616
rect 222882 -1852 258326 -1616
rect 258562 -1852 258646 -1616
rect 258882 -1852 294326 -1616
rect 294562 -1852 294646 -1616
rect 294882 -1852 330326 -1616
rect 330562 -1852 330646 -1616
rect 330882 -1852 366326 -1616
rect 366562 -1852 366646 -1616
rect 366882 -1852 402326 -1616
rect 402562 -1852 402646 -1616
rect 402882 -1852 438326 -1616
rect 438562 -1852 438646 -1616
rect 438882 -1852 474326 -1616
rect 474562 -1852 474646 -1616
rect 474882 -1852 510326 -1616
rect 510562 -1852 510646 -1616
rect 510882 -1852 546326 -1616
rect 546562 -1852 546646 -1616
rect 546882 -1852 582326 -1616
rect 582562 -1852 582646 -1616
rect 582882 -1852 586612 -1616
rect 586848 -1852 586932 -1616
rect 587168 -1852 587200 -1616
rect -3276 -1936 587200 -1852
rect -3276 -2172 -3244 -1936
rect -3008 -2172 -2924 -1936
rect -2688 -2172 6326 -1936
rect 6562 -2172 6646 -1936
rect 6882 -2172 42326 -1936
rect 42562 -2172 42646 -1936
rect 42882 -2172 78326 -1936
rect 78562 -2172 78646 -1936
rect 78882 -2172 114326 -1936
rect 114562 -2172 114646 -1936
rect 114882 -2172 150326 -1936
rect 150562 -2172 150646 -1936
rect 150882 -2172 186326 -1936
rect 186562 -2172 186646 -1936
rect 186882 -2172 222326 -1936
rect 222562 -2172 222646 -1936
rect 222882 -2172 258326 -1936
rect 258562 -2172 258646 -1936
rect 258882 -2172 294326 -1936
rect 294562 -2172 294646 -1936
rect 294882 -2172 330326 -1936
rect 330562 -2172 330646 -1936
rect 330882 -2172 366326 -1936
rect 366562 -2172 366646 -1936
rect 366882 -2172 402326 -1936
rect 402562 -2172 402646 -1936
rect 402882 -2172 438326 -1936
rect 438562 -2172 438646 -1936
rect 438882 -2172 474326 -1936
rect 474562 -2172 474646 -1936
rect 474882 -2172 510326 -1936
rect 510562 -2172 510646 -1936
rect 510882 -2172 546326 -1936
rect 546562 -2172 546646 -1936
rect 546882 -2172 582326 -1936
rect 582562 -2172 582646 -1936
rect 582882 -2172 586612 -1936
rect 586848 -2172 586932 -1936
rect 587168 -2172 587200 -1936
rect -3276 -2204 587200 -2172
rect -4236 -2576 588160 -2544
rect -4236 -2812 -4204 -2576
rect -3968 -2812 -3884 -2576
rect -3648 -2812 10826 -2576
rect 11062 -2812 11146 -2576
rect 11382 -2812 46826 -2576
rect 47062 -2812 47146 -2576
rect 47382 -2812 82826 -2576
rect 83062 -2812 83146 -2576
rect 83382 -2812 118826 -2576
rect 119062 -2812 119146 -2576
rect 119382 -2812 154826 -2576
rect 155062 -2812 155146 -2576
rect 155382 -2812 190826 -2576
rect 191062 -2812 191146 -2576
rect 191382 -2812 226826 -2576
rect 227062 -2812 227146 -2576
rect 227382 -2812 262826 -2576
rect 263062 -2812 263146 -2576
rect 263382 -2812 298826 -2576
rect 299062 -2812 299146 -2576
rect 299382 -2812 334826 -2576
rect 335062 -2812 335146 -2576
rect 335382 -2812 370826 -2576
rect 371062 -2812 371146 -2576
rect 371382 -2812 406826 -2576
rect 407062 -2812 407146 -2576
rect 407382 -2812 442826 -2576
rect 443062 -2812 443146 -2576
rect 443382 -2812 478826 -2576
rect 479062 -2812 479146 -2576
rect 479382 -2812 514826 -2576
rect 515062 -2812 515146 -2576
rect 515382 -2812 550826 -2576
rect 551062 -2812 551146 -2576
rect 551382 -2812 587572 -2576
rect 587808 -2812 587892 -2576
rect 588128 -2812 588160 -2576
rect -4236 -2896 588160 -2812
rect -4236 -3132 -4204 -2896
rect -3968 -3132 -3884 -2896
rect -3648 -3132 10826 -2896
rect 11062 -3132 11146 -2896
rect 11382 -3132 46826 -2896
rect 47062 -3132 47146 -2896
rect 47382 -3132 82826 -2896
rect 83062 -3132 83146 -2896
rect 83382 -3132 118826 -2896
rect 119062 -3132 119146 -2896
rect 119382 -3132 154826 -2896
rect 155062 -3132 155146 -2896
rect 155382 -3132 190826 -2896
rect 191062 -3132 191146 -2896
rect 191382 -3132 226826 -2896
rect 227062 -3132 227146 -2896
rect 227382 -3132 262826 -2896
rect 263062 -3132 263146 -2896
rect 263382 -3132 298826 -2896
rect 299062 -3132 299146 -2896
rect 299382 -3132 334826 -2896
rect 335062 -3132 335146 -2896
rect 335382 -3132 370826 -2896
rect 371062 -3132 371146 -2896
rect 371382 -3132 406826 -2896
rect 407062 -3132 407146 -2896
rect 407382 -3132 442826 -2896
rect 443062 -3132 443146 -2896
rect 443382 -3132 478826 -2896
rect 479062 -3132 479146 -2896
rect 479382 -3132 514826 -2896
rect 515062 -3132 515146 -2896
rect 515382 -3132 550826 -2896
rect 551062 -3132 551146 -2896
rect 551382 -3132 587572 -2896
rect 587808 -3132 587892 -2896
rect 588128 -3132 588160 -2896
rect -4236 -3164 588160 -3132
rect -5196 -3536 589120 -3504
rect -5196 -3772 -5164 -3536
rect -4928 -3772 -4844 -3536
rect -4608 -3772 15326 -3536
rect 15562 -3772 15646 -3536
rect 15882 -3772 51326 -3536
rect 51562 -3772 51646 -3536
rect 51882 -3772 87326 -3536
rect 87562 -3772 87646 -3536
rect 87882 -3772 123326 -3536
rect 123562 -3772 123646 -3536
rect 123882 -3772 159326 -3536
rect 159562 -3772 159646 -3536
rect 159882 -3772 195326 -3536
rect 195562 -3772 195646 -3536
rect 195882 -3772 231326 -3536
rect 231562 -3772 231646 -3536
rect 231882 -3772 267326 -3536
rect 267562 -3772 267646 -3536
rect 267882 -3772 303326 -3536
rect 303562 -3772 303646 -3536
rect 303882 -3772 339326 -3536
rect 339562 -3772 339646 -3536
rect 339882 -3772 375326 -3536
rect 375562 -3772 375646 -3536
rect 375882 -3772 411326 -3536
rect 411562 -3772 411646 -3536
rect 411882 -3772 447326 -3536
rect 447562 -3772 447646 -3536
rect 447882 -3772 483326 -3536
rect 483562 -3772 483646 -3536
rect 483882 -3772 519326 -3536
rect 519562 -3772 519646 -3536
rect 519882 -3772 555326 -3536
rect 555562 -3772 555646 -3536
rect 555882 -3772 588532 -3536
rect 588768 -3772 588852 -3536
rect 589088 -3772 589120 -3536
rect -5196 -3856 589120 -3772
rect -5196 -4092 -5164 -3856
rect -4928 -4092 -4844 -3856
rect -4608 -4092 15326 -3856
rect 15562 -4092 15646 -3856
rect 15882 -4092 51326 -3856
rect 51562 -4092 51646 -3856
rect 51882 -4092 87326 -3856
rect 87562 -4092 87646 -3856
rect 87882 -4092 123326 -3856
rect 123562 -4092 123646 -3856
rect 123882 -4092 159326 -3856
rect 159562 -4092 159646 -3856
rect 159882 -4092 195326 -3856
rect 195562 -4092 195646 -3856
rect 195882 -4092 231326 -3856
rect 231562 -4092 231646 -3856
rect 231882 -4092 267326 -3856
rect 267562 -4092 267646 -3856
rect 267882 -4092 303326 -3856
rect 303562 -4092 303646 -3856
rect 303882 -4092 339326 -3856
rect 339562 -4092 339646 -3856
rect 339882 -4092 375326 -3856
rect 375562 -4092 375646 -3856
rect 375882 -4092 411326 -3856
rect 411562 -4092 411646 -3856
rect 411882 -4092 447326 -3856
rect 447562 -4092 447646 -3856
rect 447882 -4092 483326 -3856
rect 483562 -4092 483646 -3856
rect 483882 -4092 519326 -3856
rect 519562 -4092 519646 -3856
rect 519882 -4092 555326 -3856
rect 555562 -4092 555646 -3856
rect 555882 -4092 588532 -3856
rect 588768 -4092 588852 -3856
rect 589088 -4092 589120 -3856
rect -5196 -4124 589120 -4092
rect -6156 -4496 590080 -4464
rect -6156 -4732 -6124 -4496
rect -5888 -4732 -5804 -4496
rect -5568 -4732 19826 -4496
rect 20062 -4732 20146 -4496
rect 20382 -4732 55826 -4496
rect 56062 -4732 56146 -4496
rect 56382 -4732 91826 -4496
rect 92062 -4732 92146 -4496
rect 92382 -4732 127826 -4496
rect 128062 -4732 128146 -4496
rect 128382 -4732 163826 -4496
rect 164062 -4732 164146 -4496
rect 164382 -4732 199826 -4496
rect 200062 -4732 200146 -4496
rect 200382 -4732 235826 -4496
rect 236062 -4732 236146 -4496
rect 236382 -4732 271826 -4496
rect 272062 -4732 272146 -4496
rect 272382 -4732 307826 -4496
rect 308062 -4732 308146 -4496
rect 308382 -4732 343826 -4496
rect 344062 -4732 344146 -4496
rect 344382 -4732 379826 -4496
rect 380062 -4732 380146 -4496
rect 380382 -4732 415826 -4496
rect 416062 -4732 416146 -4496
rect 416382 -4732 451826 -4496
rect 452062 -4732 452146 -4496
rect 452382 -4732 487826 -4496
rect 488062 -4732 488146 -4496
rect 488382 -4732 523826 -4496
rect 524062 -4732 524146 -4496
rect 524382 -4732 559826 -4496
rect 560062 -4732 560146 -4496
rect 560382 -4732 589492 -4496
rect 589728 -4732 589812 -4496
rect 590048 -4732 590080 -4496
rect -6156 -4816 590080 -4732
rect -6156 -5052 -6124 -4816
rect -5888 -5052 -5804 -4816
rect -5568 -5052 19826 -4816
rect 20062 -5052 20146 -4816
rect 20382 -5052 55826 -4816
rect 56062 -5052 56146 -4816
rect 56382 -5052 91826 -4816
rect 92062 -5052 92146 -4816
rect 92382 -5052 127826 -4816
rect 128062 -5052 128146 -4816
rect 128382 -5052 163826 -4816
rect 164062 -5052 164146 -4816
rect 164382 -5052 199826 -4816
rect 200062 -5052 200146 -4816
rect 200382 -5052 235826 -4816
rect 236062 -5052 236146 -4816
rect 236382 -5052 271826 -4816
rect 272062 -5052 272146 -4816
rect 272382 -5052 307826 -4816
rect 308062 -5052 308146 -4816
rect 308382 -5052 343826 -4816
rect 344062 -5052 344146 -4816
rect 344382 -5052 379826 -4816
rect 380062 -5052 380146 -4816
rect 380382 -5052 415826 -4816
rect 416062 -5052 416146 -4816
rect 416382 -5052 451826 -4816
rect 452062 -5052 452146 -4816
rect 452382 -5052 487826 -4816
rect 488062 -5052 488146 -4816
rect 488382 -5052 523826 -4816
rect 524062 -5052 524146 -4816
rect 524382 -5052 559826 -4816
rect 560062 -5052 560146 -4816
rect 560382 -5052 589492 -4816
rect 589728 -5052 589812 -4816
rect 590048 -5052 590080 -4816
rect -6156 -5084 590080 -5052
rect -7116 -5456 591040 -5424
rect -7116 -5692 -7084 -5456
rect -6848 -5692 -6764 -5456
rect -6528 -5692 24326 -5456
rect 24562 -5692 24646 -5456
rect 24882 -5692 60326 -5456
rect 60562 -5692 60646 -5456
rect 60882 -5692 96326 -5456
rect 96562 -5692 96646 -5456
rect 96882 -5692 132326 -5456
rect 132562 -5692 132646 -5456
rect 132882 -5692 168326 -5456
rect 168562 -5692 168646 -5456
rect 168882 -5692 204326 -5456
rect 204562 -5692 204646 -5456
rect 204882 -5692 240326 -5456
rect 240562 -5692 240646 -5456
rect 240882 -5692 276326 -5456
rect 276562 -5692 276646 -5456
rect 276882 -5692 312326 -5456
rect 312562 -5692 312646 -5456
rect 312882 -5692 348326 -5456
rect 348562 -5692 348646 -5456
rect 348882 -5692 384326 -5456
rect 384562 -5692 384646 -5456
rect 384882 -5692 420326 -5456
rect 420562 -5692 420646 -5456
rect 420882 -5692 456326 -5456
rect 456562 -5692 456646 -5456
rect 456882 -5692 492326 -5456
rect 492562 -5692 492646 -5456
rect 492882 -5692 528326 -5456
rect 528562 -5692 528646 -5456
rect 528882 -5692 564326 -5456
rect 564562 -5692 564646 -5456
rect 564882 -5692 590452 -5456
rect 590688 -5692 590772 -5456
rect 591008 -5692 591040 -5456
rect -7116 -5776 591040 -5692
rect -7116 -6012 -7084 -5776
rect -6848 -6012 -6764 -5776
rect -6528 -6012 24326 -5776
rect 24562 -6012 24646 -5776
rect 24882 -6012 60326 -5776
rect 60562 -6012 60646 -5776
rect 60882 -6012 96326 -5776
rect 96562 -6012 96646 -5776
rect 96882 -6012 132326 -5776
rect 132562 -6012 132646 -5776
rect 132882 -6012 168326 -5776
rect 168562 -6012 168646 -5776
rect 168882 -6012 204326 -5776
rect 204562 -6012 204646 -5776
rect 204882 -6012 240326 -5776
rect 240562 -6012 240646 -5776
rect 240882 -6012 276326 -5776
rect 276562 -6012 276646 -5776
rect 276882 -6012 312326 -5776
rect 312562 -6012 312646 -5776
rect 312882 -6012 348326 -5776
rect 348562 -6012 348646 -5776
rect 348882 -6012 384326 -5776
rect 384562 -6012 384646 -5776
rect 384882 -6012 420326 -5776
rect 420562 -6012 420646 -5776
rect 420882 -6012 456326 -5776
rect 456562 -6012 456646 -5776
rect 456882 -6012 492326 -5776
rect 492562 -6012 492646 -5776
rect 492882 -6012 528326 -5776
rect 528562 -6012 528646 -5776
rect 528882 -6012 564326 -5776
rect 564562 -6012 564646 -5776
rect 564882 -6012 590452 -5776
rect 590688 -6012 590772 -5776
rect 591008 -6012 591040 -5776
rect -7116 -6044 591040 -6012
rect -8076 -6416 592000 -6384
rect -8076 -6652 -8044 -6416
rect -7808 -6652 -7724 -6416
rect -7488 -6652 28826 -6416
rect 29062 -6652 29146 -6416
rect 29382 -6652 64826 -6416
rect 65062 -6652 65146 -6416
rect 65382 -6652 100826 -6416
rect 101062 -6652 101146 -6416
rect 101382 -6652 136826 -6416
rect 137062 -6652 137146 -6416
rect 137382 -6652 172826 -6416
rect 173062 -6652 173146 -6416
rect 173382 -6652 208826 -6416
rect 209062 -6652 209146 -6416
rect 209382 -6652 244826 -6416
rect 245062 -6652 245146 -6416
rect 245382 -6652 280826 -6416
rect 281062 -6652 281146 -6416
rect 281382 -6652 316826 -6416
rect 317062 -6652 317146 -6416
rect 317382 -6652 352826 -6416
rect 353062 -6652 353146 -6416
rect 353382 -6652 388826 -6416
rect 389062 -6652 389146 -6416
rect 389382 -6652 424826 -6416
rect 425062 -6652 425146 -6416
rect 425382 -6652 460826 -6416
rect 461062 -6652 461146 -6416
rect 461382 -6652 496826 -6416
rect 497062 -6652 497146 -6416
rect 497382 -6652 532826 -6416
rect 533062 -6652 533146 -6416
rect 533382 -6652 568826 -6416
rect 569062 -6652 569146 -6416
rect 569382 -6652 591412 -6416
rect 591648 -6652 591732 -6416
rect 591968 -6652 592000 -6416
rect -8076 -6736 592000 -6652
rect -8076 -6972 -8044 -6736
rect -7808 -6972 -7724 -6736
rect -7488 -6972 28826 -6736
rect 29062 -6972 29146 -6736
rect 29382 -6972 64826 -6736
rect 65062 -6972 65146 -6736
rect 65382 -6972 100826 -6736
rect 101062 -6972 101146 -6736
rect 101382 -6972 136826 -6736
rect 137062 -6972 137146 -6736
rect 137382 -6972 172826 -6736
rect 173062 -6972 173146 -6736
rect 173382 -6972 208826 -6736
rect 209062 -6972 209146 -6736
rect 209382 -6972 244826 -6736
rect 245062 -6972 245146 -6736
rect 245382 -6972 280826 -6736
rect 281062 -6972 281146 -6736
rect 281382 -6972 316826 -6736
rect 317062 -6972 317146 -6736
rect 317382 -6972 352826 -6736
rect 353062 -6972 353146 -6736
rect 353382 -6972 388826 -6736
rect 389062 -6972 389146 -6736
rect 389382 -6972 424826 -6736
rect 425062 -6972 425146 -6736
rect 425382 -6972 460826 -6736
rect 461062 -6972 461146 -6736
rect 461382 -6972 496826 -6736
rect 497062 -6972 497146 -6736
rect 497382 -6972 532826 -6736
rect 533062 -6972 533146 -6736
rect 533382 -6972 568826 -6736
rect 569062 -6972 569146 -6736
rect 569382 -6972 591412 -6736
rect 591648 -6972 591732 -6736
rect 591968 -6972 592000 -6736
rect -8076 -7004 592000 -6972
rect -9036 -7376 592960 -7344
rect -9036 -7612 -9004 -7376
rect -8768 -7612 -8684 -7376
rect -8448 -7612 33326 -7376
rect 33562 -7612 33646 -7376
rect 33882 -7612 69326 -7376
rect 69562 -7612 69646 -7376
rect 69882 -7612 105326 -7376
rect 105562 -7612 105646 -7376
rect 105882 -7612 141326 -7376
rect 141562 -7612 141646 -7376
rect 141882 -7612 177326 -7376
rect 177562 -7612 177646 -7376
rect 177882 -7612 213326 -7376
rect 213562 -7612 213646 -7376
rect 213882 -7612 249326 -7376
rect 249562 -7612 249646 -7376
rect 249882 -7612 285326 -7376
rect 285562 -7612 285646 -7376
rect 285882 -7612 321326 -7376
rect 321562 -7612 321646 -7376
rect 321882 -7612 357326 -7376
rect 357562 -7612 357646 -7376
rect 357882 -7612 393326 -7376
rect 393562 -7612 393646 -7376
rect 393882 -7612 429326 -7376
rect 429562 -7612 429646 -7376
rect 429882 -7612 465326 -7376
rect 465562 -7612 465646 -7376
rect 465882 -7612 501326 -7376
rect 501562 -7612 501646 -7376
rect 501882 -7612 537326 -7376
rect 537562 -7612 537646 -7376
rect 537882 -7612 573326 -7376
rect 573562 -7612 573646 -7376
rect 573882 -7612 592372 -7376
rect 592608 -7612 592692 -7376
rect 592928 -7612 592960 -7376
rect -9036 -7696 592960 -7612
rect -9036 -7932 -9004 -7696
rect -8768 -7932 -8684 -7696
rect -8448 -7932 33326 -7696
rect 33562 -7932 33646 -7696
rect 33882 -7932 69326 -7696
rect 69562 -7932 69646 -7696
rect 69882 -7932 105326 -7696
rect 105562 -7932 105646 -7696
rect 105882 -7932 141326 -7696
rect 141562 -7932 141646 -7696
rect 141882 -7932 177326 -7696
rect 177562 -7932 177646 -7696
rect 177882 -7932 213326 -7696
rect 213562 -7932 213646 -7696
rect 213882 -7932 249326 -7696
rect 249562 -7932 249646 -7696
rect 249882 -7932 285326 -7696
rect 285562 -7932 285646 -7696
rect 285882 -7932 321326 -7696
rect 321562 -7932 321646 -7696
rect 321882 -7932 357326 -7696
rect 357562 -7932 357646 -7696
rect 357882 -7932 393326 -7696
rect 393562 -7932 393646 -7696
rect 393882 -7932 429326 -7696
rect 429562 -7932 429646 -7696
rect 429882 -7932 465326 -7696
rect 465562 -7932 465646 -7696
rect 465882 -7932 501326 -7696
rect 501562 -7932 501646 -7696
rect 501882 -7932 537326 -7696
rect 537562 -7932 537646 -7696
rect 537882 -7932 573326 -7696
rect 573562 -7932 573646 -7696
rect 573882 -7932 592372 -7696
rect 592608 -7932 592692 -7696
rect 592928 -7932 592960 -7696
rect -9036 -7964 592960 -7932
use sky130_sram_2kbyte_1rw1r_32x512_8  dram_inst
timestamp 0
transform 1 0 220000 0 1 480000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  iram_inst
timestamp 0
transform 1 0 220000 0 1 160000
box 0 0 136620 83308
use rvj1_caravel_soc  rvj1_soc
timestamp 0
transform 1 0 232400 0 1 310400
box 13 0 128970 131144
use wbuart_wrap  uart_inst
timestamp 0
transform 1 0 100000 0 1 300000
box 0 0 70020 72164
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal4 s -2316 -1244 -1696 705180 4 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2316 -1244 586240 -624 8 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2316 704560 586240 705180 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 585620 -1244 586240 705180 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 1794 -7964 2414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 37794 -7964 38414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 73794 -7964 74414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 109794 -7964 110414 298000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 109794 374164 110414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 145794 -7964 146414 298000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 145794 374164 146414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 181794 -7964 182414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 217794 -7964 218414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 217794 245308 218414 478000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 217794 565308 218414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 253794 -7964 254414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 253794 245308 254414 308400 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 253794 565308 254414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 289794 -7964 290414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 289794 245308 290414 308400 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 289794 565308 290414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 -7964 326414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 245308 326414 308400 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 565308 326414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 361794 -7964 362414 308400 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 361794 443544 362414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 397794 -7964 398414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 433794 -7964 434414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 469794 -7964 470414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 505794 -7964 506414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 541794 -7964 542414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 577794 -7964 578414 711900 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 2866 592960 3486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 38866 592960 39486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 74866 592960 75486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 110866 592960 111486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 146866 592960 147486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 182866 592960 183486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 218866 592960 219486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 254866 592960 255486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 290866 592960 291486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 326866 592960 327486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 362866 592960 363486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 398866 592960 399486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 434866 592960 435486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 470866 592960 471486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 506866 592960 507486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 542866 592960 543486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 578866 592960 579486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 614866 592960 615486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 650866 592960 651486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -9036 686866 592960 687486 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s -4236 -3164 -3616 707100 4 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -4236 -3164 588160 -2544 8 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -4236 706480 588160 707100 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 587540 -3164 588160 707100 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 10794 -7964 11414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 46794 -7964 47414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 82794 -7964 83414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 118794 -7964 119414 298000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 118794 374164 119414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 154794 -7964 155414 298000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 154794 374164 155414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 190794 -7964 191414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 226794 -7964 227414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 226794 245308 227414 478000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 226794 565308 227414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 262794 -7964 263414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 262794 245308 263414 308400 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 262794 565308 263414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 298794 -7964 299414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 298794 245308 299414 308400 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 298794 565308 299414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 334794 -7964 335414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 334794 245308 335414 308400 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 334794 565308 335414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 370794 -7964 371414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 406794 -7964 407414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 442794 -7964 443414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 478794 -7964 479414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 514794 -7964 515414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 550794 -7964 551414 711900 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 11866 592960 12486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 47866 592960 48486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 83866 592960 84486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 119866 592960 120486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 155866 592960 156486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 191866 592960 192486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 227866 592960 228486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 263866 592960 264486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 299866 592960 300486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 335866 592960 336486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 371866 592960 372486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 407866 592960 408486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 443866 592960 444486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 479866 592960 480486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 515866 592960 516486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 551866 592960 552486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 587866 592960 588486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 623866 592960 624486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 659866 592960 660486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -9036 695866 592960 696486 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s -5196 -4124 -4576 708060 4 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -5196 -4124 589120 -3504 8 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -5196 707440 589120 708060 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 588500 -4124 589120 708060 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 15294 -7964 15914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 51294 -7964 51914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 87294 -7964 87914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 123294 -7964 123914 298000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 123294 374164 123914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 159294 -7964 159914 298000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 159294 374164 159914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 195294 -7964 195914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 231294 -7964 231914 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 231294 245308 231914 308400 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 231294 565308 231914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 267294 -7964 267914 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 267294 245308 267914 308400 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 267294 565308 267914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 303294 -7964 303914 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 303294 245308 303914 308400 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 303294 565308 303914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 339294 -7964 339914 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 339294 245308 339914 308400 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 339294 565308 339914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 375294 -7964 375914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 411294 -7964 411914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 447294 -7964 447914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 483294 -7964 483914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 519294 -7964 519914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 555294 -7964 555914 711900 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 16366 592960 16986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 52366 592960 52986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 88366 592960 88986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 124366 592960 124986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 160366 592960 160986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 196366 592960 196986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 232366 592960 232986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 268366 592960 268986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 304366 592960 304986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 340366 592960 340986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 376366 592960 376986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 412366 592960 412986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 448366 592960 448986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 484366 592960 484986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 520366 592960 520986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 556366 592960 556986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 592366 592960 592986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 628366 592960 628986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 664366 592960 664986 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -9036 700366 592960 700986 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s -6156 -5084 -5536 709020 4 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -6156 -5084 590080 -4464 8 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -6156 708400 590080 709020 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 589460 -5084 590080 709020 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 19794 -7964 20414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 55794 -7964 56414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 91794 -7964 92414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 127794 -7964 128414 298000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 127794 374164 128414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 163794 -7964 164414 298000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 163794 374164 164414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 199794 -7964 200414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 235794 -7964 236414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 235794 565308 236414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 271794 -7964 272414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 271794 565308 272414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 307794 -7964 308414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 307794 565308 308414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 343794 -7964 344414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 343794 565308 344414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 379794 -7964 380414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 415794 -7964 416414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 451794 -7964 452414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 487794 -7964 488414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 523794 -7964 524414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 559794 -7964 560414 711900 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 20866 592960 21486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 56866 592960 57486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 92866 592960 93486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 128866 592960 129486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 164866 592960 165486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 200866 592960 201486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 236866 592960 237486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 272866 592960 273486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 308866 592960 309486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 344866 592960 345486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 380866 592960 381486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 416866 592960 417486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 452866 592960 453486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 488866 592960 489486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 524866 592960 525486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 560866 592960 561486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 596866 592960 597486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 632866 592960 633486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -9036 668866 592960 669486 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s -8076 -7004 -7456 710940 4 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8076 -7004 592000 -6384 8 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8076 710320 592000 710940 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 591380 -7004 592000 710940 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 28794 -7964 29414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 64794 -7964 65414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 100794 -7964 101414 298000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 100794 374164 101414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 136794 -7964 137414 298000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 136794 374164 137414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 172794 -7964 173414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 208794 -7964 209414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 244794 -7964 245414 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 244794 245308 245414 308400 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 244794 565308 245414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 280794 -7964 281414 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 280794 245308 281414 308400 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 280794 565308 281414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 316794 -7964 317414 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 316794 245308 317414 308400 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 316794 565308 317414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 352794 -7964 353414 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 352794 245308 353414 308400 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 352794 565308 353414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 388794 -7964 389414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 424794 -7964 425414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 460794 -7964 461414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 496794 -7964 497414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 532794 -7964 533414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 568794 -7964 569414 711900 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 29866 592960 30486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 65866 592960 66486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 101866 592960 102486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 137866 592960 138486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 173866 592960 174486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 209866 592960 210486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 245866 592960 246486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 281866 592960 282486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 317866 592960 318486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 353866 592960 354486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 389866 592960 390486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 425866 592960 426486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 461866 592960 462486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 497866 592960 498486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 533866 592960 534486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 569866 592960 570486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 605866 592960 606486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 641866 592960 642486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -9036 677866 592960 678486 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s -9036 -7964 -8416 711900 4 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 -7964 592960 -7344 8 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 711280 592960 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 592340 -7964 592960 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 33294 -7964 33914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 69294 -7964 69914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 105294 -7964 105914 298000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 105294 374164 105914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 141294 -7964 141914 298000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 141294 374164 141914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 177294 -7964 177914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 213294 -7964 213914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 249294 -7964 249914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 249294 245308 249914 308400 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 249294 565308 249914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 285294 -7964 285914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 285294 245308 285914 308400 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 285294 565308 285914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 321294 -7964 321914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 321294 245308 321914 308400 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 321294 565308 321914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 357294 -7964 357914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 357294 245308 357914 308400 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 357294 565308 357914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 393294 -7964 393914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 429294 -7964 429914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 465294 -7964 465914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 501294 -7964 501914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 537294 -7964 537914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 573294 -7964 573914 711900 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 34366 592960 34986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 70366 592960 70986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 106366 592960 106986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 142366 592960 142986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 178366 592960 178986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 214366 592960 214986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 250366 592960 250986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 286366 592960 286986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 322366 592960 322986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 358366 592960 358986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 394366 592960 394986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 430366 592960 430986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 466366 592960 466986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 502366 592960 502986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 538366 592960 538986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 574366 592960 574986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 610366 592960 610986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 646366 592960 646986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -9036 682366 592960 682986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s -3276 -2204 -2656 706140 4 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -3276 -2204 587200 -1584 8 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -3276 705520 587200 706140 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 586580 -2204 587200 706140 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 6294 -7964 6914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 42294 -7964 42914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 78294 -7964 78914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 114294 -7964 114914 298000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 114294 374164 114914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 150294 -7964 150914 298000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 150294 374164 150914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 186294 -7964 186914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 222294 -7964 222914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 222294 245308 222914 478000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 222294 565308 222914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 258294 -7964 258914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 258294 245308 258914 308400 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 258294 565308 258914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 294294 -7964 294914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 294294 245308 294914 308400 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 294294 565308 294914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 330294 -7964 330914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 330294 245308 330914 308400 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 330294 565308 330914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 366294 -7964 366914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 402294 -7964 402914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 438294 -7964 438914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 474294 -7964 474914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 510294 -7964 510914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 546294 -7964 546914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 582294 -7964 582914 711900 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 7366 592960 7986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 43366 592960 43986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 79366 592960 79986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 115366 592960 115986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 151366 592960 151986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 187366 592960 187986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 223366 592960 223986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 259366 592960 259986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 295366 592960 295986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 331366 592960 331986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 367366 592960 367986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 403366 592960 403986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 439366 592960 439986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 475366 592960 475986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 511366 592960 511986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 547366 592960 547986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 583366 592960 583986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 619366 592960 619986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 655366 592960 655986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -9036 691366 592960 691986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s -7116 -6044 -6496 709980 4 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -7116 -6044 591040 -5424 8 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -7116 709360 591040 709980 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 590420 -6044 591040 709980 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 24294 -7964 24914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 60294 -7964 60914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 96294 -7964 96914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 132294 -7964 132914 298000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 132294 374164 132914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 168294 -7964 168914 298000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 168294 374164 168914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 204294 -7964 204914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 240294 -7964 240914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 240294 565308 240914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 276294 -7964 276914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 276294 565308 276914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 312294 -7964 312914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 312294 565308 312914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 348294 -7964 348914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 348294 565308 348914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 384294 -7964 384914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 420294 -7964 420914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 456294 -7964 456914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 492294 -7964 492914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 528294 -7964 528914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 564294 -7964 564914 711900 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 25366 592960 25986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 61366 592960 61986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 97366 592960 97986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 133366 592960 133986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 169366 592960 169986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 205366 592960 205986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 241366 592960 241986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 277366 592960 277986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 313366 592960 313986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 349366 592960 349986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 385366 592960 385986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 421366 592960 421986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 457366 592960 457986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 493366 592960 493986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 529366 592960 529986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 565366 592960 565986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 601366 592960 601986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 637366 592960 637986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -9036 673366 592960 673986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
