magic
tech sky130A
magscale 1 2
timestamp 1654606772
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 348786 700476 348792 700528
rect 348844 700516 348850 700528
rect 358906 700516 358912 700528
rect 348844 700488 358912 700516
rect 348844 700476 348850 700488
rect 358906 700476 358912 700488
rect 358964 700476 358970 700528
rect 300118 700408 300124 700460
rect 300176 700448 300182 700460
rect 357526 700448 357532 700460
rect 300176 700420 357532 700448
rect 300176 700408 300182 700420
rect 357526 700408 357532 700420
rect 357584 700408 357590 700460
rect 283834 700340 283840 700392
rect 283892 700380 283898 700392
rect 358814 700380 358820 700392
rect 283892 700352 358820 700380
rect 283892 700340 283898 700352
rect 358814 700340 358820 700352
rect 358872 700340 358878 700392
rect 359458 700340 359464 700392
rect 359516 700380 359522 700392
rect 397454 700380 397460 700392
rect 359516 700352 397460 700380
rect 359516 700340 359522 700352
rect 397454 700340 397460 700352
rect 397512 700340 397518 700392
rect 267642 700272 267648 700324
rect 267700 700312 267706 700324
rect 357434 700312 357440 700324
rect 267700 700284 357440 700312
rect 267700 700272 267706 700284
rect 357434 700272 357440 700284
rect 357492 700272 357498 700324
rect 358078 700272 358084 700324
rect 358136 700312 358142 700324
rect 559650 700312 559656 700324
rect 358136 700284 559656 700312
rect 358136 700272 358142 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 360838 699660 360844 699712
rect 360896 699700 360902 699712
rect 364978 699700 364984 699712
rect 360896 699672 364984 699700
rect 360896 699660 360902 699672
rect 364978 699660 364984 699672
rect 365036 699660 365042 699712
rect 359550 696940 359556 696992
rect 359608 696980 359614 696992
rect 580166 696980 580172 696992
rect 359608 696952 580172 696980
rect 359608 696940 359614 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 2774 683680 2780 683732
rect 2832 683720 2838 683732
rect 4798 683720 4804 683732
rect 2832 683692 4804 683720
rect 2832 683680 2838 683692
rect 4798 683680 4804 683692
rect 4856 683680 4862 683732
rect 358170 670692 358176 670744
rect 358228 670732 358234 670744
rect 580166 670732 580172 670744
rect 358228 670704 580172 670732
rect 358228 670692 358234 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3510 656888 3516 656940
rect 3568 656928 3574 656940
rect 178678 656928 178684 656940
rect 3568 656900 178684 656928
rect 3568 656888 3574 656900
rect 178678 656888 178684 656900
rect 178736 656888 178742 656940
rect 2774 632068 2780 632120
rect 2832 632108 2838 632120
rect 4890 632108 4896 632120
rect 2832 632080 4896 632108
rect 2832 632068 2838 632080
rect 4890 632068 4896 632080
rect 4948 632068 4954 632120
rect 362218 630640 362224 630692
rect 362276 630680 362282 630692
rect 580166 630680 580172 630692
rect 362276 630652 580172 630680
rect 362276 630640 362282 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 359642 616836 359648 616888
rect 359700 616876 359706 616888
rect 580166 616876 580172 616888
rect 359700 616848 580172 616876
rect 359700 616836 359706 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3326 605820 3332 605872
rect 3384 605860 3390 605872
rect 203518 605860 203524 605872
rect 3384 605832 203524 605860
rect 3384 605820 3390 605832
rect 203518 605820 203524 605832
rect 203576 605820 203582 605872
rect 362310 590656 362316 590708
rect 362368 590696 362374 590708
rect 579614 590696 579620 590708
rect 362368 590668 579620 590696
rect 362368 590656 362374 590668
rect 579614 590656 579620 590668
rect 579672 590656 579678 590708
rect 2774 579912 2780 579964
rect 2832 579952 2838 579964
rect 4982 579952 4988 579964
rect 2832 579924 4988 579952
rect 2832 579912 2838 579924
rect 4982 579912 4988 579924
rect 5040 579912 5046 579964
rect 3050 565836 3056 565888
rect 3108 565876 3114 565888
rect 31018 565876 31024 565888
rect 3108 565848 31024 565876
rect 3108 565836 3114 565848
rect 31018 565836 31024 565848
rect 31076 565836 31082 565888
rect 217962 565088 217968 565140
rect 218020 565128 218026 565140
rect 234614 565128 234620 565140
rect 218020 565100 234620 565128
rect 218020 565088 218026 565100
rect 234614 565088 234620 565100
rect 234672 565088 234678 565140
rect 331214 565088 331220 565140
rect 331272 565128 331278 565140
rect 358998 565128 359004 565140
rect 331272 565100 359004 565128
rect 331272 565088 331278 565100
rect 358998 565088 359004 565100
rect 359056 565088 359062 565140
rect 371878 563048 371884 563100
rect 371936 563088 371942 563100
rect 580166 563088 580172 563100
rect 371936 563060 580172 563088
rect 371936 563048 371942 563060
rect 580166 563048 580172 563060
rect 580224 563048 580230 563100
rect 2774 553664 2780 553716
rect 2832 553704 2838 553716
rect 5074 553704 5080 553716
rect 2832 553676 5080 553704
rect 2832 553664 2838 553676
rect 5074 553664 5080 553676
rect 5132 553664 5138 553716
rect 358262 536800 358268 536852
rect 358320 536840 358326 536852
rect 580166 536840 580172 536852
rect 358320 536812 580172 536840
rect 358320 536800 358326 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 3326 527756 3332 527808
rect 3384 527796 3390 527808
rect 8938 527796 8944 527808
rect 3384 527768 8944 527796
rect 3384 527756 3390 527768
rect 8938 527756 8944 527768
rect 8996 527756 9002 527808
rect 358354 484372 358360 484424
rect 358412 484412 358418 484424
rect 580166 484412 580172 484424
rect 358412 484384 580172 484412
rect 358412 484372 358418 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 217410 478864 217416 478916
rect 217468 478904 217474 478916
rect 220078 478904 220084 478916
rect 217468 478876 220084 478904
rect 217468 478864 217474 478876
rect 220078 478864 220084 478876
rect 220136 478864 220142 478916
rect 311894 478184 311900 478236
rect 311952 478224 311958 478236
rect 358906 478224 358912 478236
rect 311952 478196 358912 478224
rect 311952 478184 311958 478196
rect 358906 478184 358912 478196
rect 358964 478184 358970 478236
rect 3694 478116 3700 478168
rect 3752 478156 3758 478168
rect 354674 478156 354680 478168
rect 3752 478128 354680 478156
rect 3752 478116 3758 478128
rect 354674 478116 354680 478128
rect 354732 478116 354738 478168
rect 280246 476688 280252 476740
rect 280304 476728 280310 476740
rect 302234 476728 302240 476740
rect 280304 476700 302240 476728
rect 280304 476688 280310 476700
rect 302234 476688 302240 476700
rect 302292 476688 302298 476740
rect 241606 476620 241612 476672
rect 241664 476660 241670 476672
rect 252554 476660 252560 476672
rect 241664 476632 252560 476660
rect 241664 476620 241670 476632
rect 252554 476620 252560 476632
rect 252612 476620 252618 476672
rect 255406 476620 255412 476672
rect 255464 476660 255470 476672
rect 264974 476660 264980 476672
rect 255464 476632 264980 476660
rect 255464 476620 255470 476632
rect 264974 476620 264980 476632
rect 265032 476620 265038 476672
rect 281534 476620 281540 476672
rect 281592 476660 281598 476672
rect 304994 476660 305000 476672
rect 281592 476632 305000 476660
rect 281592 476620 281598 476632
rect 304994 476620 305000 476632
rect 305052 476620 305058 476672
rect 259546 476552 259552 476604
rect 259604 476592 259610 476604
rect 270494 476592 270500 476604
rect 259604 476564 270500 476592
rect 259604 476552 259610 476564
rect 270494 476552 270500 476564
rect 270552 476552 270558 476604
rect 283098 476552 283104 476604
rect 283156 476592 283162 476604
rect 307754 476592 307760 476604
rect 283156 476564 307760 476592
rect 283156 476552 283162 476564
rect 307754 476552 307760 476564
rect 307812 476552 307818 476604
rect 238754 476484 238760 476536
rect 238812 476524 238818 476536
rect 244274 476524 244280 476536
rect 238812 476496 244280 476524
rect 238812 476484 238818 476496
rect 244274 476484 244280 476496
rect 244332 476484 244338 476536
rect 249794 476524 249800 476536
rect 248386 476496 249800 476524
rect 236086 476416 236092 476468
rect 236144 476456 236150 476468
rect 247034 476456 247040 476468
rect 236144 476428 247040 476456
rect 236144 476416 236150 476428
rect 247034 476416 247040 476428
rect 247092 476416 247098 476468
rect 238846 476348 238852 476400
rect 238904 476388 238910 476400
rect 248386 476388 248414 476496
rect 249794 476484 249800 476496
rect 249852 476484 249858 476536
rect 252646 476484 252652 476536
rect 252704 476524 252710 476536
rect 263594 476524 263600 476536
rect 252704 476496 263600 476524
rect 252704 476484 252710 476496
rect 263594 476484 263600 476496
rect 263652 476484 263658 476536
rect 265066 476484 265072 476536
rect 265124 476524 265130 476536
rect 280154 476524 280160 476536
rect 265124 476496 280160 476524
rect 265124 476484 265130 476496
rect 280154 476484 280160 476496
rect 280212 476484 280218 476536
rect 284294 476484 284300 476536
rect 284352 476524 284358 476536
rect 310514 476524 310520 476536
rect 284352 476496 310520 476524
rect 284352 476484 284358 476496
rect 310514 476484 310520 476496
rect 310572 476484 310578 476536
rect 251174 476416 251180 476468
rect 251232 476456 251238 476468
rect 260834 476456 260840 476468
rect 251232 476428 260840 476456
rect 251232 476416 251238 476428
rect 260834 476416 260840 476428
rect 260892 476416 260898 476468
rect 268010 476456 268016 476468
rect 260944 476428 268016 476456
rect 238904 476360 248414 476388
rect 238904 476348 238910 476360
rect 258166 476348 258172 476400
rect 258224 476388 258230 476400
rect 260944 476388 260972 476428
rect 268010 476416 268016 476428
rect 268068 476416 268074 476468
rect 285674 476416 285680 476468
rect 285732 476456 285738 476468
rect 313274 476456 313280 476468
rect 285732 476428 313280 476456
rect 285732 476416 285738 476428
rect 313274 476416 313280 476428
rect 313332 476416 313338 476468
rect 273254 476388 273260 476400
rect 258224 476360 260972 476388
rect 261036 476360 273260 476388
rect 258224 476348 258230 476360
rect 234706 476280 234712 476332
rect 234764 476320 234770 476332
rect 242894 476320 242900 476332
rect 234764 476292 242900 476320
rect 234764 476280 234770 476292
rect 242894 476280 242900 476292
rect 242952 476280 242958 476332
rect 245746 476280 245752 476332
rect 245804 476320 245810 476332
rect 255314 476320 255320 476332
rect 245804 476292 255320 476320
rect 245804 476280 245810 476292
rect 255314 476280 255320 476292
rect 255372 476280 255378 476332
rect 255424 476292 256924 476320
rect 241514 476212 241520 476264
rect 241572 476252 241578 476264
rect 244274 476252 244280 476264
rect 241572 476224 244280 476252
rect 241572 476212 241578 476224
rect 244274 476212 244280 476224
rect 244332 476212 244338 476264
rect 248414 476212 248420 476264
rect 248472 476252 248478 476264
rect 255424 476252 255452 476292
rect 248472 476224 255452 476252
rect 248472 476212 248478 476224
rect 242802 476144 242808 476196
rect 242860 476184 242866 476196
rect 244918 476184 244924 476196
rect 242860 476156 244924 476184
rect 242860 476144 242866 476156
rect 244918 476144 244924 476156
rect 244976 476144 244982 476196
rect 252370 476144 252376 476196
rect 252428 476184 252434 476196
rect 256694 476184 256700 476196
rect 252428 476156 256700 476184
rect 252428 476144 252434 476156
rect 256694 476144 256700 476156
rect 256752 476144 256758 476196
rect 256896 476184 256924 476292
rect 260926 476280 260932 476332
rect 260984 476320 260990 476332
rect 261036 476320 261064 476360
rect 273254 476348 273260 476360
rect 273312 476348 273318 476400
rect 287238 476348 287244 476400
rect 287296 476388 287302 476400
rect 314654 476388 314660 476400
rect 287296 476360 314660 476388
rect 287296 476348 287302 476360
rect 314654 476348 314660 476360
rect 314712 476348 314718 476400
rect 260984 476292 261064 476320
rect 260984 476280 260990 476292
rect 263686 476280 263692 476332
rect 263744 476320 263750 476332
rect 277854 476320 277860 476332
rect 263744 476292 277860 476320
rect 263744 476280 263750 476292
rect 277854 476280 277860 476292
rect 277912 476280 277918 476332
rect 288526 476280 288532 476332
rect 288584 476320 288590 476332
rect 317414 476320 317420 476332
rect 288584 476292 317420 476320
rect 288584 476280 288590 476292
rect 317414 476280 317420 476292
rect 317472 476280 317478 476332
rect 262398 476212 262404 476264
rect 262456 476252 262462 476264
rect 276014 476252 276020 476264
rect 262456 476224 276020 476252
rect 262456 476212 262462 476224
rect 276014 476212 276020 476224
rect 276072 476212 276078 476264
rect 292758 476212 292764 476264
rect 292816 476252 292822 476264
rect 322934 476252 322940 476264
rect 292816 476224 322940 476252
rect 292816 476212 292822 476224
rect 322934 476212 322940 476224
rect 322992 476212 322998 476264
rect 258258 476184 258264 476196
rect 256896 476156 258264 476184
rect 258258 476144 258264 476156
rect 258316 476144 258322 476196
rect 267734 476144 267740 476196
rect 267792 476184 267798 476196
rect 282914 476184 282920 476196
rect 267792 476156 282920 476184
rect 267792 476144 267798 476156
rect 282914 476144 282920 476156
rect 282972 476144 282978 476196
rect 289998 476144 290004 476196
rect 290056 476184 290062 476196
rect 320174 476184 320180 476196
rect 290056 476156 320180 476184
rect 290056 476144 290062 476156
rect 320174 476144 320180 476156
rect 320232 476144 320238 476196
rect 234614 476076 234620 476128
rect 234672 476116 234678 476128
rect 235902 476116 235908 476128
rect 234672 476088 235908 476116
rect 234672 476076 234678 476088
rect 235902 476076 235908 476088
rect 235960 476076 235966 476128
rect 241422 476076 241428 476128
rect 241480 476116 241486 476128
rect 242894 476116 242900 476128
rect 241480 476088 242900 476116
rect 241480 476076 241486 476088
rect 242894 476076 242900 476088
rect 242952 476076 242958 476128
rect 244274 476076 244280 476128
rect 244332 476116 244338 476128
rect 245654 476116 245660 476128
rect 244332 476088 245660 476116
rect 244332 476076 244338 476088
rect 245654 476076 245660 476088
rect 245712 476076 245718 476128
rect 251082 476076 251088 476128
rect 251140 476116 251146 476128
rect 252554 476116 252560 476128
rect 251140 476088 252560 476116
rect 251140 476076 251146 476088
rect 252554 476076 252560 476088
rect 252612 476076 252618 476128
rect 263502 476076 263508 476128
rect 263560 476116 263566 476128
rect 266998 476116 267004 476128
rect 263560 476088 267004 476116
rect 263560 476076 263566 476088
rect 266998 476076 267004 476088
rect 267056 476076 267062 476128
rect 280062 476076 280068 476128
rect 280120 476116 280126 476128
rect 282178 476116 282184 476128
rect 280120 476088 282184 476116
rect 280120 476076 280126 476088
rect 282178 476076 282184 476088
rect 282236 476076 282242 476128
rect 293954 476076 293960 476128
rect 294012 476116 294018 476128
rect 325786 476116 325792 476128
rect 294012 476088 325792 476116
rect 294012 476076 294018 476088
rect 325786 476076 325792 476088
rect 325844 476076 325850 476128
rect 219066 475396 219072 475448
rect 219124 475436 219130 475448
rect 249886 475436 249892 475448
rect 219124 475408 249892 475436
rect 219124 475396 219130 475408
rect 249886 475396 249892 475408
rect 249944 475396 249950 475448
rect 217594 475328 217600 475380
rect 217652 475368 217658 475380
rect 253934 475368 253940 475380
rect 217652 475340 253940 475368
rect 217652 475328 217658 475340
rect 253934 475328 253940 475340
rect 253992 475328 253998 475380
rect 3326 474716 3332 474768
rect 3384 474756 3390 474768
rect 333974 474756 333980 474768
rect 3384 474728 333980 474756
rect 3384 474716 3390 474728
rect 333974 474716 333980 474728
rect 334032 474716 334038 474768
rect 217502 473968 217508 474020
rect 217560 474008 217566 474020
rect 251266 474008 251272 474020
rect 217560 473980 251272 474008
rect 217560 473968 217566 473980
rect 251266 473968 251272 473980
rect 251324 473968 251330 474020
rect 219158 472608 219164 472660
rect 219216 472648 219222 472660
rect 247126 472648 247132 472660
rect 219216 472620 247132 472648
rect 219216 472608 219222 472620
rect 247126 472608 247132 472620
rect 247184 472608 247190 472660
rect 3418 462340 3424 462392
rect 3476 462380 3482 462392
rect 335354 462380 335360 462392
rect 3476 462352 335360 462380
rect 3476 462340 3482 462352
rect 335354 462340 335360 462352
rect 335412 462340 335418 462392
rect 271966 461660 271972 461712
rect 272024 461700 272030 461712
rect 289906 461700 289912 461712
rect 272024 461672 289912 461700
rect 272024 461660 272030 461672
rect 289906 461660 289912 461672
rect 289964 461660 289970 461712
rect 273254 461592 273260 461644
rect 273312 461632 273318 461644
rect 292666 461632 292672 461644
rect 273312 461604 292672 461632
rect 273312 461592 273318 461604
rect 292666 461592 292672 461604
rect 292724 461592 292730 461644
rect 274542 460300 274548 460352
rect 274600 460340 274606 460352
rect 285122 460340 285128 460352
rect 274600 460312 285128 460340
rect 274600 460300 274606 460312
rect 285122 460300 285128 460312
rect 285180 460300 285186 460352
rect 273162 460232 273168 460284
rect 273220 460272 273226 460284
rect 283006 460272 283012 460284
rect 273220 460244 283012 460272
rect 273220 460232 273226 460244
rect 283006 460232 283012 460244
rect 283064 460232 283070 460284
rect 270586 460164 270592 460216
rect 270644 460204 270650 460216
rect 287146 460204 287152 460216
rect 270644 460176 287152 460204
rect 270644 460164 270650 460176
rect 287146 460164 287152 460176
rect 287204 460164 287210 460216
rect 266262 458940 266268 458992
rect 266320 458980 266326 458992
rect 274634 458980 274640 458992
rect 266320 458952 274640 458980
rect 266320 458940 266326 458952
rect 274634 458940 274640 458952
rect 274692 458940 274698 458992
rect 267550 458872 267556 458924
rect 267608 458912 267614 458924
rect 276014 458912 276020 458924
rect 267608 458884 276020 458912
rect 267608 458872 267614 458884
rect 276014 458872 276020 458884
rect 276072 458872 276078 458924
rect 271782 458804 271788 458856
rect 271840 458844 271846 458856
rect 282086 458844 282092 458856
rect 271840 458816 282092 458844
rect 271840 458804 271846 458816
rect 282086 458804 282092 458816
rect 282144 458804 282150 458856
rect 269022 457716 269028 457768
rect 269080 457756 269086 457768
rect 279050 457756 279056 457768
rect 269080 457728 279056 457756
rect 269080 457716 269086 457728
rect 279050 457716 279056 457728
rect 279108 457716 279114 457768
rect 270402 457648 270408 457700
rect 270460 457688 270466 457700
rect 280522 457688 280528 457700
rect 270460 457660 280528 457688
rect 270460 457648 270466 457660
rect 280522 457648 280528 457660
rect 280580 457648 280586 457700
rect 275186 457580 275192 457632
rect 275244 457620 275250 457632
rect 295334 457620 295340 457632
rect 275244 457592 295340 457620
rect 275244 457580 275250 457592
rect 295334 457580 295340 457592
rect 295392 457580 295398 457632
rect 276566 457512 276572 457564
rect 276624 457552 276630 457564
rect 298094 457552 298100 457564
rect 276624 457524 298100 457552
rect 276624 457512 276630 457524
rect 298094 457512 298100 457524
rect 298152 457512 298158 457564
rect 217870 457444 217876 457496
rect 217928 457484 217934 457496
rect 256786 457484 256792 457496
rect 217928 457456 256792 457484
rect 217928 457444 217934 457456
rect 256786 457444 256792 457456
rect 256844 457444 256850 457496
rect 267642 457444 267648 457496
rect 267700 457484 267706 457496
rect 277394 457484 277400 457496
rect 267700 457456 277400 457484
rect 267700 457444 267706 457456
rect 277394 457444 277400 457456
rect 277452 457444 277458 457496
rect 277946 457444 277952 457496
rect 278004 457484 278010 457496
rect 300854 457484 300860 457496
rect 278004 457456 300860 457484
rect 278004 457444 278010 457456
rect 300854 457444 300860 457456
rect 300912 457444 300918 457496
rect 300854 456220 300860 456272
rect 300912 456260 300918 456272
rect 362218 456260 362224 456272
rect 300912 456232 362224 456260
rect 300912 456220 300918 456232
rect 362218 456220 362224 456232
rect 362276 456220 362282 456272
rect 219250 456152 219256 456204
rect 219308 456192 219314 456204
rect 240962 456192 240968 456204
rect 219308 456164 240968 456192
rect 219308 456152 219314 456164
rect 240962 456152 240968 456164
rect 241020 456152 241026 456204
rect 278682 456152 278688 456204
rect 278740 456192 278746 456204
rect 291378 456192 291384 456204
rect 278740 456164 291384 456192
rect 278740 456152 278746 456164
rect 291378 456152 291384 456164
rect 291436 456152 291442 456204
rect 303154 456152 303160 456204
rect 303212 456192 303218 456204
rect 580258 456192 580264 456204
rect 303212 456164 580264 456192
rect 303212 456152 303218 456164
rect 580258 456152 580264 456164
rect 580316 456152 580322 456204
rect 219342 456084 219348 456136
rect 219400 456124 219406 456136
rect 244366 456124 244372 456136
rect 219400 456096 244372 456124
rect 219400 456084 219406 456096
rect 244366 456084 244372 456096
rect 244424 456084 244430 456136
rect 269206 456084 269212 456136
rect 269264 456124 269270 456136
rect 285766 456124 285772 456136
rect 269264 456096 285772 456124
rect 269264 456084 269270 456096
rect 285766 456084 285772 456096
rect 285824 456084 285830 456136
rect 298370 456084 298376 456136
rect 298428 456124 298434 456136
rect 580442 456124 580448 456136
rect 298428 456096 580448 456124
rect 298428 456084 298434 456096
rect 580442 456084 580448 456096
rect 580500 456084 580506 456136
rect 3602 456016 3608 456068
rect 3660 456056 3666 456068
rect 333514 456056 333520 456068
rect 3660 456028 333520 456056
rect 3660 456016 3666 456028
rect 333514 456016 333520 456028
rect 333572 456016 333578 456068
rect 218054 454928 218060 454980
rect 218112 454968 218118 454980
rect 317414 454968 317420 454980
rect 218112 454940 317420 454968
rect 218112 454928 218118 454940
rect 317414 454928 317420 454940
rect 317472 454928 317478 454980
rect 31018 454860 31024 454912
rect 31076 454900 31082 454912
rect 331214 454900 331220 454912
rect 31076 454872 331220 454900
rect 31076 454860 31082 454872
rect 331214 454860 331220 454872
rect 331272 454860 331278 454912
rect 337378 454860 337384 454912
rect 337436 454900 337442 454912
rect 359458 454900 359464 454912
rect 337436 454872 359464 454900
rect 337436 454860 337442 454872
rect 359458 454860 359464 454872
rect 359516 454860 359522 454912
rect 3326 454792 3332 454844
rect 3384 454832 3390 454844
rect 325694 454832 325700 454844
rect 3384 454804 325700 454832
rect 3384 454792 3390 454804
rect 325694 454792 325700 454804
rect 325752 454792 325758 454844
rect 325786 454792 325792 454844
rect 325844 454832 325850 454844
rect 362310 454832 362316 454844
rect 325844 454804 362316 454832
rect 325844 454792 325850 454804
rect 362310 454792 362316 454804
rect 362368 454792 362374 454844
rect 3510 454724 3516 454776
rect 3568 454764 3574 454776
rect 328730 454764 328736 454776
rect 3568 454736 328736 454764
rect 3568 454724 3574 454736
rect 328730 454724 328736 454736
rect 328788 454724 328794 454776
rect 329834 454724 329840 454776
rect 329892 454764 329898 454776
rect 359550 454764 359556 454776
rect 329892 454736 359556 454764
rect 329892 454724 329898 454736
rect 359550 454724 359556 454736
rect 359608 454724 359614 454776
rect 5074 454656 5080 454708
rect 5132 454696 5138 454708
rect 354766 454696 354772 454708
rect 5132 454668 354772 454696
rect 5132 454656 5138 454668
rect 354766 454656 354772 454668
rect 354824 454656 354830 454708
rect 323394 453636 323400 453688
rect 323452 453676 323458 453688
rect 358262 453676 358268 453688
rect 323452 453648 358268 453676
rect 323452 453636 323458 453648
rect 358262 453636 358268 453648
rect 358320 453636 358326 453688
rect 321002 453568 321008 453620
rect 321060 453608 321066 453620
rect 358354 453608 358360 453620
rect 321060 453580 358360 453608
rect 321060 453568 321066 453580
rect 358354 453568 358360 453580
rect 358412 453568 358418 453620
rect 310882 453500 310888 453552
rect 310940 453540 310946 453552
rect 360838 453540 360844 453552
rect 310940 453512 360844 453540
rect 310940 453500 310946 453512
rect 360838 453500 360844 453512
rect 360896 453500 360902 453552
rect 203518 453432 203524 453484
rect 203576 453472 203582 453484
rect 353754 453472 353760 453484
rect 203576 453444 353760 453472
rect 203576 453432 203582 453444
rect 353754 453432 353760 453444
rect 353812 453432 353818 453484
rect 178678 453364 178684 453416
rect 178736 453404 178742 453416
rect 353386 453404 353392 453416
rect 178736 453376 353392 453404
rect 178736 453364 178742 453376
rect 353386 453364 353392 453376
rect 353444 453364 353450 453416
rect 6914 453296 6920 453348
rect 6972 453336 6978 453348
rect 351362 453336 351368 453348
rect 6972 453308 351368 453336
rect 6972 453296 6978 453308
rect 351362 453296 351368 453308
rect 351420 453296 351426 453348
rect 303890 452208 303896 452260
rect 303948 452248 303954 452260
rect 358078 452248 358084 452260
rect 303948 452220 358084 452248
rect 303948 452208 303954 452220
rect 358078 452208 358084 452220
rect 358136 452208 358142 452260
rect 308490 452140 308496 452192
rect 308548 452180 308554 452192
rect 429194 452180 429200 452192
rect 308548 452152 429200 452180
rect 308548 452140 308554 452152
rect 429194 452140 429200 452152
rect 429252 452140 429258 452192
rect 306374 452072 306380 452124
rect 306432 452112 306438 452124
rect 494054 452112 494060 452124
rect 306432 452084 494060 452112
rect 306432 452072 306438 452084
rect 494054 452072 494060 452084
rect 494112 452072 494118 452124
rect 71774 452004 71780 452056
rect 71832 452044 71838 452056
rect 349246 452044 349252 452056
rect 71832 452016 349252 452044
rect 71832 452004 71838 452016
rect 349246 452004 349252 452016
rect 349304 452004 349310 452056
rect 8938 451936 8944 451988
rect 8996 451976 9002 451988
rect 331858 451976 331864 451988
rect 8996 451948 331864 451976
rect 8996 451936 9002 451948
rect 331858 451936 331864 451948
rect 331916 451936 331922 451988
rect 4982 451868 4988 451920
rect 5040 451908 5046 451920
rect 329926 451908 329932 451920
rect 5040 451880 329932 451908
rect 5040 451868 5046 451880
rect 329926 451868 329932 451880
rect 329984 451868 329990 451920
rect 301958 450780 301964 450832
rect 302016 450820 302022 450832
rect 358170 450820 358176 450832
rect 302016 450792 358176 450820
rect 302016 450780 302022 450792
rect 358170 450780 358176 450792
rect 358228 450780 358234 450832
rect 299658 450712 299664 450764
rect 299716 450752 299722 450764
rect 359642 450752 359648 450764
rect 299716 450724 359648 450752
rect 299716 450712 299722 450724
rect 359642 450712 359648 450724
rect 359700 450712 359706 450764
rect 217686 450644 217692 450696
rect 217744 450684 217750 450696
rect 234246 450684 234252 450696
rect 217744 450656 234252 450684
rect 217744 450644 217750 450656
rect 234246 450644 234252 450656
rect 234304 450644 234310 450696
rect 297266 450644 297272 450696
rect 297324 450684 297330 450696
rect 371878 450684 371884 450696
rect 297324 450656 371884 450684
rect 297324 450644 297330 450656
rect 371878 450644 371884 450656
rect 371936 450644 371942 450696
rect 4798 450576 4804 450628
rect 4856 450616 4862 450628
rect 325326 450616 325332 450628
rect 4856 450588 325332 450616
rect 4856 450576 4862 450588
rect 325326 450576 325332 450588
rect 325384 450576 325390 450628
rect 4890 450508 4896 450560
rect 4948 450548 4954 450560
rect 327626 450548 327632 450560
rect 4948 450520 327632 450548
rect 4948 450508 4954 450520
rect 327626 450508 327632 450520
rect 327684 450508 327690 450560
rect 335446 450508 335452 450560
rect 335504 450548 335510 450560
rect 462314 450548 462320 450560
rect 335504 450520 462320 450548
rect 335504 450508 335510 450520
rect 462314 450508 462320 450520
rect 462372 450508 462378 450560
rect 310514 449488 310520 449540
rect 310572 449528 310578 449540
rect 412634 449528 412640 449540
rect 310572 449500 412640 449528
rect 310572 449488 310578 449500
rect 412634 449488 412640 449500
rect 412692 449488 412698 449540
rect 153194 449420 153200 449472
rect 153252 449460 153258 449472
rect 319898 449460 319904 449472
rect 153252 449432 319904 449460
rect 153252 449420 153258 449432
rect 319898 449420 319904 449432
rect 319956 449420 319962 449472
rect 308214 449352 308220 449404
rect 308272 449392 308278 449404
rect 477494 449392 477500 449404
rect 308272 449364 477500 449392
rect 308272 449352 308278 449364
rect 477494 449352 477500 449364
rect 477552 449352 477558 449404
rect 88334 449284 88340 449336
rect 88392 449324 88398 449336
rect 322198 449324 322204 449336
rect 88392 449296 322204 449324
rect 88392 449284 88398 449296
rect 322198 449284 322204 449296
rect 322256 449284 322262 449336
rect 305822 449216 305828 449268
rect 305880 449256 305886 449268
rect 542354 449256 542360 449268
rect 305880 449228 542360 449256
rect 305880 449216 305886 449228
rect 542354 449216 542360 449228
rect 542412 449216 542418 449268
rect 23474 449148 23480 449200
rect 23532 449188 23538 449200
rect 324498 449188 324504 449200
rect 23532 449160 324504 449188
rect 23532 449148 23538 449160
rect 324498 449148 324504 449160
rect 324556 449148 324562 449200
rect 201494 448128 201500 448180
rect 201552 448168 201558 448180
rect 344738 448168 344744 448180
rect 201552 448140 344744 448168
rect 201552 448128 201558 448140
rect 344738 448128 344744 448140
rect 344796 448128 344802 448180
rect 169754 448060 169760 448112
rect 169812 448100 169818 448112
rect 318334 448100 318340 448112
rect 169812 448072 318340 448100
rect 169812 448060 169818 448072
rect 318334 448060 318340 448072
rect 318392 448060 318398 448112
rect 136634 447992 136640 448044
rect 136692 448032 136698 448044
rect 347038 448032 347044 448044
rect 136692 448004 347044 448032
rect 136692 447992 136698 448004
rect 347038 447992 347044 448004
rect 347096 447992 347102 448044
rect 104894 447924 104900 447976
rect 104952 447964 104958 447976
rect 320634 447964 320640 447976
rect 104952 447936 320640 447964
rect 104952 447924 104958 447936
rect 320634 447924 320640 447936
rect 320692 447924 320698 447976
rect 333054 447924 333060 447976
rect 333112 447964 333118 447976
rect 527174 447964 527180 447976
rect 333112 447936 527180 447964
rect 333112 447924 333118 447936
rect 527174 447924 527180 447936
rect 527232 447924 527238 447976
rect 40034 447856 40040 447908
rect 40092 447896 40098 447908
rect 322934 447896 322940 447908
rect 40092 447868 322940 447896
rect 40092 447856 40098 447868
rect 322934 447856 322940 447868
rect 322992 447856 322998 447908
rect 328454 447856 328460 447908
rect 328512 447896 328518 447908
rect 580350 447896 580356 447908
rect 328512 447868 580356 447896
rect 328512 447856 328518 447868
rect 580350 447856 580356 447868
rect 580408 447856 580414 447908
rect 2866 447788 2872 447840
rect 2924 447828 2930 447840
rect 356422 447828 356428 447840
rect 2924 447800 356428 447828
rect 2924 447788 2930 447800
rect 356422 447788 356428 447800
rect 356480 447788 356486 447840
rect 244274 447244 244280 447296
rect 244332 447284 244338 447296
rect 244918 447284 244924 447296
rect 244332 447256 244924 447284
rect 244332 447244 244338 447256
rect 244918 447244 244924 447256
rect 244976 447244 244982 447296
rect 249794 447244 249800 447296
rect 249852 447284 249858 447296
rect 250254 447284 250260 447296
rect 249852 447256 250260 447284
rect 249852 447244 249858 447256
rect 250254 447244 250260 447256
rect 250312 447244 250318 447296
rect 283006 447244 283012 447296
rect 283064 447284 283070 447296
rect 283742 447284 283748 447296
rect 283064 447256 283748 447284
rect 283064 447244 283070 447256
rect 283742 447244 283748 447256
rect 283800 447244 283806 447296
rect 325694 447244 325700 447296
rect 325752 447284 325758 447296
rect 326614 447284 326620 447296
rect 325752 447256 326620 447284
rect 325752 447244 325758 447256
rect 326614 447244 326620 447256
rect 326672 447244 326678 447296
rect 329834 447244 329840 447296
rect 329892 447284 329898 447296
rect 330478 447284 330484 447296
rect 329892 447256 330484 447284
rect 329892 447244 329898 447256
rect 330478 447244 330484 447256
rect 330536 447244 330542 447296
rect 354674 447244 354680 447296
rect 354732 447284 354738 447296
rect 355318 447284 355324 447296
rect 354732 447256 355324 447284
rect 354732 447244 354738 447256
rect 355318 447244 355324 447256
rect 355376 447244 355382 447296
rect 245010 447040 245016 447092
rect 245068 447080 245074 447092
rect 246758 447080 246764 447092
rect 245068 447052 246764 447080
rect 245068 447040 245074 447052
rect 246758 447040 246764 447052
rect 246816 447040 246822 447092
rect 252462 447040 252468 447092
rect 252520 447080 252526 447092
rect 255314 447080 255320 447092
rect 252520 447052 255320 447080
rect 252520 447040 252526 447052
rect 255314 447040 255320 447052
rect 255372 447040 255378 447092
rect 262858 447040 262864 447092
rect 262916 447080 262922 447092
rect 270034 447080 270040 447092
rect 262916 447052 270040 447080
rect 262916 447040 262922 447052
rect 270034 447040 270040 447052
rect 270092 447040 270098 447092
rect 253842 446972 253848 447024
rect 253900 447012 253906 447024
rect 259178 447012 259184 447024
rect 253900 446984 259184 447012
rect 253900 446972 253906 446984
rect 259178 446972 259184 446984
rect 259236 446972 259242 447024
rect 259362 446972 259368 447024
rect 259420 447012 259426 447024
rect 265434 447012 265440 447024
rect 259420 446984 265440 447012
rect 259420 446972 259426 446984
rect 265434 446972 265440 446984
rect 265492 446972 265498 447024
rect 268470 447012 268476 447024
rect 267706 446984 268476 447012
rect 255222 446904 255228 446956
rect 255280 446944 255286 446956
rect 260374 446944 260380 446956
rect 255280 446916 260380 446944
rect 255280 446904 255286 446916
rect 260374 446904 260380 446916
rect 260432 446904 260438 446956
rect 261478 446904 261484 446956
rect 261536 446944 261542 446956
rect 267706 446944 267734 446984
rect 268470 446972 268476 446984
rect 268528 446972 268534 447024
rect 261536 446916 267734 446944
rect 261536 446904 261542 446916
rect 217962 446836 217968 446888
rect 218020 446876 218026 446888
rect 315942 446876 315948 446888
rect 218020 446848 315948 446876
rect 218020 446836 218026 446848
rect 315942 446836 315948 446848
rect 316000 446836 316006 446888
rect 210418 446768 210424 446820
rect 210476 446808 210482 446820
rect 345934 446808 345940 446820
rect 210476 446780 345940 446808
rect 210476 446768 210482 446780
rect 345934 446768 345940 446780
rect 345992 446768 345998 446820
rect 266998 446632 267004 446684
rect 267056 446672 267062 446684
rect 271598 446672 271604 446684
rect 267056 446644 271604 446672
rect 267056 446632 267062 446644
rect 271598 446632 271604 446644
rect 271656 446632 271662 446684
rect 282178 446632 282184 446684
rect 282236 446672 282242 446684
rect 293402 446672 293408 446684
rect 282236 446644 293408 446672
rect 282236 446632 282242 446644
rect 293402 446632 293408 446644
rect 293460 446632 293466 446684
rect 340046 446632 340052 446684
rect 340104 446672 340110 446684
rect 358998 446672 359004 446684
rect 340104 446644 359004 446672
rect 340104 446632 340110 446644
rect 358998 446632 359004 446644
rect 359056 446632 359062 446684
rect 256602 446564 256608 446616
rect 256660 446604 256666 446616
rect 262306 446604 262312 446616
rect 256660 446576 262312 446604
rect 256660 446564 256666 446576
rect 262306 446564 262312 446576
rect 262364 446564 262370 446616
rect 276658 446564 276664 446616
rect 276716 446604 276722 446616
rect 288710 446604 288716 446616
rect 276716 446576 288716 446604
rect 276716 446564 276722 446576
rect 288710 446564 288716 446576
rect 288768 446564 288774 446616
rect 307386 446564 307392 446616
rect 307444 446604 307450 446616
rect 340874 446604 340880 446616
rect 307444 446576 340880 446604
rect 307444 446564 307450 446576
rect 340874 446564 340880 446576
rect 340932 446564 340938 446616
rect 342438 446564 342444 446616
rect 342496 446604 342502 446616
rect 357434 446604 357440 446616
rect 342496 446576 357440 446604
rect 342496 446564 342502 446576
rect 357434 446564 357440 446576
rect 357492 446564 357498 446616
rect 220078 446496 220084 446548
rect 220136 446536 220142 446548
rect 232774 446536 232780 446548
rect 220136 446508 232780 446536
rect 220136 446496 220142 446508
rect 232774 446496 232780 446508
rect 232832 446496 232838 446548
rect 260742 446496 260748 446548
rect 260800 446536 260806 446548
rect 266998 446536 267004 446548
rect 260800 446508 267004 446536
rect 260800 446496 260806 446508
rect 266998 446496 267004 446508
rect 267056 446496 267062 446548
rect 275278 446496 275284 446548
rect 275336 446536 275342 446548
rect 287146 446536 287152 446548
rect 275336 446508 287152 446536
rect 275336 446496 275342 446508
rect 287146 446496 287152 446508
rect 287204 446496 287210 446548
rect 315206 446496 315212 446548
rect 315264 446536 315270 446548
rect 358814 446536 358820 446548
rect 315264 446508 358820 446536
rect 315264 446496 315270 446508
rect 358814 446496 358820 446508
rect 358872 446496 358878 446548
rect 217778 446428 217784 446480
rect 217836 446468 217842 446480
rect 233510 446468 233516 446480
rect 217836 446440 233516 446468
rect 217836 446428 217842 446440
rect 233510 446428 233516 446440
rect 233568 446428 233574 446480
rect 257982 446428 257988 446480
rect 258040 446468 258046 446480
rect 263870 446468 263876 446480
rect 258040 446440 263876 446468
rect 258040 446428 258046 446440
rect 263870 446428 263876 446440
rect 263928 446428 263934 446480
rect 264882 446428 264888 446480
rect 264940 446468 264946 446480
rect 273162 446468 273168 446480
rect 264940 446440 273168 446468
rect 264940 446428 264946 446440
rect 273162 446428 273168 446440
rect 273220 446428 273226 446480
rect 278038 446428 278044 446480
rect 278096 446468 278102 446480
rect 290274 446468 290280 446480
rect 278096 446440 290280 446468
rect 278096 446428 278102 446440
rect 290274 446428 290280 446440
rect 290332 446428 290338 446480
rect 313642 446428 313648 446480
rect 313700 446468 313706 446480
rect 357526 446468 357532 446480
rect 313700 446440 357532 446468
rect 313700 446428 313706 446440
rect 357526 446428 357532 446440
rect 357584 446428 357590 446480
rect 256694 446360 256700 446412
rect 256752 446400 256758 446412
rect 257246 446400 257252 446412
rect 256752 446372 257252 446400
rect 256752 446360 256758 446372
rect 257246 446360 257252 446372
rect 257304 446360 257310 446412
rect 309778 446360 309784 446412
rect 309836 446400 309842 446412
rect 346302 446400 346308 446412
rect 309836 446372 346308 446400
rect 309836 446360 309842 446372
rect 346302 446360 346308 446372
rect 346360 446360 346366 446412
rect 318702 446292 318708 446344
rect 318760 446332 318766 446344
rect 357986 446332 357992 446344
rect 318760 446304 357992 446332
rect 318760 446292 318766 446304
rect 357986 446292 357992 446304
rect 358044 446292 358050 446344
rect 314378 446224 314384 446276
rect 314436 446264 314442 446276
rect 364978 446264 364984 446276
rect 314436 446236 364984 446264
rect 314436 446224 314442 446236
rect 364978 446224 364984 446236
rect 365036 446224 365042 446276
rect 288342 446156 288348 446208
rect 288400 446196 288406 446208
rect 359550 446196 359556 446208
rect 288400 446168 359556 446196
rect 288400 446156 288406 446168
rect 359550 446156 359556 446168
rect 359608 446156 359614 446208
rect 232314 446088 232320 446140
rect 232372 446128 232378 446140
rect 338482 446128 338488 446140
rect 232372 446100 338488 446128
rect 232372 446088 232378 446100
rect 338482 446088 338488 446100
rect 338540 446088 338546 446140
rect 233786 446020 233792 446072
rect 233844 446060 233850 446072
rect 343174 446060 343180 446072
rect 233844 446032 343180 446060
rect 233844 446020 233850 446032
rect 343174 446020 343180 446032
rect 343232 446020 343238 446072
rect 343266 446020 343272 446072
rect 343324 446060 343330 446072
rect 357158 446060 357164 446072
rect 343324 446032 357164 446060
rect 343324 446020 343330 446032
rect 357158 446020 357164 446032
rect 357216 446020 357222 446072
rect 231118 445952 231124 446004
rect 231176 445992 231182 446004
rect 347866 445992 347872 446004
rect 231176 445964 347872 445992
rect 231176 445952 231182 445964
rect 347866 445952 347872 445964
rect 347924 445952 347930 446004
rect 232222 445884 232228 445936
rect 232280 445924 232286 445936
rect 352558 445924 352564 445936
rect 232280 445896 352564 445924
rect 232280 445884 232286 445896
rect 352558 445884 352564 445896
rect 352616 445884 352622 445936
rect 233878 445816 233884 445868
rect 233936 445856 233942 445868
rect 360286 445856 360292 445868
rect 233936 445828 360292 445856
rect 233936 445816 233942 445828
rect 360286 445816 360292 445828
rect 360344 445816 360350 445868
rect 305086 445748 305092 445800
rect 305144 445788 305150 445800
rect 338758 445788 338764 445800
rect 305144 445760 338764 445788
rect 305144 445748 305150 445760
rect 338758 445748 338764 445760
rect 338816 445748 338822 445800
rect 351914 445748 351920 445800
rect 351972 445788 351978 445800
rect 358722 445788 358728 445800
rect 351972 445760 358728 445788
rect 351972 445748 351978 445760
rect 358722 445748 358728 445760
rect 358780 445748 358786 445800
rect 4890 445136 4896 445188
rect 4948 445176 4954 445188
rect 345566 445176 345572 445188
rect 4948 445148 345572 445176
rect 4948 445136 4954 445148
rect 345566 445136 345572 445148
rect 345624 445136 345630 445188
rect 346302 445136 346308 445188
rect 346360 445176 346366 445188
rect 580626 445176 580632 445188
rect 346360 445148 580632 445176
rect 346360 445136 346366 445148
rect 580626 445136 580632 445148
rect 580684 445136 580690 445188
rect 40678 445068 40684 445120
rect 40736 445108 40742 445120
rect 337010 445108 337016 445120
rect 40736 445080 337016 445108
rect 40736 445068 40742 445080
rect 337010 445068 337016 445080
rect 337068 445068 337074 445120
rect 340874 445068 340880 445120
rect 340932 445108 340938 445120
rect 580534 445108 580540 445120
rect 340932 445080 580540 445108
rect 340932 445068 340938 445080
rect 580534 445068 580540 445080
rect 580592 445068 580598 445120
rect 3878 445000 3884 445052
rect 3936 445040 3942 445052
rect 318702 445040 318708 445052
rect 3936 445012 318708 445040
rect 3936 445000 3942 445012
rect 318702 445000 318708 445012
rect 318760 445000 318766 445052
rect 338758 445000 338764 445052
rect 338816 445040 338822 445052
rect 580442 445040 580448 445052
rect 338816 445012 580448 445040
rect 338816 445000 338822 445012
rect 580442 445000 580448 445012
rect 580500 445000 580506 445052
rect 312078 444932 312084 444984
rect 312136 444972 312142 444984
rect 367738 444972 367744 444984
rect 312136 444944 367744 444972
rect 312136 444932 312142 444944
rect 367738 444932 367744 444944
rect 367796 444932 367802 444984
rect 231210 444864 231216 444916
rect 231268 444904 231274 444916
rect 340874 444904 340880 444916
rect 231268 444876 340880 444904
rect 231268 444864 231274 444876
rect 340874 444864 340880 444876
rect 340932 444864 340938 444916
rect 228358 444796 228364 444848
rect 228416 444836 228422 444848
rect 344002 444836 344008 444848
rect 228416 444808 344008 444836
rect 228416 444796 228422 444808
rect 344002 444796 344008 444808
rect 344060 444796 344066 444848
rect 218422 444728 218428 444780
rect 218480 444768 218486 444780
rect 348602 444768 348608 444780
rect 218480 444740 348608 444768
rect 218480 444728 218486 444740
rect 348602 444728 348608 444740
rect 348660 444728 348666 444780
rect 174538 444660 174544 444712
rect 174596 444700 174602 444712
rect 341610 444700 341616 444712
rect 174596 444672 341616 444700
rect 174596 444660 174602 444672
rect 341610 444660 341616 444672
rect 341668 444660 341674 444712
rect 106918 444592 106924 444644
rect 106976 444632 106982 444644
rect 339310 444632 339316 444644
rect 106976 444604 339316 444632
rect 106976 444592 106982 444604
rect 339310 444592 339316 444604
rect 339368 444592 339374 444644
rect 316770 444524 316776 444576
rect 316828 444564 316834 444576
rect 365070 444564 365076 444576
rect 316828 444536 365076 444564
rect 316828 444524 316834 444536
rect 365070 444524 365076 444536
rect 365128 444524 365134 444576
rect 43438 444456 43444 444508
rect 43496 444496 43502 444508
rect 350166 444496 350172 444508
rect 43496 444468 350172 444496
rect 43496 444456 43502 444468
rect 350166 444456 350172 444468
rect 350224 444456 350230 444508
rect 319070 444388 319076 444440
rect 319128 444428 319134 444440
rect 365162 444428 365168 444440
rect 319128 444400 365168 444428
rect 319128 444388 319134 444400
rect 365162 444388 365168 444400
rect 365220 444388 365226 444440
rect 288342 444088 288348 444100
rect 277366 444060 288348 444088
rect 3786 443912 3792 443964
rect 3844 443952 3850 443964
rect 233786 443952 233792 443964
rect 3844 443924 233792 443952
rect 3844 443912 3850 443924
rect 233786 443912 233792 443924
rect 233844 443912 233850 443964
rect 3510 443844 3516 443896
rect 3568 443884 3574 443896
rect 233878 443884 233884 443896
rect 3568 443856 233884 443884
rect 3568 443844 3574 443856
rect 233878 443844 233884 443856
rect 233936 443844 233942 443896
rect 3602 443776 3608 443828
rect 3660 443816 3666 443828
rect 277366 443816 277394 444060
rect 288342 444048 288348 444060
rect 288400 444048 288406 444100
rect 3660 443788 277394 443816
rect 3660 443776 3666 443788
rect 3970 443708 3976 443760
rect 4028 443748 4034 443760
rect 343266 443748 343272 443760
rect 4028 443720 343272 443748
rect 4028 443708 4034 443720
rect 343266 443708 343272 443720
rect 343324 443708 343330 443760
rect 3694 443640 3700 443692
rect 3752 443680 3758 443692
rect 351914 443680 351920 443692
rect 3752 443652 351920 443680
rect 3752 443640 3758 443652
rect 351914 443640 351920 443652
rect 351972 443640 351978 443692
rect 320818 443572 320824 443624
rect 320876 443612 320882 443624
rect 320876 443584 325694 443612
rect 320876 443572 320882 443584
rect 298066 443516 303016 443544
rect 298066 443204 298094 443516
rect 298186 443436 298192 443488
rect 298244 443436 298250 443488
rect 296686 443176 298094 443204
rect 180058 443096 180064 443148
rect 180116 443136 180122 443148
rect 296686 443136 296714 443176
rect 180116 443108 296714 443136
rect 180116 443096 180122 443108
rect 298204 443068 298232 443436
rect 302988 443272 303016 443516
rect 316006 443516 322336 443544
rect 303154 443436 303160 443488
rect 303212 443436 303218 443488
rect 303172 443340 303200 443436
rect 316006 443340 316034 443516
rect 320818 443436 320824 443488
rect 320876 443436 320882 443488
rect 303172 443312 316034 443340
rect 302988 443244 307754 443272
rect 307726 443068 307754 443244
rect 320836 443136 320864 443436
rect 322308 443204 322336 443516
rect 325666 443476 325694 443584
rect 360838 443476 360844 443488
rect 325666 443448 327074 443476
rect 327046 443408 327074 443448
rect 354646 443448 360844 443476
rect 327046 443380 329834 443408
rect 329806 443340 329834 443380
rect 329806 443312 331168 443340
rect 328426 443244 329834 443272
rect 328426 443204 328454 443244
rect 322308 443176 328454 443204
rect 311820 443108 320864 443136
rect 311820 443068 311848 443108
rect 298204 443040 303200 443068
rect 307726 443040 311848 443068
rect 312004 443040 317276 443068
rect 303172 442994 303200 443040
rect 312004 443000 312032 443040
rect 303080 442966 303200 442994
rect 309106 442972 312032 443000
rect 317248 443000 317276 443040
rect 317248 442972 321554 443000
rect 303080 442932 303108 442966
rect 309106 442932 309134 442972
rect 303080 442904 309134 442932
rect 321526 442796 321554 442972
rect 329806 442932 329834 443244
rect 331140 443136 331168 443312
rect 332566 443176 335354 443204
rect 332566 443136 332594 443176
rect 331140 443108 332594 443136
rect 335326 443136 335354 443176
rect 354646 443136 354674 443448
rect 360838 443436 360844 443448
rect 360896 443436 360902 443488
rect 335326 443108 354674 443136
rect 580350 443068 580356 443080
rect 330956 443040 580356 443068
rect 330956 442932 330984 443040
rect 580350 443028 580356 443040
rect 580408 443028 580414 443080
rect 580258 443000 580264 443012
rect 329806 442904 330984 442932
rect 331186 442972 580264 443000
rect 331186 442796 331214 442972
rect 580258 442960 580264 442972
rect 580316 442960 580322 443012
rect 321526 442768 331214 442796
rect 3418 433984 3424 434036
rect 3476 434024 3482 434036
rect 232222 434024 232228 434036
rect 3476 433996 232228 434024
rect 3476 433984 3482 433996
rect 232222 433984 232228 433996
rect 232280 433984 232286 434036
rect 365162 431876 365168 431928
rect 365220 431916 365226 431928
rect 580166 431916 580172 431928
rect 365220 431888 580172 431916
rect 365220 431876 365226 431888
rect 580166 431876 580172 431888
rect 580224 431876 580230 431928
rect 3326 423580 3332 423632
rect 3384 423620 3390 423632
rect 40678 423620 40684 423632
rect 3384 423592 40684 423620
rect 3384 423580 3390 423592
rect 40678 423580 40684 423592
rect 40736 423580 40742 423632
rect 3326 411204 3332 411256
rect 3384 411244 3390 411256
rect 232222 411244 232228 411256
rect 3384 411216 232228 411244
rect 3384 411204 3390 411216
rect 232222 411204 232228 411216
rect 232280 411204 232286 411256
rect 365070 379448 365076 379500
rect 365128 379488 365134 379500
rect 579614 379488 579620 379500
rect 365128 379460 579620 379488
rect 365128 379448 365134 379460
rect 579614 379448 579620 379460
rect 579672 379448 579678 379500
rect 3326 372512 3332 372564
rect 3384 372552 3390 372564
rect 106918 372552 106924 372564
rect 3384 372524 106924 372552
rect 3384 372512 3390 372524
rect 106918 372512 106924 372524
rect 106976 372512 106982 372564
rect 3326 358708 3332 358760
rect 3384 358748 3390 358760
rect 231210 358748 231216 358760
rect 3384 358720 231216 358748
rect 3384 358708 3390 358720
rect 231210 358708 231216 358720
rect 231268 358708 231274 358760
rect 364978 325592 364984 325644
rect 365036 325632 365042 325644
rect 579982 325632 579988 325644
rect 365036 325604 579988 325632
rect 365036 325592 365042 325604
rect 579982 325592 579988 325604
rect 580040 325592 580046 325644
rect 3326 320084 3332 320136
rect 3384 320124 3390 320136
rect 174538 320124 174544 320136
rect 3384 320096 174544 320124
rect 3384 320084 3390 320096
rect 174538 320084 174544 320096
rect 174596 320084 174602 320136
rect 304994 310496 305000 310548
rect 305052 310536 305058 310548
rect 305178 310536 305184 310548
rect 305052 310508 305184 310536
rect 305052 310496 305058 310508
rect 305178 310496 305184 310508
rect 305236 310496 305242 310548
rect 309410 310496 309416 310548
rect 309468 310536 309474 310548
rect 309778 310536 309784 310548
rect 309468 310508 309784 310536
rect 309468 310496 309474 310508
rect 309778 310496 309784 310508
rect 309836 310496 309842 310548
rect 310790 310496 310796 310548
rect 310848 310536 310854 310548
rect 311158 310536 311164 310548
rect 310848 310508 311164 310536
rect 310848 310496 310854 310508
rect 311158 310496 311164 310508
rect 311216 310496 311222 310548
rect 312170 310496 312176 310548
rect 312228 310536 312234 310548
rect 312538 310536 312544 310548
rect 312228 310508 312544 310536
rect 312228 310496 312234 310508
rect 312538 310496 312544 310508
rect 312596 310496 312602 310548
rect 215202 309068 215208 309120
rect 215260 309108 215266 309120
rect 279694 309108 279700 309120
rect 215260 309080 279700 309108
rect 215260 309068 215266 309080
rect 279694 309068 279700 309080
rect 279752 309068 279758 309120
rect 323762 309068 323768 309120
rect 323820 309108 323826 309120
rect 358998 309108 359004 309120
rect 323820 309080 359004 309108
rect 323820 309068 323826 309080
rect 358998 309068 359004 309080
rect 359056 309068 359062 309120
rect 216490 309000 216496 309052
rect 216548 309040 216554 309052
rect 280430 309040 280436 309052
rect 216548 309012 280436 309040
rect 216548 309000 216554 309012
rect 280430 309000 280436 309012
rect 280488 309000 280494 309052
rect 324498 309000 324504 309052
rect 324556 309040 324562 309052
rect 361482 309040 361488 309052
rect 324556 309012 361488 309040
rect 324556 309000 324562 309012
rect 361482 309000 361488 309012
rect 361540 309000 361546 309052
rect 189718 308932 189724 308984
rect 189776 308972 189782 308984
rect 255958 308972 255964 308984
rect 189776 308944 255964 308972
rect 189776 308932 189782 308944
rect 255958 308932 255964 308944
rect 256016 308932 256022 308984
rect 316402 308932 316408 308984
rect 316460 308972 316466 308984
rect 326338 308972 326344 308984
rect 316460 308944 326344 308972
rect 316460 308932 316466 308944
rect 326338 308932 326344 308944
rect 326396 308932 326402 308984
rect 331122 308932 331128 308984
rect 331180 308972 331186 308984
rect 331490 308972 331496 308984
rect 331180 308944 331496 308972
rect 331180 308932 331186 308944
rect 331490 308932 331496 308944
rect 331548 308932 331554 308984
rect 354214 308932 354220 308984
rect 354272 308972 354278 308984
rect 367278 308972 367284 308984
rect 354272 308944 367284 308972
rect 354272 308932 354278 308944
rect 367278 308932 367284 308944
rect 367336 308932 367342 308984
rect 182818 308864 182824 308916
rect 182876 308904 182882 308916
rect 254578 308904 254584 308916
rect 182876 308876 254584 308904
rect 182876 308864 182882 308876
rect 254578 308864 254584 308876
rect 254636 308864 254642 308916
rect 294966 308864 294972 308916
rect 295024 308904 295030 308916
rect 356882 308904 356888 308916
rect 295024 308876 356888 308904
rect 295024 308864 295030 308876
rect 356882 308864 356888 308876
rect 356940 308864 356946 308916
rect 356974 308864 356980 308916
rect 357032 308904 357038 308916
rect 369118 308904 369124 308916
rect 357032 308876 369124 308904
rect 357032 308864 357038 308876
rect 369118 308864 369124 308876
rect 369176 308864 369182 308916
rect 213822 308796 213828 308848
rect 213880 308836 213886 308848
rect 287330 308836 287336 308848
rect 213880 308808 287336 308836
rect 213880 308796 213886 308808
rect 287330 308796 287336 308808
rect 287388 308796 287394 308848
rect 294230 308796 294236 308848
rect 294288 308836 294294 308848
rect 356146 308836 356152 308848
rect 294288 308808 356152 308836
rect 294288 308796 294294 308808
rect 356146 308796 356152 308808
rect 356204 308796 356210 308848
rect 178678 308728 178684 308780
rect 178736 308768 178742 308780
rect 253198 308768 253204 308780
rect 178736 308740 253204 308768
rect 178736 308728 178742 308740
rect 253198 308728 253204 308740
rect 253256 308728 253262 308780
rect 294506 308728 294512 308780
rect 294564 308768 294570 308780
rect 357066 308768 357072 308780
rect 294564 308740 357072 308768
rect 294564 308728 294570 308740
rect 357066 308728 357072 308740
rect 357124 308728 357130 308780
rect 68278 308660 68284 308712
rect 68336 308700 68342 308712
rect 236362 308700 236368 308712
rect 68336 308672 236368 308700
rect 68336 308660 68342 308672
rect 236362 308660 236368 308672
rect 236420 308660 236426 308712
rect 266630 308700 266636 308712
rect 253906 308672 266636 308700
rect 50338 308592 50344 308644
rect 50396 308632 50402 308644
rect 240778 308632 240784 308644
rect 50396 308604 240784 308632
rect 50396 308592 50402 308604
rect 240778 308592 240784 308604
rect 240836 308592 240842 308644
rect 253382 308592 253388 308644
rect 253440 308632 253446 308644
rect 253906 308632 253934 308672
rect 266630 308660 266636 308672
rect 266688 308660 266694 308712
rect 291286 308660 291292 308712
rect 291344 308700 291350 308712
rect 355318 308700 355324 308712
rect 291344 308672 355324 308700
rect 291344 308660 291350 308672
rect 355318 308660 355324 308672
rect 355376 308660 355382 308712
rect 356514 308660 356520 308712
rect 356572 308700 356578 308712
rect 356572 308672 369854 308700
rect 356572 308660 356578 308672
rect 253440 308604 253934 308632
rect 253440 308592 253446 308604
rect 292666 308592 292672 308644
rect 292724 308632 292730 308644
rect 357250 308632 357256 308644
rect 292724 308604 357256 308632
rect 292724 308592 292730 308604
rect 357250 308592 357256 308604
rect 357308 308592 357314 308644
rect 46198 308524 46204 308576
rect 46256 308564 46262 308576
rect 239398 308564 239404 308576
rect 46256 308536 239404 308564
rect 46256 308524 46262 308536
rect 239398 308524 239404 308536
rect 239456 308524 239462 308576
rect 248598 308524 248604 308576
rect 248656 308564 248662 308576
rect 249150 308564 249156 308576
rect 248656 308536 249156 308564
rect 248656 308524 248662 308536
rect 249150 308524 249156 308536
rect 249208 308524 249214 308576
rect 290550 308524 290556 308576
rect 290608 308564 290614 308576
rect 355410 308564 355416 308576
rect 290608 308536 355416 308564
rect 290608 308524 290614 308536
rect 355410 308524 355416 308536
rect 355468 308524 355474 308576
rect 358354 308524 358360 308576
rect 358412 308564 358418 308576
rect 368842 308564 368848 308576
rect 358412 308536 368848 308564
rect 358412 308524 358418 308536
rect 368842 308524 368848 308536
rect 368900 308524 368906 308576
rect 369826 308564 369854 308672
rect 370130 308564 370136 308576
rect 369826 308536 370136 308564
rect 370130 308524 370136 308536
rect 370188 308524 370194 308576
rect 32398 308456 32404 308508
rect 32456 308496 32462 308508
rect 233050 308496 233056 308508
rect 32456 308468 233056 308496
rect 32456 308456 32462 308468
rect 233050 308456 233056 308468
rect 233108 308456 233114 308508
rect 233326 308456 233332 308508
rect 233384 308496 233390 308508
rect 234154 308496 234160 308508
rect 233384 308468 234160 308496
rect 233384 308456 233390 308468
rect 234154 308456 234160 308468
rect 234212 308456 234218 308508
rect 247218 308456 247224 308508
rect 247276 308496 247282 308508
rect 247954 308496 247960 308508
rect 247276 308468 247960 308496
rect 247276 308456 247282 308468
rect 247954 308456 247960 308468
rect 248012 308456 248018 308508
rect 248414 308456 248420 308508
rect 248472 308496 248478 308508
rect 248782 308496 248788 308508
rect 248472 308468 248788 308496
rect 248472 308456 248478 308468
rect 248782 308456 248788 308468
rect 248840 308456 248846 308508
rect 252738 308456 252744 308508
rect 252796 308496 252802 308508
rect 253014 308496 253020 308508
rect 252796 308468 253020 308496
rect 252796 308456 252802 308468
rect 253014 308456 253020 308468
rect 253072 308456 253078 308508
rect 271874 308456 271880 308508
rect 271932 308496 271938 308508
rect 272150 308496 272156 308508
rect 271932 308468 272156 308496
rect 271932 308456 271938 308468
rect 272150 308456 272156 308468
rect 272208 308456 272214 308508
rect 290826 308456 290832 308508
rect 290884 308496 290890 308508
rect 357158 308496 357164 308508
rect 290884 308468 357164 308496
rect 290884 308456 290890 308468
rect 357158 308456 357164 308468
rect 357216 308456 357222 308508
rect 25498 308388 25504 308440
rect 25556 308428 25562 308440
rect 231762 308428 231768 308440
rect 25556 308400 231768 308428
rect 25556 308388 25562 308400
rect 231762 308388 231768 308400
rect 231820 308388 231826 308440
rect 231946 308388 231952 308440
rect 232004 308428 232010 308440
rect 232774 308428 232780 308440
rect 232004 308400 232780 308428
rect 232004 308388 232010 308400
rect 232774 308388 232780 308400
rect 232832 308388 232838 308440
rect 233234 308388 233240 308440
rect 233292 308428 233298 308440
rect 233694 308428 233700 308440
rect 233292 308400 233700 308428
rect 233292 308388 233298 308400
rect 233694 308388 233700 308400
rect 233752 308388 233758 308440
rect 247126 308388 247132 308440
rect 247184 308428 247190 308440
rect 247862 308428 247868 308440
rect 247184 308400 247868 308428
rect 247184 308388 247190 308400
rect 247862 308388 247868 308400
rect 247920 308388 247926 308440
rect 248690 308388 248696 308440
rect 248748 308428 248754 308440
rect 249518 308428 249524 308440
rect 248748 308400 249524 308428
rect 248748 308388 248754 308400
rect 249518 308388 249524 308400
rect 249576 308388 249582 308440
rect 249886 308388 249892 308440
rect 249944 308428 249950 308440
rect 250530 308428 250536 308440
rect 249944 308400 250536 308428
rect 249944 308388 249950 308400
rect 250530 308388 250536 308400
rect 250588 308388 250594 308440
rect 251542 308388 251548 308440
rect 251600 308428 251606 308440
rect 252278 308428 252284 308440
rect 251600 308400 252284 308428
rect 251600 308388 251606 308400
rect 252278 308388 252284 308400
rect 252336 308388 252342 308440
rect 252646 308388 252652 308440
rect 252704 308428 252710 308440
rect 253290 308428 253296 308440
rect 252704 308400 253296 308428
rect 252704 308388 252710 308400
rect 253290 308388 253296 308400
rect 253348 308388 253354 308440
rect 264974 308388 264980 308440
rect 265032 308428 265038 308440
rect 265342 308428 265348 308440
rect 265032 308400 265348 308428
rect 265032 308388 265038 308400
rect 265342 308388 265348 308400
rect 265400 308388 265406 308440
rect 266446 308388 266452 308440
rect 266504 308428 266510 308440
rect 266814 308428 266820 308440
rect 266504 308400 266820 308428
rect 266504 308388 266510 308400
rect 266814 308388 266820 308400
rect 266872 308388 266878 308440
rect 269206 308388 269212 308440
rect 269264 308428 269270 308440
rect 270034 308428 270040 308440
rect 269264 308400 270040 308428
rect 269264 308388 269270 308400
rect 270034 308388 270040 308400
rect 270092 308388 270098 308440
rect 270678 308388 270684 308440
rect 270736 308428 270742 308440
rect 271506 308428 271512 308440
rect 270736 308400 271512 308428
rect 270736 308388 270742 308400
rect 271506 308388 271512 308400
rect 271564 308388 271570 308440
rect 271966 308388 271972 308440
rect 272024 308428 272030 308440
rect 272794 308428 272800 308440
rect 272024 308400 272800 308428
rect 272024 308388 272030 308400
rect 272794 308388 272800 308400
rect 272852 308388 272858 308440
rect 357802 308428 357808 308440
rect 292546 308400 357808 308428
rect 218974 308320 218980 308372
rect 219032 308360 219038 308372
rect 279050 308360 279056 308372
rect 219032 308332 279056 308360
rect 219032 308320 219038 308332
rect 279050 308320 279056 308332
rect 279108 308320 279114 308372
rect 219066 308252 219072 308304
rect 219124 308292 219130 308304
rect 277670 308292 277676 308304
rect 219124 308264 277676 308292
rect 219124 308252 219130 308264
rect 277670 308252 277676 308264
rect 277728 308252 277734 308304
rect 218882 308184 218888 308236
rect 218940 308224 218946 308236
rect 218940 308196 253934 308224
rect 218940 308184 218946 308196
rect 244366 308116 244372 308168
rect 244424 308156 244430 308168
rect 244734 308156 244740 308168
rect 244424 308128 244740 308156
rect 244424 308116 244430 308128
rect 244734 308116 244740 308128
rect 244792 308116 244798 308168
rect 245930 308116 245936 308168
rect 245988 308156 245994 308168
rect 246574 308156 246580 308168
rect 245988 308128 246580 308156
rect 245988 308116 245994 308128
rect 246574 308116 246580 308128
rect 246632 308116 246638 308168
rect 249978 308116 249984 308168
rect 250036 308156 250042 308168
rect 250254 308156 250260 308168
rect 250036 308128 250260 308156
rect 250036 308116 250042 308128
rect 250254 308116 250260 308128
rect 250312 308116 250318 308168
rect 252830 308116 252836 308168
rect 252888 308156 252894 308168
rect 253658 308156 253664 308168
rect 252888 308128 253664 308156
rect 252888 308116 252894 308128
rect 253658 308116 253664 308128
rect 253716 308116 253722 308168
rect 231762 308048 231768 308100
rect 231820 308088 231826 308100
rect 236178 308088 236184 308100
rect 231820 308060 236184 308088
rect 231820 308048 231826 308060
rect 236178 308048 236184 308060
rect 236236 308048 236242 308100
rect 244550 308048 244556 308100
rect 244608 308088 244614 308100
rect 245194 308088 245200 308100
rect 244608 308060 245200 308088
rect 244608 308048 244614 308060
rect 245194 308048 245200 308060
rect 245252 308048 245258 308100
rect 246022 308048 246028 308100
rect 246080 308088 246086 308100
rect 246942 308088 246948 308100
rect 246080 308060 246948 308088
rect 246080 308048 246086 308060
rect 246942 308048 246948 308060
rect 247000 308048 247006 308100
rect 253906 308088 253934 308196
rect 263502 308184 263508 308236
rect 263560 308224 263566 308236
rect 264054 308224 264060 308236
rect 263560 308196 264060 308224
rect 263560 308184 263566 308196
rect 264054 308184 264060 308196
rect 264112 308184 264118 308236
rect 266538 308184 266544 308236
rect 266596 308224 266602 308236
rect 267366 308224 267372 308236
rect 266596 308196 267372 308224
rect 266596 308184 266602 308196
rect 267366 308184 267372 308196
rect 267424 308184 267430 308236
rect 268010 308184 268016 308236
rect 268068 308224 268074 308236
rect 268746 308224 268752 308236
rect 268068 308196 268752 308224
rect 268068 308184 268074 308196
rect 268746 308184 268752 308196
rect 268804 308184 268810 308236
rect 269298 308184 269304 308236
rect 269356 308224 269362 308236
rect 270126 308224 270132 308236
rect 269356 308196 270132 308224
rect 269356 308184 269362 308196
rect 270126 308184 270132 308196
rect 270184 308184 270190 308236
rect 270494 308184 270500 308236
rect 270552 308224 270558 308236
rect 270954 308224 270960 308236
rect 270552 308196 270960 308224
rect 270552 308184 270558 308196
rect 270954 308184 270960 308196
rect 271012 308184 271018 308236
rect 289906 308184 289912 308236
rect 289964 308224 289970 308236
rect 292546 308224 292574 308400
rect 357802 308388 357808 308400
rect 357860 308388 357866 308440
rect 358814 308388 358820 308440
rect 358872 308428 358878 308440
rect 370498 308428 370504 308440
rect 358872 308400 370504 308428
rect 358872 308388 358878 308400
rect 370498 308388 370504 308400
rect 370556 308388 370562 308440
rect 356146 308320 356152 308372
rect 356204 308360 356210 308372
rect 356974 308360 356980 308372
rect 356204 308332 356980 308360
rect 356204 308320 356210 308332
rect 356974 308320 356980 308332
rect 357032 308320 357038 308372
rect 358262 308320 358268 308372
rect 358320 308360 358326 308372
rect 360010 308360 360016 308372
rect 358320 308332 360016 308360
rect 358320 308320 358326 308332
rect 360010 308320 360016 308332
rect 360068 308320 360074 308372
rect 355594 308252 355600 308304
rect 355652 308292 355658 308304
rect 367922 308292 367928 308304
rect 355652 308264 367928 308292
rect 355652 308252 355658 308264
rect 367922 308252 367928 308264
rect 367980 308252 367986 308304
rect 289964 308196 292574 308224
rect 289964 308184 289970 308196
rect 355134 308184 355140 308236
rect 355192 308224 355198 308236
rect 367554 308224 367560 308236
rect 355192 308196 367560 308224
rect 355192 308184 355198 308196
rect 367554 308184 367560 308196
rect 367612 308184 367618 308236
rect 263686 308116 263692 308168
rect 263744 308156 263750 308168
rect 264330 308156 264336 308168
rect 263744 308128 264336 308156
rect 263744 308116 263750 308128
rect 264330 308116 264336 308128
rect 264388 308116 264394 308168
rect 265250 308116 265256 308168
rect 265308 308156 265314 308168
rect 265986 308156 265992 308168
rect 265308 308128 265992 308156
rect 265308 308116 265314 308128
rect 265986 308116 265992 308128
rect 266044 308116 266050 308168
rect 276290 308156 276296 308168
rect 268212 308128 276296 308156
rect 268212 308088 268240 308128
rect 276290 308116 276296 308128
rect 276348 308116 276354 308168
rect 359642 308116 359648 308168
rect 359700 308156 359706 308168
rect 362310 308156 362316 308168
rect 359700 308128 362316 308156
rect 359700 308116 359706 308128
rect 362310 308116 362316 308128
rect 362368 308116 362374 308168
rect 253906 308060 268240 308088
rect 270494 308048 270500 308100
rect 270552 308088 270558 308100
rect 271414 308088 271420 308100
rect 270552 308060 271420 308088
rect 270552 308048 270558 308060
rect 271414 308048 271420 308060
rect 271472 308048 271478 308100
rect 326338 308048 326344 308100
rect 326396 308088 326402 308100
rect 331766 308088 331772 308100
rect 326396 308060 331772 308088
rect 326396 308048 326402 308060
rect 331766 308048 331772 308060
rect 331824 308048 331830 308100
rect 350994 308048 351000 308100
rect 351052 308088 351058 308100
rect 359458 308088 359464 308100
rect 351052 308060 359464 308088
rect 351052 308048 351058 308060
rect 359458 308048 359464 308060
rect 359516 308048 359522 308100
rect 360194 308048 360200 308100
rect 360252 308088 360258 308100
rect 368750 308088 368756 308100
rect 360252 308060 368756 308088
rect 360252 308048 360258 308060
rect 368750 308048 368756 308060
rect 368808 308048 368814 308100
rect 233050 307980 233056 308032
rect 233108 308020 233114 308032
rect 238018 308020 238024 308032
rect 233108 307992 238024 308020
rect 233108 307980 233114 307992
rect 238018 307980 238024 307992
rect 238076 307980 238082 308032
rect 244366 307980 244372 308032
rect 244424 308020 244430 308032
rect 245102 308020 245108 308032
rect 244424 307992 245108 308020
rect 244424 307980 244430 307992
rect 245102 307980 245108 307992
rect 245160 307980 245166 308032
rect 249978 307980 249984 308032
rect 250036 308020 250042 308032
rect 250898 308020 250904 308032
rect 250036 307992 250904 308020
rect 250036 307980 250042 307992
rect 250898 307980 250904 307992
rect 250956 307980 250962 308032
rect 263778 307980 263784 308032
rect 263836 308020 263842 308032
rect 264698 308020 264704 308032
rect 263836 307992 264704 308020
rect 263836 307980 263842 307992
rect 264698 307980 264704 307992
rect 264756 307980 264762 308032
rect 267734 307980 267740 308032
rect 267792 308020 267798 308032
rect 268102 308020 268108 308032
rect 267792 307992 268108 308020
rect 267792 307980 267798 307992
rect 268102 307980 268108 307992
rect 268160 307980 268166 308032
rect 356054 307980 356060 308032
rect 356112 308020 356118 308032
rect 366450 308020 366456 308032
rect 356112 307992 366456 308020
rect 356112 307980 356118 307992
rect 366450 307980 366456 307992
rect 366508 307980 366514 308032
rect 256786 307912 256792 307964
rect 256844 307952 256850 307964
rect 257338 307952 257344 307964
rect 256844 307924 257344 307952
rect 256844 307912 256850 307924
rect 257338 307912 257344 307924
rect 257396 307912 257402 307964
rect 354674 307912 354680 307964
rect 354732 307952 354738 307964
rect 354732 307924 360056 307952
rect 354732 307912 354738 307924
rect 253198 307844 253204 307896
rect 253256 307884 253262 307896
rect 258994 307884 259000 307896
rect 253256 307856 259000 307884
rect 253256 307844 253262 307856
rect 258994 307844 259000 307856
rect 259052 307844 259058 307896
rect 360028 307884 360056 307924
rect 360102 307912 360108 307964
rect 360160 307952 360166 307964
rect 362770 307952 362776 307964
rect 360160 307924 362776 307952
rect 360160 307912 360166 307924
rect 362770 307912 362776 307924
rect 362828 307912 362834 307964
rect 360028 307856 360194 307884
rect 257338 307776 257344 307828
rect 257396 307816 257402 307828
rect 258258 307816 258264 307828
rect 257396 307788 258264 307816
rect 257396 307776 257402 307788
rect 258258 307776 258264 307788
rect 258316 307776 258322 307828
rect 260282 307776 260288 307828
rect 260340 307816 260346 307828
rect 262398 307816 262404 307828
rect 260340 307788 262404 307816
rect 260340 307776 260346 307788
rect 262398 307776 262404 307788
rect 262456 307776 262462 307828
rect 358170 307776 358176 307828
rect 358228 307816 358234 307828
rect 359550 307816 359556 307828
rect 358228 307788 359556 307816
rect 358228 307776 358234 307788
rect 359550 307776 359556 307788
rect 359608 307776 359614 307828
rect 360166 307816 360194 307856
rect 360930 307844 360936 307896
rect 360988 307884 360994 307896
rect 363690 307884 363696 307896
rect 360988 307856 363696 307884
rect 360988 307844 360994 307856
rect 363690 307844 363696 307856
rect 363748 307844 363754 307896
rect 360166 307788 360976 307816
rect 360948 307748 360976 307788
rect 361022 307776 361028 307828
rect 361080 307816 361086 307828
rect 361574 307816 361580 307828
rect 361080 307788 361580 307816
rect 361080 307776 361086 307788
rect 361574 307776 361580 307788
rect 361632 307776 361638 307828
rect 367370 307816 367376 307828
rect 361684 307788 367376 307816
rect 361684 307748 361712 307788
rect 367370 307776 367376 307788
rect 367428 307776 367434 307828
rect 360948 307720 361712 307748
rect 251358 307640 251364 307692
rect 251416 307680 251422 307692
rect 251910 307680 251916 307692
rect 251416 307652 251916 307680
rect 251416 307640 251422 307652
rect 251910 307640 251916 307652
rect 251968 307640 251974 307692
rect 267734 307640 267740 307692
rect 267792 307680 267798 307692
rect 268654 307680 268660 307692
rect 267792 307652 268660 307680
rect 267792 307640 267798 307652
rect 268654 307640 268660 307652
rect 268712 307640 268718 307692
rect 359826 307640 359832 307692
rect 359884 307680 359890 307692
rect 361390 307680 361396 307692
rect 359884 307652 361396 307680
rect 359884 307640 359890 307652
rect 361390 307640 361396 307652
rect 361448 307640 361454 307692
rect 266630 307504 266636 307556
rect 266688 307544 266694 307556
rect 266906 307544 266912 307556
rect 266688 307516 266912 307544
rect 266688 307504 266694 307516
rect 266906 307504 266912 307516
rect 266964 307504 266970 307556
rect 264974 307232 264980 307284
rect 265032 307272 265038 307284
rect 265894 307272 265900 307284
rect 265032 307244 265900 307272
rect 265032 307232 265038 307244
rect 265894 307232 265900 307244
rect 265952 307232 265958 307284
rect 202874 307164 202880 307216
rect 202932 307204 202938 307216
rect 271874 307204 271880 307216
rect 202932 307176 271880 307204
rect 202932 307164 202938 307176
rect 271874 307164 271880 307176
rect 271932 307164 271938 307216
rect 314838 307164 314844 307216
rect 314896 307204 314902 307216
rect 422294 307204 422300 307216
rect 314896 307176 422300 307204
rect 314896 307164 314902 307176
rect 422294 307164 422300 307176
rect 422352 307164 422358 307216
rect 189074 307096 189080 307148
rect 189132 307136 189138 307148
rect 269482 307136 269488 307148
rect 189132 307108 269488 307136
rect 189132 307096 189138 307108
rect 269482 307096 269488 307108
rect 269540 307096 269546 307148
rect 269574 307096 269580 307148
rect 269632 307096 269638 307148
rect 272058 307096 272064 307148
rect 272116 307136 272122 307148
rect 272242 307136 272248 307148
rect 272116 307108 272248 307136
rect 272116 307096 272122 307108
rect 272242 307096 272248 307108
rect 272300 307096 272306 307148
rect 321922 307096 321928 307148
rect 321980 307136 321986 307148
rect 458174 307136 458180 307148
rect 321980 307108 458180 307136
rect 321980 307096 321986 307108
rect 458174 307096 458180 307108
rect 458232 307096 458238 307148
rect 67634 307028 67640 307080
rect 67692 307068 67698 307080
rect 245562 307068 245568 307080
rect 67692 307040 245568 307068
rect 67692 307028 67698 307040
rect 245562 307028 245568 307040
rect 245620 307028 245626 307080
rect 245746 306960 245752 307012
rect 245804 307000 245810 307012
rect 246482 307000 246488 307012
rect 245804 306972 246488 307000
rect 245804 306960 245810 306972
rect 246482 306960 246488 306972
rect 246540 306960 246546 307012
rect 254302 306960 254308 307012
rect 254360 307000 254366 307012
rect 254486 307000 254492 307012
rect 254360 306972 254492 307000
rect 254360 306960 254366 306972
rect 254486 306960 254492 306972
rect 254544 306960 254550 307012
rect 261018 306960 261024 307012
rect 261076 306960 261082 307012
rect 261036 306808 261064 306960
rect 269592 306944 269620 307096
rect 480254 307068 480260 307080
rect 331186 307040 480260 307068
rect 272058 306960 272064 307012
rect 272116 307000 272122 307012
rect 272886 307000 272892 307012
rect 272116 306972 272892 307000
rect 272116 306960 272122 306972
rect 272886 306960 272892 306972
rect 272944 306960 272950 307012
rect 300854 306960 300860 307012
rect 300912 307000 300918 307012
rect 301130 307000 301136 307012
rect 300912 306972 301136 307000
rect 300912 306960 300918 306972
rect 301130 306960 301136 306972
rect 301188 306960 301194 307012
rect 317782 306960 317788 307012
rect 317840 306960 317846 307012
rect 326062 306960 326068 307012
rect 326120 307000 326126 307012
rect 331186 307000 331214 307040
rect 480254 307028 480260 307040
rect 480312 307028 480318 307080
rect 326120 306972 331214 307000
rect 326120 306960 326126 306972
rect 336826 306960 336832 307012
rect 336884 307000 336890 307012
rect 337010 307000 337016 307012
rect 336884 306972 337016 307000
rect 336884 306960 336890 306972
rect 337010 306960 337016 306972
rect 337068 306960 337074 307012
rect 269574 306892 269580 306944
rect 269632 306892 269638 306944
rect 317800 306808 317828 306960
rect 261018 306756 261024 306808
rect 261076 306756 261082 306808
rect 317782 306756 317788 306808
rect 317840 306756 317846 306808
rect 243262 306688 243268 306740
rect 243320 306688 243326 306740
rect 243280 306536 243308 306688
rect 299566 306552 299572 306604
rect 299624 306592 299630 306604
rect 300210 306592 300216 306604
rect 299624 306564 300216 306592
rect 299624 306552 299630 306564
rect 300210 306552 300216 306564
rect 300268 306552 300274 306604
rect 328638 306552 328644 306604
rect 328696 306592 328702 306604
rect 329006 306592 329012 306604
rect 328696 306564 329012 306592
rect 328696 306552 328702 306564
rect 329006 306552 329012 306564
rect 329064 306552 329070 306604
rect 332686 306552 332692 306604
rect 332744 306592 332750 306604
rect 332870 306592 332876 306604
rect 332744 306564 332876 306592
rect 332744 306552 332750 306564
rect 332870 306552 332876 306564
rect 332928 306552 332934 306604
rect 236086 306484 236092 306536
rect 236144 306524 236150 306536
rect 237282 306524 237288 306536
rect 236144 306496 237288 306524
rect 236144 306484 236150 306496
rect 237282 306484 237288 306496
rect 237340 306484 237346 306536
rect 243262 306484 243268 306536
rect 243320 306484 243326 306536
rect 279970 306524 279976 306536
rect 270466 306496 279976 306524
rect 234798 306416 234804 306468
rect 234856 306456 234862 306468
rect 235902 306456 235908 306468
rect 234856 306428 235908 306456
rect 234856 306416 234862 306428
rect 235902 306416 235908 306428
rect 235960 306416 235966 306468
rect 236178 306416 236184 306468
rect 236236 306456 236242 306468
rect 236822 306456 236828 306468
rect 236236 306428 236828 306456
rect 236236 306416 236242 306428
rect 236822 306416 236828 306428
rect 236880 306416 236886 306468
rect 237558 306416 237564 306468
rect 237616 306456 237622 306468
rect 237834 306456 237840 306468
rect 237616 306428 237840 306456
rect 237616 306416 237622 306428
rect 237834 306416 237840 306428
rect 237892 306416 237898 306468
rect 240226 306416 240232 306468
rect 240284 306456 240290 306468
rect 241054 306456 241060 306468
rect 240284 306428 241060 306456
rect 240284 306416 240290 306428
rect 241054 306416 241060 306428
rect 241112 306416 241118 306468
rect 243078 306416 243084 306468
rect 243136 306456 243142 306468
rect 244182 306456 244188 306468
rect 243136 306428 244188 306456
rect 243136 306416 243142 306428
rect 244182 306416 244188 306428
rect 244240 306416 244246 306468
rect 254026 306416 254032 306468
rect 254084 306456 254090 306468
rect 254670 306456 254676 306468
rect 254084 306428 254676 306456
rect 254084 306416 254090 306428
rect 254670 306416 254676 306428
rect 254728 306416 254734 306468
rect 255406 306416 255412 306468
rect 255464 306456 255470 306468
rect 256050 306456 256056 306468
rect 255464 306428 256056 306456
rect 255464 306416 255470 306428
rect 256050 306416 256056 306428
rect 256108 306416 256114 306468
rect 256970 306416 256976 306468
rect 257028 306456 257034 306468
rect 257430 306456 257436 306468
rect 257028 306428 257436 306456
rect 257028 306416 257034 306428
rect 257430 306416 257436 306428
rect 257488 306416 257494 306468
rect 259454 306416 259460 306468
rect 259512 306456 259518 306468
rect 259822 306456 259828 306468
rect 259512 306428 259828 306456
rect 259512 306416 259518 306428
rect 259822 306416 259828 306428
rect 259880 306416 259886 306468
rect 260834 306416 260840 306468
rect 260892 306456 260898 306468
rect 261202 306456 261208 306468
rect 260892 306428 261208 306456
rect 260892 306416 260898 306428
rect 261202 306416 261208 306428
rect 261260 306416 261266 306468
rect 234706 306348 234712 306400
rect 234764 306388 234770 306400
rect 235534 306388 235540 306400
rect 234764 306360 235540 306388
rect 234764 306348 234770 306360
rect 235534 306348 235540 306360
rect 235592 306348 235598 306400
rect 236270 306348 236276 306400
rect 236328 306388 236334 306400
rect 236914 306388 236920 306400
rect 236328 306360 236920 306388
rect 236328 306348 236334 306360
rect 236914 306348 236920 306360
rect 236972 306348 236978 306400
rect 237466 306348 237472 306400
rect 237524 306388 237530 306400
rect 238202 306388 238208 306400
rect 237524 306360 238208 306388
rect 237524 306348 237530 306360
rect 238202 306348 238208 306360
rect 238260 306348 238266 306400
rect 238846 306348 238852 306400
rect 238904 306388 238910 306400
rect 239582 306388 239588 306400
rect 238904 306360 239588 306388
rect 238904 306348 238910 306360
rect 239582 306348 239588 306360
rect 239640 306348 239646 306400
rect 240410 306348 240416 306400
rect 240468 306388 240474 306400
rect 240962 306388 240968 306400
rect 240468 306360 240968 306388
rect 240468 306348 240474 306360
rect 240962 306348 240968 306360
rect 241020 306348 241026 306400
rect 241606 306348 241612 306400
rect 241664 306388 241670 306400
rect 242342 306388 242348 306400
rect 241664 306360 242348 306388
rect 241664 306348 241670 306360
rect 242342 306348 242348 306360
rect 242400 306348 242406 306400
rect 242986 306348 242992 306400
rect 243044 306388 243050 306400
rect 243722 306388 243728 306400
rect 243044 306360 243728 306388
rect 243044 306348 243050 306360
rect 243722 306348 243728 306360
rect 243780 306348 243786 306400
rect 254210 306348 254216 306400
rect 254268 306388 254274 306400
rect 255038 306388 255044 306400
rect 254268 306360 255044 306388
rect 254268 306348 254274 306360
rect 255038 306348 255044 306360
rect 255096 306348 255102 306400
rect 255498 306348 255504 306400
rect 255556 306388 255562 306400
rect 255774 306388 255780 306400
rect 255556 306360 255780 306388
rect 255556 306348 255562 306360
rect 255774 306348 255780 306360
rect 255832 306348 255838 306400
rect 257154 306348 257160 306400
rect 257212 306388 257218 306400
rect 257798 306388 257804 306400
rect 257212 306360 257804 306388
rect 257212 306348 257218 306360
rect 257798 306348 257804 306360
rect 257856 306348 257862 306400
rect 261110 306348 261116 306400
rect 261168 306388 261174 306400
rect 261570 306388 261576 306400
rect 261168 306360 261576 306388
rect 261168 306348 261174 306360
rect 261570 306348 261576 306360
rect 261628 306348 261634 306400
rect 262398 306348 262404 306400
rect 262456 306388 262462 306400
rect 263318 306388 263324 306400
rect 262456 306360 263324 306388
rect 262456 306348 262462 306360
rect 263318 306348 263324 306360
rect 263376 306348 263382 306400
rect 216398 306280 216404 306332
rect 216456 306320 216462 306332
rect 270466 306320 270494 306496
rect 279970 306484 279976 306496
rect 280028 306484 280034 306536
rect 288526 306484 288532 306536
rect 288584 306524 288590 306536
rect 288584 306496 288940 306524
rect 288584 306484 288590 306496
rect 273070 306416 273076 306468
rect 273128 306456 273134 306468
rect 273128 306428 280154 306456
rect 273128 306416 273134 306428
rect 273346 306348 273352 306400
rect 273404 306388 273410 306400
rect 273806 306388 273812 306400
rect 273404 306360 273812 306388
rect 273404 306348 273410 306360
rect 273806 306348 273812 306360
rect 273864 306348 273870 306400
rect 216456 306292 270494 306320
rect 216456 306280 216462 306292
rect 273530 306280 273536 306332
rect 273588 306320 273594 306332
rect 274174 306320 274180 306332
rect 273588 306292 274180 306320
rect 273588 306280 273594 306292
rect 274174 306280 274180 306292
rect 274232 306280 274238 306332
rect 280126 306320 280154 306428
rect 280982 306416 280988 306468
rect 281040 306456 281046 306468
rect 285950 306456 285956 306468
rect 281040 306428 285956 306456
rect 281040 306416 281046 306428
rect 285950 306416 285956 306428
rect 286008 306416 286014 306468
rect 288802 306416 288808 306468
rect 288860 306416 288866 306468
rect 284294 306348 284300 306400
rect 284352 306388 284358 306400
rect 285490 306388 285496 306400
rect 284352 306360 285496 306388
rect 284352 306348 284358 306360
rect 285490 306348 285496 306360
rect 285548 306348 285554 306400
rect 281810 306320 281816 306332
rect 280126 306292 281816 306320
rect 281810 306280 281816 306292
rect 281868 306280 281874 306332
rect 284662 306280 284668 306332
rect 284720 306320 284726 306332
rect 285122 306320 285128 306332
rect 284720 306292 285128 306320
rect 284720 306280 284726 306292
rect 285122 306280 285128 306292
rect 285180 306280 285186 306332
rect 286042 306280 286048 306332
rect 286100 306320 286106 306332
rect 286870 306320 286876 306332
rect 286100 306292 286876 306320
rect 286100 306280 286106 306292
rect 286870 306280 286876 306292
rect 286928 306280 286934 306332
rect 218698 306212 218704 306264
rect 218756 306252 218762 306264
rect 273070 306252 273076 306264
rect 218756 306224 273076 306252
rect 218756 306212 218762 306224
rect 273070 306212 273076 306224
rect 273128 306212 273134 306264
rect 284386 306212 284392 306264
rect 284444 306252 284450 306264
rect 284570 306252 284576 306264
rect 284444 306224 284576 306252
rect 284444 306212 284450 306224
rect 284570 306212 284576 306224
rect 284628 306212 284634 306264
rect 285766 306212 285772 306264
rect 285824 306252 285830 306264
rect 286134 306252 286140 306264
rect 285824 306224 286140 306252
rect 285824 306212 285830 306224
rect 286134 306212 286140 306224
rect 286192 306212 286198 306264
rect 288618 306212 288624 306264
rect 288676 306252 288682 306264
rect 288820 306252 288848 306416
rect 288912 306264 288940 306496
rect 296806 306484 296812 306536
rect 296864 306524 296870 306536
rect 297174 306524 297180 306536
rect 296864 306496 297180 306524
rect 296864 306484 296870 306496
rect 297174 306484 297180 306496
rect 297232 306484 297238 306536
rect 342714 306524 342720 306536
rect 342272 306496 342720 306524
rect 292942 306456 292948 306468
rect 292684 306428 292948 306456
rect 292684 306400 292712 306428
rect 292942 306416 292948 306428
rect 293000 306416 293006 306468
rect 327074 306416 327080 306468
rect 327132 306456 327138 306468
rect 327442 306456 327448 306468
rect 327132 306428 327448 306456
rect 327132 306416 327138 306428
rect 327442 306416 327448 306428
rect 327500 306416 327506 306468
rect 289814 306348 289820 306400
rect 289872 306388 289878 306400
rect 291010 306388 291016 306400
rect 289872 306360 291016 306388
rect 289872 306348 289878 306360
rect 291010 306348 291016 306360
rect 291068 306348 291074 306400
rect 292666 306348 292672 306400
rect 292724 306348 292730 306400
rect 298094 306348 298100 306400
rect 298152 306388 298158 306400
rect 298646 306388 298652 306400
rect 298152 306360 298652 306388
rect 298152 306348 298158 306360
rect 298646 306348 298652 306360
rect 298704 306348 298710 306400
rect 302418 306348 302424 306400
rect 302476 306388 302482 306400
rect 302878 306388 302884 306400
rect 302476 306360 302884 306388
rect 302476 306348 302482 306360
rect 302878 306348 302884 306360
rect 302936 306348 302942 306400
rect 305086 306348 305092 306400
rect 305144 306388 305150 306400
rect 306006 306388 306012 306400
rect 305144 306360 306012 306388
rect 305144 306348 305150 306360
rect 306006 306348 306012 306360
rect 306064 306348 306070 306400
rect 307846 306348 307852 306400
rect 307904 306388 307910 306400
rect 308766 306388 308772 306400
rect 307904 306360 308772 306388
rect 307904 306348 307910 306360
rect 308766 306348 308772 306360
rect 308824 306348 308830 306400
rect 316126 306348 316132 306400
rect 316184 306388 316190 306400
rect 316954 306388 316960 306400
rect 316184 306360 316960 306388
rect 316184 306348 316190 306360
rect 316954 306348 316960 306360
rect 317012 306348 317018 306400
rect 321646 306348 321652 306400
rect 321704 306388 321710 306400
rect 322474 306388 322480 306400
rect 321704 306360 322480 306388
rect 321704 306348 321710 306360
rect 322474 306348 322480 306360
rect 322532 306348 322538 306400
rect 324314 306348 324320 306400
rect 324372 306388 324378 306400
rect 325234 306388 325240 306400
rect 324372 306360 325240 306388
rect 324372 306348 324378 306360
rect 325234 306348 325240 306360
rect 325292 306348 325298 306400
rect 328454 306348 328460 306400
rect 328512 306388 328518 306400
rect 329282 306388 329288 306400
rect 328512 306360 329288 306388
rect 328512 306348 328518 306360
rect 329282 306348 329288 306360
rect 329340 306348 329346 306400
rect 329926 306348 329932 306400
rect 329984 306388 329990 306400
rect 330202 306388 330208 306400
rect 329984 306360 330208 306388
rect 329984 306348 329990 306360
rect 330202 306348 330208 306360
rect 330260 306348 330266 306400
rect 331582 306348 331588 306400
rect 331640 306388 331646 306400
rect 331950 306388 331956 306400
rect 331640 306360 331956 306388
rect 331640 306348 331646 306360
rect 331950 306348 331956 306360
rect 332008 306348 332014 306400
rect 289906 306280 289912 306332
rect 289964 306320 289970 306332
rect 290182 306320 290188 306332
rect 289964 306292 290188 306320
rect 289964 306280 289970 306292
rect 290182 306280 290188 306292
rect 290240 306280 290246 306332
rect 291286 306280 291292 306332
rect 291344 306320 291350 306332
rect 291930 306320 291936 306332
rect 291344 306292 291936 306320
rect 291344 306280 291350 306292
rect 291930 306280 291936 306292
rect 291988 306280 291994 306332
rect 293954 306280 293960 306332
rect 294012 306320 294018 306332
rect 295150 306320 295156 306332
rect 294012 306292 295156 306320
rect 294012 306280 294018 306292
rect 295150 306280 295156 306292
rect 295208 306280 295214 306332
rect 298278 306280 298284 306332
rect 298336 306320 298342 306332
rect 298738 306320 298744 306332
rect 298336 306292 298744 306320
rect 298336 306280 298342 306292
rect 298738 306280 298744 306292
rect 298796 306280 298802 306332
rect 299566 306280 299572 306332
rect 299624 306320 299630 306332
rect 300486 306320 300492 306332
rect 299624 306292 300492 306320
rect 299624 306280 299630 306292
rect 300486 306280 300492 306292
rect 300544 306280 300550 306332
rect 300946 306280 300952 306332
rect 301004 306320 301010 306332
rect 301958 306320 301964 306332
rect 301004 306292 301964 306320
rect 301004 306280 301010 306292
rect 301958 306280 301964 306292
rect 302016 306280 302022 306332
rect 302602 306280 302608 306332
rect 302660 306320 302666 306332
rect 303246 306320 303252 306332
rect 302660 306292 303252 306320
rect 302660 306280 302666 306292
rect 303246 306280 303252 306292
rect 303304 306280 303310 306332
rect 305178 306280 305184 306332
rect 305236 306320 305242 306332
rect 306098 306320 306104 306332
rect 305236 306292 306104 306320
rect 305236 306280 305242 306292
rect 306098 306280 306104 306292
rect 306156 306280 306162 306332
rect 306374 306280 306380 306332
rect 306432 306320 306438 306332
rect 307478 306320 307484 306332
rect 306432 306292 307484 306320
rect 306432 306280 306438 306292
rect 307478 306280 307484 306292
rect 307536 306280 307542 306332
rect 307754 306280 307760 306332
rect 307812 306320 307818 306332
rect 308306 306320 308312 306332
rect 307812 306292 308312 306320
rect 307812 306280 307818 306292
rect 308306 306280 308312 306292
rect 308364 306280 308370 306332
rect 309226 306280 309232 306332
rect 309284 306320 309290 306332
rect 310146 306320 310152 306332
rect 309284 306292 310152 306320
rect 309284 306280 309290 306292
rect 310146 306280 310152 306292
rect 310204 306280 310210 306332
rect 310514 306280 310520 306332
rect 310572 306320 310578 306332
rect 311526 306320 311532 306332
rect 310572 306292 311532 306320
rect 310572 306280 310578 306292
rect 311526 306280 311532 306292
rect 311584 306280 311590 306332
rect 311986 306280 311992 306332
rect 312044 306320 312050 306332
rect 312906 306320 312912 306332
rect 312044 306292 312912 306320
rect 312044 306280 312050 306292
rect 312906 306280 312912 306292
rect 312964 306280 312970 306332
rect 314746 306280 314752 306332
rect 314804 306320 314810 306332
rect 315574 306320 315580 306332
rect 314804 306292 315580 306320
rect 314804 306280 314810 306292
rect 315574 306280 315580 306292
rect 315632 306280 315638 306332
rect 316034 306280 316040 306332
rect 316092 306320 316098 306332
rect 316862 306320 316868 306332
rect 316092 306292 316868 306320
rect 316092 306280 316098 306292
rect 316862 306280 316868 306292
rect 316920 306280 316926 306332
rect 317690 306280 317696 306332
rect 317748 306320 317754 306332
rect 318242 306320 318248 306332
rect 317748 306292 318248 306320
rect 317748 306280 317754 306292
rect 318242 306280 318248 306292
rect 318300 306280 318306 306332
rect 318794 306280 318800 306332
rect 318852 306320 318858 306332
rect 320082 306320 320088 306332
rect 318852 306292 320088 306320
rect 318852 306280 318858 306292
rect 320082 306280 320088 306292
rect 320140 306280 320146 306332
rect 320174 306280 320180 306332
rect 320232 306320 320238 306332
rect 321462 306320 321468 306332
rect 320232 306292 321468 306320
rect 320232 306280 320238 306292
rect 321462 306280 321468 306292
rect 321520 306280 321526 306332
rect 321554 306280 321560 306332
rect 321612 306320 321618 306332
rect 322382 306320 322388 306332
rect 321612 306292 322388 306320
rect 321612 306280 321618 306292
rect 322382 306280 322388 306292
rect 322440 306280 322446 306332
rect 323026 306280 323032 306332
rect 323084 306320 323090 306332
rect 323394 306320 323400 306332
rect 323084 306292 323400 306320
rect 323084 306280 323090 306292
rect 323394 306280 323400 306292
rect 323452 306280 323458 306332
rect 324406 306280 324412 306332
rect 324464 306320 324470 306332
rect 325142 306320 325148 306332
rect 324464 306292 325148 306320
rect 324464 306280 324470 306292
rect 325142 306280 325148 306292
rect 325200 306280 325206 306332
rect 325786 306280 325792 306332
rect 325844 306320 325850 306332
rect 326614 306320 326620 306332
rect 325844 306292 326620 306320
rect 325844 306280 325850 306292
rect 326614 306280 326620 306292
rect 326672 306280 326678 306332
rect 327166 306280 327172 306332
rect 327224 306320 327230 306332
rect 327994 306320 328000 306332
rect 327224 306292 328000 306320
rect 327224 306280 327230 306292
rect 327994 306280 328000 306292
rect 328052 306280 328058 306332
rect 328638 306280 328644 306332
rect 328696 306320 328702 306332
rect 329374 306320 329380 306332
rect 328696 306292 329380 306320
rect 328696 306280 328702 306292
rect 329374 306280 329380 306292
rect 329432 306280 329438 306332
rect 329834 306280 329840 306332
rect 329892 306320 329898 306332
rect 330294 306320 330300 306332
rect 329892 306292 330300 306320
rect 329892 306280 329898 306292
rect 330294 306280 330300 306292
rect 330352 306280 330358 306332
rect 331490 306280 331496 306332
rect 331548 306320 331554 306332
rect 331858 306320 331864 306332
rect 331548 306292 331864 306320
rect 331548 306280 331554 306292
rect 331858 306280 331864 306292
rect 331916 306280 331922 306332
rect 335630 306280 335636 306332
rect 335688 306320 335694 306332
rect 335998 306320 336004 306332
rect 335688 306292 336004 306320
rect 335688 306280 335694 306292
rect 335998 306280 336004 306292
rect 336056 306280 336062 306332
rect 337102 306280 337108 306332
rect 337160 306320 337166 306332
rect 337470 306320 337476 306332
rect 337160 306292 337476 306320
rect 337160 306280 337166 306292
rect 337470 306280 337476 306292
rect 337528 306280 337534 306332
rect 341150 306280 341156 306332
rect 341208 306320 341214 306332
rect 341518 306320 341524 306332
rect 341208 306292 341524 306320
rect 341208 306280 341214 306292
rect 341518 306280 341524 306292
rect 341576 306280 341582 306332
rect 342272 306264 342300 306496
rect 342714 306484 342720 306496
rect 342772 306484 342778 306536
rect 342622 306416 342628 306468
rect 342680 306416 342686 306468
rect 343634 306416 343640 306468
rect 343692 306456 343698 306468
rect 344002 306456 344008 306468
rect 343692 306428 344008 306456
rect 343692 306416 343698 306428
rect 344002 306416 344008 306428
rect 344060 306416 344066 306468
rect 357710 306416 357716 306468
rect 357768 306456 357774 306468
rect 357986 306456 357992 306468
rect 357768 306428 357992 306456
rect 357768 306416 357774 306428
rect 357986 306416 357992 306428
rect 358044 306416 358050 306468
rect 358354 306416 358360 306468
rect 358412 306456 358418 306468
rect 360010 306456 360016 306468
rect 358412 306428 360016 306456
rect 358412 306416 358418 306428
rect 360010 306416 360016 306428
rect 360068 306416 360074 306468
rect 360286 306416 360292 306468
rect 360344 306456 360350 306468
rect 360746 306456 360752 306468
rect 360344 306428 360752 306456
rect 360344 306416 360350 306428
rect 360746 306416 360752 306428
rect 360804 306416 360810 306468
rect 288676 306224 288848 306252
rect 288676 306212 288682 306224
rect 288894 306212 288900 306264
rect 288952 306212 288958 306264
rect 291470 306212 291476 306264
rect 291528 306252 291534 306264
rect 292390 306252 292396 306264
rect 291528 306224 292396 306252
rect 291528 306212 291534 306224
rect 292390 306212 292396 306224
rect 292448 306212 292454 306264
rect 292850 306212 292856 306264
rect 292908 306252 292914 306264
rect 293770 306252 293776 306264
rect 292908 306224 293776 306252
rect 292908 306212 292914 306224
rect 293770 306212 293776 306224
rect 293828 306212 293834 306264
rect 296898 306212 296904 306264
rect 296956 306252 296962 306264
rect 297542 306252 297548 306264
rect 296956 306224 297548 306252
rect 296956 306212 296962 306224
rect 297542 306212 297548 306224
rect 297600 306212 297606 306264
rect 298186 306212 298192 306264
rect 298244 306252 298250 306264
rect 299198 306252 299204 306264
rect 298244 306224 299204 306252
rect 298244 306212 298250 306224
rect 299198 306212 299204 306224
rect 299256 306212 299262 306264
rect 302326 306212 302332 306264
rect 302384 306252 302390 306264
rect 303338 306252 303344 306264
rect 302384 306224 303344 306252
rect 302384 306212 302390 306224
rect 303338 306212 303344 306224
rect 303396 306212 303402 306264
rect 303614 306212 303620 306264
rect 303672 306252 303678 306264
rect 304074 306252 304080 306264
rect 303672 306224 304080 306252
rect 303672 306212 303678 306224
rect 304074 306212 304080 306224
rect 304132 306212 304138 306264
rect 321738 306212 321744 306264
rect 321796 306252 321802 306264
rect 322014 306252 322020 306264
rect 321796 306224 322020 306252
rect 321796 306212 321802 306224
rect 322014 306212 322020 306224
rect 322072 306212 322078 306264
rect 323118 306212 323124 306264
rect 323176 306252 323182 306264
rect 323854 306252 323860 306264
rect 323176 306224 323860 306252
rect 323176 306212 323182 306224
rect 323854 306212 323860 306224
rect 323912 306212 323918 306264
rect 325970 306212 325976 306264
rect 326028 306252 326034 306264
rect 326982 306252 326988 306264
rect 326028 306224 326988 306252
rect 326028 306212 326034 306224
rect 326982 306212 326988 306224
rect 327040 306212 327046 306264
rect 327258 306212 327264 306264
rect 327316 306252 327322 306264
rect 327534 306252 327540 306264
rect 327316 306224 327540 306252
rect 327316 306212 327322 306224
rect 327534 306212 327540 306224
rect 327592 306212 327598 306264
rect 328822 306212 328828 306264
rect 328880 306252 328886 306264
rect 329742 306252 329748 306264
rect 328880 306224 329748 306252
rect 328880 306212 328886 306224
rect 329742 306212 329748 306224
rect 329800 306212 329806 306264
rect 331306 306212 331312 306264
rect 331364 306252 331370 306264
rect 332318 306252 332324 306264
rect 331364 306224 332324 306252
rect 331364 306212 331370 306224
rect 332318 306212 332324 306224
rect 332376 306212 332382 306264
rect 332594 306212 332600 306264
rect 332652 306252 332658 306264
rect 332962 306252 332968 306264
rect 332652 306224 332968 306252
rect 332652 306212 332658 306224
rect 332962 306212 332968 306224
rect 333020 306212 333026 306264
rect 340966 306212 340972 306264
rect 341024 306252 341030 306264
rect 341334 306252 341340 306264
rect 341024 306224 341340 306252
rect 341024 306212 341030 306224
rect 341334 306212 341340 306224
rect 341392 306212 341398 306264
rect 342254 306212 342260 306264
rect 342312 306212 342318 306264
rect 214558 306144 214564 306196
rect 214616 306184 214622 306196
rect 277854 306184 277860 306196
rect 214616 306156 277860 306184
rect 214616 306144 214622 306156
rect 277854 306144 277860 306156
rect 277912 306144 277918 306196
rect 285858 306144 285864 306196
rect 285916 306184 285922 306196
rect 286502 306184 286508 306196
rect 285916 306156 286508 306184
rect 285916 306144 285922 306156
rect 286502 306144 286508 306156
rect 286560 306144 286566 306196
rect 288710 306144 288716 306196
rect 288768 306184 288774 306196
rect 289630 306184 289636 306196
rect 288768 306156 289636 306184
rect 288768 306144 288774 306156
rect 289630 306144 289636 306156
rect 289688 306144 289694 306196
rect 294046 306144 294052 306196
rect 294104 306184 294110 306196
rect 294690 306184 294696 306196
rect 294104 306156 294696 306184
rect 294104 306144 294110 306156
rect 294690 306144 294696 306156
rect 294748 306144 294754 306196
rect 296806 306144 296812 306196
rect 296864 306184 296870 306196
rect 297910 306184 297916 306196
rect 296864 306156 297916 306184
rect 296864 306144 296870 306156
rect 297910 306144 297916 306156
rect 297968 306144 297974 306196
rect 303982 306144 303988 306196
rect 304040 306184 304046 306196
rect 304718 306184 304724 306196
rect 304040 306156 304724 306184
rect 304040 306144 304046 306156
rect 304718 306144 304724 306156
rect 304776 306144 304782 306196
rect 319162 306144 319168 306196
rect 319220 306184 319226 306196
rect 319622 306184 319628 306196
rect 319220 306156 319628 306184
rect 319220 306144 319226 306156
rect 319622 306144 319628 306156
rect 319680 306144 319686 306196
rect 320542 306144 320548 306196
rect 320600 306184 320606 306196
rect 321094 306184 321100 306196
rect 320600 306156 321100 306184
rect 320600 306144 320606 306156
rect 321094 306144 321100 306156
rect 321152 306144 321158 306196
rect 321830 306144 321836 306196
rect 321888 306184 321894 306196
rect 322842 306184 322848 306196
rect 321888 306156 322848 306184
rect 321888 306144 321894 306156
rect 322842 306144 322848 306156
rect 322900 306144 322906 306196
rect 327350 306144 327356 306196
rect 327408 306184 327414 306196
rect 328362 306184 328368 306196
rect 327408 306156 328368 306184
rect 327408 306144 327414 306156
rect 328362 306144 328368 306156
rect 328420 306144 328426 306196
rect 333974 306144 333980 306196
rect 334032 306184 334038 306196
rect 334434 306184 334440 306196
rect 334032 306156 334440 306184
rect 334032 306144 334038 306156
rect 334434 306144 334440 306156
rect 334492 306144 334498 306196
rect 335354 306144 335360 306196
rect 335412 306184 335418 306196
rect 335814 306184 335820 306196
rect 335412 306156 335820 306184
rect 335412 306144 335418 306156
rect 335814 306144 335820 306156
rect 335872 306144 335878 306196
rect 337010 306144 337016 306196
rect 337068 306184 337074 306196
rect 337838 306184 337844 306196
rect 337068 306156 337844 306184
rect 337068 306144 337074 306156
rect 337838 306144 337844 306156
rect 337896 306144 337902 306196
rect 338206 306144 338212 306196
rect 338264 306184 338270 306196
rect 338574 306184 338580 306196
rect 338264 306156 338580 306184
rect 338264 306144 338270 306156
rect 338574 306144 338580 306156
rect 338632 306144 338638 306196
rect 339494 306144 339500 306196
rect 339552 306184 339558 306196
rect 339954 306184 339960 306196
rect 339552 306156 339960 306184
rect 339552 306144 339558 306156
rect 339954 306144 339960 306156
rect 340012 306144 340018 306196
rect 340874 306144 340880 306196
rect 340932 306184 340938 306196
rect 341978 306184 341984 306196
rect 340932 306156 341984 306184
rect 340932 306144 340938 306156
rect 341978 306144 341984 306156
rect 342036 306144 342042 306196
rect 216306 306076 216312 306128
rect 216364 306116 216370 306128
rect 281074 306116 281080 306128
rect 216364 306088 281080 306116
rect 216364 306076 216370 306088
rect 281074 306076 281080 306088
rect 281132 306076 281138 306128
rect 284386 306076 284392 306128
rect 284444 306116 284450 306128
rect 285030 306116 285036 306128
rect 284444 306088 285036 306116
rect 284444 306076 284450 306088
rect 285030 306076 285036 306088
rect 285088 306076 285094 306128
rect 288526 306076 288532 306128
rect 288584 306116 288590 306128
rect 289170 306116 289176 306128
rect 288584 306088 289176 306116
rect 288584 306076 288590 306088
rect 289170 306076 289176 306088
rect 289228 306076 289234 306128
rect 295334 306076 295340 306128
rect 295392 306116 295398 306128
rect 295702 306116 295708 306128
rect 295392 306088 295708 306116
rect 295392 306076 295398 306088
rect 295702 306076 295708 306088
rect 295760 306076 295766 306128
rect 299842 306076 299848 306128
rect 299900 306116 299906 306128
rect 300578 306116 300584 306128
rect 299900 306088 300584 306116
rect 299900 306076 299906 306088
rect 300578 306076 300584 306088
rect 300636 306076 300642 306128
rect 303798 306076 303804 306128
rect 303856 306116 303862 306128
rect 304626 306116 304632 306128
rect 303856 306088 304632 306116
rect 303856 306076 303862 306088
rect 304626 306076 304632 306088
rect 304684 306076 304690 306128
rect 313458 306076 313464 306128
rect 313516 306116 313522 306128
rect 314286 306116 314292 306128
rect 313516 306088 314292 306116
rect 313516 306076 313522 306088
rect 314286 306076 314292 306088
rect 314344 306076 314350 306128
rect 319070 306076 319076 306128
rect 319128 306116 319134 306128
rect 319714 306116 319720 306128
rect 319128 306088 319720 306116
rect 319128 306076 319134 306088
rect 319714 306076 319720 306088
rect 319772 306076 319778 306128
rect 330018 306076 330024 306128
rect 330076 306116 330082 306128
rect 330754 306116 330760 306128
rect 330076 306088 330760 306116
rect 330076 306076 330082 306088
rect 330754 306076 330760 306088
rect 330812 306076 330818 306128
rect 332594 306076 332600 306128
rect 332652 306116 332658 306128
rect 333330 306116 333336 306128
rect 332652 306088 333336 306116
rect 332652 306076 332658 306088
rect 333330 306076 333336 306088
rect 333388 306076 333394 306128
rect 334158 306076 334164 306128
rect 334216 306116 334222 306128
rect 335078 306116 335084 306128
rect 334216 306088 335084 306116
rect 334216 306076 334222 306088
rect 335078 306076 335084 306088
rect 335136 306076 335142 306128
rect 336734 306076 336740 306128
rect 336792 306116 336798 306128
rect 337378 306116 337384 306128
rect 336792 306088 337384 306116
rect 336792 306076 336798 306088
rect 337378 306076 337384 306088
rect 337436 306076 337442 306128
rect 338390 306076 338396 306128
rect 338448 306116 338454 306128
rect 339218 306116 339224 306128
rect 338448 306088 339224 306116
rect 338448 306076 338454 306088
rect 339218 306076 339224 306088
rect 339276 306076 339282 306128
rect 339586 306076 339592 306128
rect 339644 306116 339650 306128
rect 340598 306116 340604 306128
rect 339644 306088 340604 306116
rect 339644 306076 339650 306088
rect 340598 306076 340604 306088
rect 340656 306076 340662 306128
rect 342640 306116 342668 306416
rect 360194 306388 360200 306400
rect 357406 306360 360200 306388
rect 355870 306280 355876 306332
rect 355928 306320 355934 306332
rect 357406 306320 357434 306360
rect 360194 306348 360200 306360
rect 360252 306348 360258 306400
rect 360470 306348 360476 306400
rect 360528 306388 360534 306400
rect 361114 306388 361120 306400
rect 360528 306360 361120 306388
rect 360528 306348 360534 306360
rect 361114 306348 361120 306360
rect 361172 306348 361178 306400
rect 363046 306348 363052 306400
rect 363104 306388 363110 306400
rect 363230 306388 363236 306400
rect 363104 306360 363236 306388
rect 363104 306348 363110 306360
rect 363230 306348 363236 306360
rect 363288 306348 363294 306400
rect 371418 306320 371424 306332
rect 355928 306292 357434 306320
rect 358556 306292 371424 306320
rect 355928 306280 355934 306292
rect 343726 306212 343732 306264
rect 343784 306252 343790 306264
rect 344738 306252 344744 306264
rect 343784 306224 344744 306252
rect 343784 306212 343790 306224
rect 344738 306212 344744 306224
rect 344796 306212 344802 306264
rect 345014 306212 345020 306264
rect 345072 306252 345078 306264
rect 345474 306252 345480 306264
rect 345072 306224 345480 306252
rect 345072 306212 345078 306224
rect 345474 306212 345480 306224
rect 345532 306212 345538 306264
rect 357618 306212 357624 306264
rect 357676 306252 357682 306264
rect 358078 306252 358084 306264
rect 357676 306224 358084 306252
rect 357676 306212 357682 306224
rect 358078 306212 358084 306224
rect 358136 306212 358142 306264
rect 354950 306144 354956 306196
rect 355008 306184 355014 306196
rect 358556 306184 358584 306292
rect 371418 306280 371424 306292
rect 371476 306280 371482 306332
rect 359918 306252 359924 306264
rect 355008 306156 358584 306184
rect 358648 306224 359924 306252
rect 355008 306144 355014 306156
rect 342806 306116 342812 306128
rect 342640 306088 342812 306116
rect 342806 306076 342812 306088
rect 342864 306076 342870 306128
rect 357802 306076 357808 306128
rect 357860 306116 357866 306128
rect 358078 306116 358084 306128
rect 357860 306088 358084 306116
rect 357860 306076 357866 306088
rect 358078 306076 358084 306088
rect 358136 306076 358142 306128
rect 358648 306116 358676 306224
rect 359918 306212 359924 306224
rect 359976 306212 359982 306264
rect 360194 306212 360200 306264
rect 360252 306252 360258 306264
rect 371326 306252 371332 306264
rect 360252 306224 371332 306252
rect 360252 306212 360258 306224
rect 371326 306212 371332 306224
rect 371384 306212 371390 306264
rect 369210 306184 369216 306196
rect 358556 306088 358676 306116
rect 358740 306156 369216 306184
rect 215018 306008 215024 306060
rect 215076 306048 215082 306060
rect 279234 306048 279240 306060
rect 215076 306020 279240 306048
rect 215076 306008 215082 306020
rect 279234 306008 279240 306020
rect 279292 306008 279298 306060
rect 288802 306008 288808 306060
rect 288860 306048 288866 306060
rect 289262 306048 289268 306060
rect 288860 306020 289268 306048
rect 288860 306008 288866 306020
rect 289262 306008 289268 306020
rect 289320 306008 289326 306060
rect 295610 306008 295616 306060
rect 295668 306048 295674 306060
rect 296530 306048 296536 306060
rect 295668 306020 296536 306048
rect 295668 306008 295674 306020
rect 296530 306008 296536 306020
rect 296588 306008 296594 306060
rect 303614 306008 303620 306060
rect 303672 306048 303678 306060
rect 304258 306048 304264 306060
rect 303672 306020 304264 306048
rect 303672 306008 303678 306020
rect 304258 306008 304264 306020
rect 304316 306008 304322 306060
rect 332778 306008 332784 306060
rect 332836 306048 332842 306060
rect 333698 306048 333704 306060
rect 332836 306020 333704 306048
rect 332836 306008 332842 306020
rect 333698 306008 333704 306020
rect 333756 306008 333762 306060
rect 333974 306008 333980 306060
rect 334032 306048 334038 306060
rect 334710 306048 334716 306060
rect 334032 306020 334716 306048
rect 334032 306008 334038 306020
rect 334710 306008 334716 306020
rect 334768 306008 334774 306060
rect 338206 306008 338212 306060
rect 338264 306048 338270 306060
rect 338850 306048 338856 306060
rect 338264 306020 338856 306048
rect 338264 306008 338270 306020
rect 338850 306008 338856 306020
rect 338908 306008 338914 306060
rect 342346 306008 342352 306060
rect 342404 306048 342410 306060
rect 343358 306048 343364 306060
rect 342404 306020 343364 306048
rect 342404 306008 342410 306020
rect 343358 306008 343364 306020
rect 343416 306008 343422 306060
rect 355502 306008 355508 306060
rect 355560 306048 355566 306060
rect 358556 306048 358584 306088
rect 355560 306020 358584 306048
rect 355560 306008 355566 306020
rect 214650 305940 214656 305992
rect 214708 305980 214714 305992
rect 280614 305980 280620 305992
rect 214708 305952 280620 305980
rect 214708 305940 214714 305952
rect 280614 305940 280620 305952
rect 280672 305940 280678 305992
rect 295334 305940 295340 305992
rect 295392 305980 295398 305992
rect 296162 305980 296168 305992
rect 295392 305952 296168 305980
rect 295392 305940 295398 305952
rect 296162 305940 296168 305952
rect 296220 305940 296226 305992
rect 354030 305940 354036 305992
rect 354088 305980 354094 305992
rect 358354 305980 358360 305992
rect 354088 305952 358360 305980
rect 354088 305940 354094 305952
rect 358354 305940 358360 305952
rect 358412 305940 358418 305992
rect 358740 305980 358768 306156
rect 369210 306144 369216 306156
rect 369268 306144 369274 306196
rect 359918 306076 359924 306128
rect 359976 306116 359982 306128
rect 371878 306116 371884 306128
rect 359976 306088 371884 306116
rect 359976 306076 359982 306088
rect 371878 306076 371884 306088
rect 371936 306076 371942 306128
rect 360010 306008 360016 306060
rect 360068 306048 360074 306060
rect 371510 306048 371516 306060
rect 360068 306020 371516 306048
rect 360068 306008 360074 306020
rect 371510 306008 371516 306020
rect 371568 306008 371574 306060
rect 358464 305952 358768 305980
rect 213730 305872 213736 305924
rect 213788 305912 213794 305924
rect 282730 305912 282736 305924
rect 213788 305884 282736 305912
rect 213788 305872 213794 305884
rect 282730 305872 282736 305884
rect 282788 305872 282794 305924
rect 352834 305872 352840 305924
rect 352892 305912 352898 305924
rect 358464 305912 358492 305952
rect 358814 305940 358820 305992
rect 358872 305980 358878 305992
rect 369026 305980 369032 305992
rect 358872 305952 369032 305980
rect 358872 305940 358878 305952
rect 369026 305940 369032 305952
rect 369084 305940 369090 305992
rect 352892 305884 358492 305912
rect 352892 305872 352898 305884
rect 358538 305872 358544 305924
rect 358596 305912 358602 305924
rect 370406 305912 370412 305924
rect 358596 305884 370412 305912
rect 358596 305872 358602 305884
rect 370406 305872 370412 305884
rect 370464 305872 370470 305924
rect 214466 305804 214472 305856
rect 214524 305844 214530 305856
rect 283466 305844 283472 305856
rect 214524 305816 283472 305844
rect 214524 305804 214530 305816
rect 283466 305804 283472 305816
rect 283524 305804 283530 305856
rect 354490 305804 354496 305856
rect 354548 305844 354554 305856
rect 371786 305844 371792 305856
rect 354548 305816 371792 305844
rect 354548 305804 354554 305816
rect 371786 305804 371792 305816
rect 371844 305804 371850 305856
rect 216122 305736 216128 305788
rect 216180 305776 216186 305788
rect 288066 305776 288072 305788
rect 216180 305748 288072 305776
rect 216180 305736 216186 305748
rect 288066 305736 288072 305748
rect 288124 305736 288130 305788
rect 350074 305736 350080 305788
rect 350132 305776 350138 305788
rect 368934 305776 368940 305788
rect 350132 305748 368940 305776
rect 350132 305736 350138 305748
rect 368934 305736 368940 305748
rect 368992 305736 368998 305788
rect 214742 305668 214748 305720
rect 214800 305708 214806 305720
rect 287606 305708 287612 305720
rect 214800 305680 287612 305708
rect 214800 305668 214806 305680
rect 287606 305668 287612 305680
rect 287664 305668 287670 305720
rect 352190 305668 352196 305720
rect 352248 305708 352254 305720
rect 358538 305708 358544 305720
rect 352248 305680 358544 305708
rect 352248 305668 352254 305680
rect 358538 305668 358544 305680
rect 358596 305668 358602 305720
rect 358722 305668 358728 305720
rect 358780 305708 358786 305720
rect 370314 305708 370320 305720
rect 358780 305680 370320 305708
rect 358780 305668 358786 305680
rect 370314 305668 370320 305680
rect 370372 305668 370378 305720
rect 217686 305600 217692 305652
rect 217744 305640 217750 305652
rect 345658 305640 345664 305652
rect 217744 305612 345664 305640
rect 217744 305600 217750 305612
rect 345658 305600 345664 305612
rect 345716 305600 345722 305652
rect 346578 305600 346584 305652
rect 346636 305640 346642 305652
rect 369302 305640 369308 305652
rect 346636 305612 369308 305640
rect 346636 305600 346642 305612
rect 369302 305600 369308 305612
rect 369360 305600 369366 305652
rect 215110 305532 215116 305584
rect 215168 305572 215174 305584
rect 276474 305572 276480 305584
rect 215168 305544 276480 305572
rect 215168 305532 215174 305544
rect 276474 305532 276480 305544
rect 276532 305532 276538 305584
rect 348234 305532 348240 305584
rect 348292 305572 348298 305584
rect 363782 305572 363788 305584
rect 348292 305544 363788 305572
rect 348292 305532 348298 305544
rect 363782 305532 363788 305544
rect 363840 305532 363846 305584
rect 216582 305464 216588 305516
rect 216640 305504 216646 305516
rect 278590 305504 278596 305516
rect 216640 305476 278596 305504
rect 216640 305464 216646 305476
rect 278590 305464 278596 305476
rect 278648 305464 278654 305516
rect 357342 305464 357348 305516
rect 357400 305504 357406 305516
rect 371694 305504 371700 305516
rect 357400 305476 371700 305504
rect 357400 305464 357406 305476
rect 371694 305464 371700 305476
rect 371752 305464 371758 305516
rect 216214 305396 216220 305448
rect 216272 305436 216278 305448
rect 277210 305436 277216 305448
rect 216272 305408 277216 305436
rect 216272 305396 216278 305408
rect 277210 305396 277216 305408
rect 277268 305396 277274 305448
rect 351454 305396 351460 305448
rect 351512 305436 351518 305448
rect 358814 305436 358820 305448
rect 351512 305408 358820 305436
rect 351512 305396 351518 305408
rect 358814 305396 358820 305408
rect 358872 305396 358878 305448
rect 359090 305396 359096 305448
rect 359148 305436 359154 305448
rect 359734 305436 359740 305448
rect 359148 305408 359740 305436
rect 359148 305396 359154 305408
rect 359734 305396 359740 305408
rect 359792 305396 359798 305448
rect 365070 305436 365076 305448
rect 360166 305408 365076 305436
rect 234982 305328 234988 305380
rect 235040 305368 235046 305380
rect 235442 305368 235448 305380
rect 235040 305340 235448 305368
rect 235040 305328 235046 305340
rect 235442 305328 235448 305340
rect 235500 305328 235506 305380
rect 237650 305328 237656 305380
rect 237708 305368 237714 305380
rect 238294 305368 238300 305380
rect 237708 305340 238300 305368
rect 237708 305328 237714 305340
rect 238294 305328 238300 305340
rect 238352 305328 238358 305380
rect 239122 305328 239128 305380
rect 239180 305368 239186 305380
rect 240042 305368 240048 305380
rect 239180 305340 240048 305368
rect 239180 305328 239186 305340
rect 240042 305328 240048 305340
rect 240100 305328 240106 305380
rect 241790 305328 241796 305380
rect 241848 305368 241854 305380
rect 242434 305368 242440 305380
rect 241848 305340 242440 305368
rect 241848 305328 241854 305340
rect 242434 305328 242440 305340
rect 242492 305328 242498 305380
rect 253934 305328 253940 305380
rect 253992 305368 253998 305380
rect 254302 305368 254308 305380
rect 253992 305340 254308 305368
rect 253992 305328 253998 305340
rect 254302 305328 254308 305340
rect 254360 305328 254366 305380
rect 255498 305328 255504 305380
rect 255556 305368 255562 305380
rect 256418 305368 256424 305380
rect 255556 305340 256424 305368
rect 255556 305328 255562 305340
rect 256418 305328 256424 305340
rect 256476 305328 256482 305380
rect 258258 305328 258264 305380
rect 258316 305368 258322 305380
rect 259178 305368 259184 305380
rect 258316 305340 259184 305368
rect 258316 305328 258322 305340
rect 259178 305328 259184 305340
rect 259236 305328 259242 305380
rect 259730 305328 259736 305380
rect 259788 305368 259794 305380
rect 260558 305368 260564 305380
rect 259788 305340 260564 305368
rect 259788 305328 259794 305340
rect 260558 305328 260564 305340
rect 260616 305328 260622 305380
rect 260834 305328 260840 305380
rect 260892 305368 260898 305380
rect 261294 305368 261300 305380
rect 260892 305340 261300 305368
rect 260892 305328 260898 305340
rect 261294 305328 261300 305340
rect 261352 305328 261358 305380
rect 262214 305328 262220 305380
rect 262272 305368 262278 305380
rect 262582 305368 262588 305380
rect 262272 305340 262588 305368
rect 262272 305328 262278 305340
rect 262582 305328 262588 305340
rect 262640 305328 262646 305380
rect 353294 305328 353300 305380
rect 353352 305368 353358 305380
rect 360166 305368 360194 305408
rect 365070 305396 365076 305408
rect 365128 305396 365134 305448
rect 353352 305340 360194 305368
rect 353352 305328 353358 305340
rect 237742 305260 237748 305312
rect 237800 305300 237806 305312
rect 238662 305300 238668 305312
rect 237800 305272 238668 305300
rect 237800 305260 237806 305272
rect 238662 305260 238668 305272
rect 238720 305260 238726 305312
rect 259546 305260 259552 305312
rect 259604 305300 259610 305312
rect 260190 305300 260196 305312
rect 259604 305272 260196 305300
rect 259604 305260 259610 305272
rect 260190 305260 260196 305272
rect 260248 305260 260254 305312
rect 260926 305260 260932 305312
rect 260984 305300 260990 305312
rect 261938 305300 261944 305312
rect 260984 305272 261944 305300
rect 260984 305260 260990 305272
rect 261938 305260 261944 305272
rect 261996 305260 262002 305312
rect 350810 305260 350816 305312
rect 350868 305300 350874 305312
rect 358722 305300 358728 305312
rect 350868 305272 358728 305300
rect 350868 305260 350874 305272
rect 358722 305260 358728 305272
rect 358780 305260 358786 305312
rect 359458 305056 359464 305108
rect 359516 305096 359522 305108
rect 360102 305096 360108 305108
rect 359516 305068 360108 305096
rect 359516 305056 359522 305068
rect 360102 305056 360108 305068
rect 360160 305056 360166 305108
rect 335446 304648 335452 304700
rect 335504 304688 335510 304700
rect 336458 304688 336464 304700
rect 335504 304660 336464 304688
rect 335504 304648 335510 304660
rect 336458 304648 336464 304660
rect 336516 304648 336522 304700
rect 317414 304512 317420 304564
rect 317472 304552 317478 304564
rect 318334 304552 318340 304564
rect 317472 304524 318340 304552
rect 317472 304512 317478 304524
rect 318334 304512 318340 304524
rect 318392 304512 318398 304564
rect 308582 304376 308588 304428
rect 308640 304416 308646 304428
rect 390554 304416 390560 304428
rect 308640 304388 390560 304416
rect 308640 304376 308646 304388
rect 390554 304376 390560 304388
rect 390612 304376 390618 304428
rect 301038 304308 301044 304360
rect 301096 304348 301102 304360
rect 301222 304348 301228 304360
rect 301096 304320 301228 304348
rect 301096 304308 301102 304320
rect 301222 304308 301228 304320
rect 301280 304308 301286 304360
rect 314102 304308 314108 304360
rect 314160 304348 314166 304360
rect 418154 304348 418160 304360
rect 314160 304320 418160 304348
rect 314160 304308 314166 304320
rect 418154 304308 418160 304320
rect 418212 304308 418218 304360
rect 217410 304240 217416 304292
rect 217468 304280 217474 304292
rect 352650 304280 352656 304292
rect 217468 304252 352656 304280
rect 217468 304240 217474 304252
rect 352650 304240 352656 304252
rect 352708 304240 352714 304292
rect 317598 304172 317604 304224
rect 317656 304212 317662 304224
rect 317874 304212 317880 304224
rect 317656 304184 317880 304212
rect 317656 304172 317662 304184
rect 317874 304172 317880 304184
rect 317932 304172 317938 304224
rect 322934 304172 322940 304224
rect 322992 304212 322998 304224
rect 323302 304212 323308 304224
rect 322992 304184 323308 304212
rect 322992 304172 322998 304184
rect 323302 304172 323308 304184
rect 323360 304172 323366 304224
rect 324590 304172 324596 304224
rect 324648 304212 324654 304224
rect 325602 304212 325608 304224
rect 324648 304184 325608 304212
rect 324648 304172 324654 304184
rect 325602 304172 325608 304184
rect 325660 304172 325666 304224
rect 255314 304104 255320 304156
rect 255372 304144 255378 304156
rect 255682 304144 255688 304156
rect 255372 304116 255688 304144
rect 255372 304104 255378 304116
rect 255682 304104 255688 304116
rect 255740 304104 255746 304156
rect 258074 303696 258080 303748
rect 258132 303736 258138 303748
rect 258350 303736 258356 303748
rect 258132 303708 258356 303736
rect 258132 303696 258138 303708
rect 258350 303696 258356 303708
rect 258408 303696 258414 303748
rect 320266 303696 320272 303748
rect 320324 303736 320330 303748
rect 320634 303736 320640 303748
rect 320324 303708 320640 303736
rect 320324 303696 320330 303708
rect 320634 303696 320640 303708
rect 320692 303696 320698 303748
rect 212442 303560 212448 303612
rect 212500 303600 212506 303612
rect 280154 303600 280160 303612
rect 212500 303572 280160 303600
rect 212500 303560 212506 303572
rect 280154 303560 280160 303572
rect 280212 303560 280218 303612
rect 353570 303560 353576 303612
rect 353628 303600 353634 303612
rect 372798 303600 372804 303612
rect 353628 303572 372804 303600
rect 353628 303560 353634 303572
rect 372798 303560 372804 303572
rect 372856 303560 372862 303612
rect 213546 303492 213552 303544
rect 213604 303532 213610 303544
rect 282086 303532 282092 303544
rect 213604 303504 282092 303532
rect 213604 303492 213610 303504
rect 282086 303492 282092 303504
rect 282144 303492 282150 303544
rect 352374 303492 352380 303544
rect 352432 303532 352438 303544
rect 372890 303532 372896 303544
rect 352432 303504 372896 303532
rect 352432 303492 352438 303504
rect 372890 303492 372896 303504
rect 372948 303492 372954 303544
rect 213086 303424 213092 303476
rect 213144 303464 213150 303476
rect 282546 303464 282552 303476
rect 213144 303436 282552 303464
rect 213144 303424 213150 303436
rect 282546 303424 282552 303436
rect 282604 303424 282610 303476
rect 351730 303424 351736 303476
rect 351788 303464 351794 303476
rect 371602 303464 371608 303476
rect 351788 303436 371608 303464
rect 351788 303424 351794 303436
rect 371602 303424 371608 303436
rect 371660 303424 371666 303476
rect 217962 303356 217968 303408
rect 218020 303396 218026 303408
rect 288250 303396 288256 303408
rect 218020 303368 288256 303396
rect 218020 303356 218026 303368
rect 288250 303356 288256 303368
rect 288308 303356 288314 303408
rect 347590 303356 347596 303408
rect 347648 303396 347654 303408
rect 371970 303396 371976 303408
rect 347648 303368 371976 303396
rect 347648 303356 347654 303368
rect 371970 303356 371976 303368
rect 372028 303356 372034 303408
rect 213638 303288 213644 303340
rect 213696 303328 213702 303340
rect 283098 303328 283104 303340
rect 213696 303300 283104 303328
rect 213696 303288 213702 303300
rect 283098 303288 283104 303300
rect 283156 303288 283162 303340
rect 306650 303288 306656 303340
rect 306708 303328 306714 303340
rect 379514 303328 379520 303340
rect 306708 303300 379520 303328
rect 306708 303288 306714 303300
rect 379514 303288 379520 303300
rect 379572 303288 379578 303340
rect 211062 303220 211068 303272
rect 211120 303260 211126 303272
rect 282270 303260 282276 303272
rect 211120 303232 282276 303260
rect 211120 303220 211126 303232
rect 282270 303220 282276 303232
rect 282328 303220 282334 303272
rect 307202 303220 307208 303272
rect 307260 303260 307266 303272
rect 382274 303260 382280 303272
rect 307260 303232 382280 303260
rect 307260 303220 307266 303232
rect 382274 303220 382280 303232
rect 382332 303220 382338 303272
rect 212350 303152 212356 303204
rect 212408 303192 212414 303204
rect 283006 303192 283012 303204
rect 212408 303164 283012 303192
rect 212408 303152 212414 303164
rect 283006 303152 283012 303164
rect 283064 303152 283070 303204
rect 301038 303152 301044 303204
rect 301096 303192 301102 303204
rect 301866 303192 301872 303204
rect 301096 303164 301872 303192
rect 301096 303152 301102 303164
rect 301866 303152 301872 303164
rect 301924 303152 301930 303204
rect 308030 303152 308036 303204
rect 308088 303192 308094 303204
rect 386414 303192 386420 303204
rect 308088 303164 386420 303192
rect 308088 303152 308094 303164
rect 386414 303152 386420 303164
rect 386472 303152 386478 303204
rect 213362 303084 213368 303136
rect 213420 303124 213426 303136
rect 346854 303124 346860 303136
rect 213420 303096 346860 303124
rect 213420 303084 213426 303096
rect 346854 303084 346860 303096
rect 346912 303084 346918 303136
rect 348510 303084 348516 303136
rect 348568 303124 348574 303136
rect 370682 303124 370688 303136
rect 348568 303096 370688 303124
rect 348568 303084 348574 303096
rect 370682 303084 370688 303096
rect 370740 303084 370746 303136
rect 306558 303016 306564 303068
rect 306616 303056 306622 303068
rect 307386 303056 307392 303068
rect 306616 303028 307392 303056
rect 306616 303016 306622 303028
rect 307386 303016 307392 303028
rect 307444 303016 307450 303068
rect 353110 303016 353116 303068
rect 353168 303056 353174 303068
rect 374270 303056 374276 303068
rect 353168 303028 374276 303056
rect 353168 303016 353174 303028
rect 374270 303016 374276 303028
rect 374328 303016 374334 303068
rect 211890 302948 211896 303000
rect 211948 302988 211954 303000
rect 347774 302988 347780 303000
rect 211948 302960 347780 302988
rect 211948 302948 211954 302960
rect 347774 302948 347780 302960
rect 347832 302948 347838 303000
rect 349614 302948 349620 303000
rect 349672 302988 349678 303000
rect 372706 302988 372712 303000
rect 349672 302960 372712 302988
rect 349672 302948 349678 302960
rect 372706 302948 372712 302960
rect 372764 302948 372770 303000
rect 210602 302880 210608 302932
rect 210660 302920 210666 302932
rect 348050 302920 348056 302932
rect 210660 302892 348056 302920
rect 210660 302880 210666 302892
rect 348050 302880 348056 302892
rect 348108 302880 348114 302932
rect 348694 302880 348700 302932
rect 348752 302920 348758 302932
rect 374178 302920 374184 302932
rect 348752 302892 374184 302920
rect 348752 302880 348758 302892
rect 374178 302880 374184 302892
rect 374236 302880 374242 302932
rect 217870 302812 217876 302864
rect 217928 302852 217934 302864
rect 283926 302852 283932 302864
rect 217928 302824 283932 302852
rect 217928 302812 217934 302824
rect 283926 302812 283932 302824
rect 283984 302812 283990 302864
rect 349430 302812 349436 302864
rect 349488 302852 349494 302864
rect 367646 302852 367652 302864
rect 349488 302824 367652 302852
rect 349488 302812 349494 302824
rect 367646 302812 367652 302824
rect 367704 302812 367710 302864
rect 215938 302744 215944 302796
rect 215996 302784 216002 302796
rect 280890 302784 280896 302796
rect 215996 302756 280896 302784
rect 215996 302744 216002 302756
rect 280890 302744 280896 302756
rect 280948 302744 280954 302796
rect 350350 302744 350356 302796
rect 350408 302784 350414 302796
rect 366542 302784 366548 302796
rect 350408 302756 366548 302784
rect 350408 302744 350414 302756
rect 366542 302744 366548 302756
rect 366600 302744 366606 302796
rect 218790 302676 218796 302728
rect 218848 302716 218854 302728
rect 281534 302716 281540 302728
rect 218848 302688 281540 302716
rect 218848 302676 218854 302688
rect 281534 302676 281540 302688
rect 281592 302676 281598 302728
rect 356330 302676 356336 302728
rect 356388 302716 356394 302728
rect 370590 302716 370596 302728
rect 356388 302688 370596 302716
rect 356388 302676 356394 302688
rect 370590 302676 370596 302688
rect 370648 302676 370654 302728
rect 217502 302608 217508 302660
rect 217560 302648 217566 302660
rect 351914 302648 351920 302660
rect 217560 302620 351920 302648
rect 217560 302608 217566 302620
rect 351914 302608 351920 302620
rect 351972 302608 351978 302660
rect 305270 302336 305276 302388
rect 305328 302376 305334 302388
rect 305546 302376 305552 302388
rect 305328 302348 305552 302376
rect 305328 302336 305334 302348
rect 305546 302336 305552 302348
rect 305604 302336 305610 302388
rect 305638 301792 305644 301844
rect 305696 301832 305702 301844
rect 375374 301832 375380 301844
rect 305696 301804 375380 301832
rect 305696 301792 305702 301804
rect 375374 301792 375380 301804
rect 375432 301792 375438 301844
rect 217594 301724 217600 301776
rect 217652 301764 217658 301776
rect 345014 301764 345020 301776
rect 217652 301736 345020 301764
rect 217652 301724 217658 301736
rect 345014 301724 345020 301736
rect 345072 301724 345078 301776
rect 217042 301656 217048 301708
rect 217100 301696 217106 301708
rect 350626 301696 350632 301708
rect 217100 301668 350632 301696
rect 217100 301656 217106 301668
rect 350626 301656 350632 301668
rect 350684 301656 350690 301708
rect 341610 301588 341616 301640
rect 341668 301628 341674 301640
rect 560294 301628 560300 301640
rect 341668 301600 560300 301628
rect 341668 301588 341674 301600
rect 560294 301588 560300 301600
rect 560352 301588 560358 301640
rect 342806 301520 342812 301572
rect 342864 301560 342870 301572
rect 564434 301560 564440 301572
rect 342864 301532 564440 301560
rect 342864 301520 342870 301532
rect 564434 301520 564440 301532
rect 564492 301520 564498 301572
rect 344370 301452 344376 301504
rect 344428 301492 344434 301504
rect 574094 301492 574100 301504
rect 344428 301464 574100 301492
rect 344428 301452 344434 301464
rect 574094 301452 574100 301464
rect 574152 301452 574158 301504
rect 243170 300840 243176 300892
rect 243228 300880 243234 300892
rect 243354 300880 243360 300892
rect 243228 300852 243360 300880
rect 243228 300840 243234 300852
rect 243354 300840 243360 300852
rect 243412 300840 243418 300892
rect 216030 300772 216036 300824
rect 216088 300812 216094 300824
rect 285858 300812 285864 300824
rect 216088 300784 285864 300812
rect 216088 300772 216094 300784
rect 285858 300772 285864 300784
rect 285916 300772 285922 300824
rect 214374 300704 214380 300756
rect 214432 300744 214438 300756
rect 285766 300744 285772 300756
rect 214432 300716 285772 300744
rect 214432 300704 214438 300716
rect 285766 300704 285772 300716
rect 285824 300704 285830 300756
rect 212166 300636 212172 300688
rect 212224 300676 212230 300688
rect 284294 300676 284300 300688
rect 212224 300648 284300 300676
rect 212224 300636 212230 300648
rect 284294 300636 284300 300648
rect 284352 300636 284358 300688
rect 213178 300568 213184 300620
rect 213236 300608 213242 300620
rect 280982 300608 280988 300620
rect 213236 300580 280988 300608
rect 213236 300568 213242 300580
rect 280982 300568 280988 300580
rect 281040 300568 281046 300620
rect 210970 300500 210976 300552
rect 211028 300540 211034 300552
rect 284386 300540 284392 300552
rect 211028 300512 284392 300540
rect 211028 300500 211034 300512
rect 284386 300500 284392 300512
rect 284444 300500 284450 300552
rect 210878 300432 210884 300484
rect 210936 300472 210942 300484
rect 284754 300472 284760 300484
rect 210936 300444 284760 300472
rect 210936 300432 210942 300444
rect 284754 300432 284760 300444
rect 284812 300432 284818 300484
rect 305362 300432 305368 300484
rect 305420 300472 305426 300484
rect 372614 300472 372620 300484
rect 305420 300444 372620 300472
rect 305420 300432 305426 300444
rect 372614 300432 372620 300444
rect 372672 300432 372678 300484
rect 212258 300364 212264 300416
rect 212316 300404 212322 300416
rect 285674 300404 285680 300416
rect 212316 300376 285680 300404
rect 212316 300364 212322 300376
rect 285674 300364 285680 300376
rect 285732 300364 285738 300416
rect 321922 300364 321928 300416
rect 321980 300404 321986 300416
rect 456794 300404 456800 300416
rect 321980 300376 456800 300404
rect 321980 300364 321986 300376
rect 456794 300364 456800 300376
rect 456852 300364 456858 300416
rect 210510 300296 210516 300348
rect 210568 300336 210574 300348
rect 350534 300336 350540 300348
rect 210568 300308 350540 300336
rect 210568 300296 210574 300308
rect 350534 300296 350540 300308
rect 350592 300296 350598 300348
rect 210694 300228 210700 300280
rect 210752 300268 210758 300280
rect 284662 300268 284668 300280
rect 210752 300240 284668 300268
rect 210752 300228 210758 300240
rect 284662 300228 284668 300240
rect 284720 300228 284726 300280
rect 338574 300228 338580 300280
rect 338632 300268 338638 300280
rect 542354 300268 542360 300280
rect 338632 300240 542360 300268
rect 338632 300228 338638 300240
rect 542354 300228 542360 300240
rect 542412 300228 542418 300280
rect 210786 300160 210792 300212
rect 210844 300200 210850 300212
rect 284478 300200 284484 300212
rect 210844 300172 284484 300200
rect 210844 300160 210850 300172
rect 284478 300160 284484 300172
rect 284536 300160 284542 300212
rect 339770 300160 339776 300212
rect 339828 300200 339834 300212
rect 549254 300200 549260 300212
rect 339828 300172 549260 300200
rect 339828 300160 339834 300172
rect 549254 300160 549260 300172
rect 549312 300160 549318 300212
rect 213454 300092 213460 300144
rect 213512 300132 213518 300144
rect 288434 300132 288440 300144
rect 213512 300104 288440 300132
rect 213512 300092 213518 300104
rect 288434 300092 288440 300104
rect 288492 300092 288498 300144
rect 340230 300092 340236 300144
rect 340288 300132 340294 300144
rect 553394 300132 553400 300144
rect 340288 300104 553400 300132
rect 340288 300092 340294 300104
rect 553394 300092 553400 300104
rect 553452 300092 553458 300144
rect 215846 300024 215852 300076
rect 215904 300064 215910 300076
rect 286410 300064 286416 300076
rect 215904 300036 286416 300064
rect 215904 300024 215910 300036
rect 286410 300024 286416 300036
rect 286468 300024 286474 300076
rect 217778 299956 217784 300008
rect 217836 299996 217842 300008
rect 283282 299996 283288 300008
rect 217836 299968 283288 299996
rect 217836 299956 217842 299968
rect 283282 299956 283288 299968
rect 283340 299956 283346 300008
rect 219342 299888 219348 299940
rect 219400 299928 219406 299940
rect 284570 299928 284576 299940
rect 219400 299900 284576 299928
rect 219400 299888 219406 299900
rect 284570 299888 284576 299900
rect 284628 299888 284634 299940
rect 321002 298936 321008 298988
rect 321060 298976 321066 298988
rect 454034 298976 454040 298988
rect 321060 298948 454040 298976
rect 321060 298936 321066 298948
rect 454034 298936 454040 298948
rect 454092 298936 454098 298988
rect 336090 298868 336096 298920
rect 336148 298908 336154 298920
rect 531314 298908 531320 298920
rect 336148 298880 531320 298908
rect 336148 298868 336154 298880
rect 531314 298868 531320 298880
rect 531372 298868 531378 298920
rect 337194 298800 337200 298852
rect 337252 298840 337258 298852
rect 535454 298840 535460 298852
rect 337252 298812 535460 298840
rect 337252 298800 337258 298812
rect 535454 298800 535460 298812
rect 535512 298800 535518 298852
rect 337102 298732 337108 298784
rect 337160 298772 337166 298784
rect 539594 298772 539600 298784
rect 337160 298744 539600 298772
rect 337160 298732 337166 298744
rect 539594 298732 539600 298744
rect 539652 298732 539658 298784
rect 330662 297576 330668 297628
rect 330720 297616 330726 297628
rect 503714 297616 503720 297628
rect 330720 297588 503720 297616
rect 330720 297576 330726 297588
rect 503714 297576 503720 297588
rect 503772 297576 503778 297628
rect 331674 297508 331680 297560
rect 331732 297548 331738 297560
rect 506474 297548 506480 297560
rect 331732 297520 506480 297548
rect 331732 297508 331738 297520
rect 506474 297508 506480 297520
rect 506532 297508 506538 297560
rect 331582 297440 331588 297492
rect 331640 297480 331646 297492
rect 510614 297480 510620 297492
rect 331640 297452 510620 297480
rect 331640 297440 331646 297452
rect 510614 297440 510620 297452
rect 510672 297440 510678 297492
rect 342622 297372 342628 297424
rect 342680 297412 342686 297424
rect 567194 297412 567200 297424
rect 342680 297384 567200 297412
rect 342680 297372 342686 297384
rect 567194 297372 567200 297384
rect 567252 297372 567258 297424
rect 218606 296216 218612 296268
rect 218664 296256 218670 296268
rect 349154 296256 349160 296268
rect 218664 296228 349160 296256
rect 218664 296216 218670 296228
rect 349154 296216 349160 296228
rect 349212 296216 349218 296268
rect 327534 296148 327540 296200
rect 327592 296188 327598 296200
rect 489914 296188 489920 296200
rect 327592 296160 489920 296188
rect 327592 296148 327598 296160
rect 489914 296148 489920 296160
rect 489972 296148 489978 296200
rect 328914 296080 328920 296132
rect 328972 296120 328978 296132
rect 492674 296120 492680 296132
rect 328972 296092 492680 296120
rect 328972 296080 328978 296092
rect 492674 296080 492680 296092
rect 492732 296080 492738 296132
rect 330110 296012 330116 296064
rect 330168 296052 330174 296064
rect 499574 296052 499580 296064
rect 330168 296024 499580 296052
rect 330168 296012 330174 296024
rect 499574 296012 499580 296024
rect 499632 296012 499638 296064
rect 341242 295944 341248 295996
rect 341300 295984 341306 295996
rect 556154 295984 556160 295996
rect 341300 295956 556160 295984
rect 341300 295944 341306 295956
rect 556154 295944 556160 295956
rect 556212 295944 556218 295996
rect 218514 294856 218520 294908
rect 218572 294896 218578 294908
rect 348234 294896 348240 294908
rect 218572 294868 348240 294896
rect 218572 294856 218578 294868
rect 348234 294856 348240 294868
rect 348292 294856 348298 294908
rect 321830 294788 321836 294840
rect 321888 294828 321894 294840
rect 463694 294828 463700 294840
rect 321888 294800 463700 294828
rect 321888 294788 321894 294800
rect 463694 294788 463700 294800
rect 463752 294788 463758 294840
rect 324682 294720 324688 294772
rect 324740 294760 324746 294772
rect 473354 294760 473360 294772
rect 324740 294732 473360 294760
rect 324740 294720 324746 294732
rect 473354 294720 473360 294732
rect 473412 294720 473418 294772
rect 326062 294652 326068 294704
rect 326120 294692 326126 294704
rect 481634 294692 481640 294704
rect 326120 294664 481640 294692
rect 326120 294652 326126 294664
rect 481634 294652 481640 294664
rect 481692 294652 481698 294704
rect 124214 294584 124220 294636
rect 124272 294624 124278 294636
rect 256694 294624 256700 294636
rect 124272 294596 256700 294624
rect 124272 294584 124278 294596
rect 256694 294584 256700 294596
rect 256752 294584 256758 294636
rect 335722 294584 335728 294636
rect 335780 294624 335786 294636
rect 528554 294624 528560 294636
rect 335780 294596 528560 294624
rect 335780 294584 335786 294596
rect 528554 294584 528560 294596
rect 528612 294584 528618 294636
rect 314930 293428 314936 293480
rect 314988 293468 314994 293480
rect 427814 293468 427820 293480
rect 314988 293440 427820 293468
rect 314988 293428 314994 293440
rect 427814 293428 427820 293440
rect 427872 293428 427878 293480
rect 117314 293360 117320 293412
rect 117372 293400 117378 293412
rect 255682 293400 255688 293412
rect 117372 293372 255688 293400
rect 117372 293360 117378 293372
rect 255682 293360 255688 293372
rect 255740 293360 255746 293412
rect 317874 293360 317880 293412
rect 317932 293400 317938 293412
rect 441614 293400 441620 293412
rect 317932 293372 441620 293400
rect 317932 293360 317938 293372
rect 441614 293360 441620 293372
rect 441672 293360 441678 293412
rect 110414 293292 110420 293344
rect 110472 293332 110478 293344
rect 254302 293332 254308 293344
rect 110472 293304 254308 293332
rect 110472 293292 110478 293304
rect 254302 293292 254308 293304
rect 254360 293292 254366 293344
rect 321738 293292 321744 293344
rect 321796 293332 321802 293344
rect 459554 293332 459560 293344
rect 321796 293304 459560 293332
rect 321796 293292 321802 293304
rect 459554 293292 459560 293304
rect 459612 293292 459618 293344
rect 102134 293224 102140 293276
rect 102192 293264 102198 293276
rect 252922 293264 252928 293276
rect 102192 293236 252928 293264
rect 102192 293224 102198 293236
rect 252922 293224 252928 293236
rect 252980 293224 252986 293276
rect 324590 293224 324596 293276
rect 324648 293264 324654 293276
rect 477494 293264 477500 293276
rect 324648 293236 477500 293264
rect 324648 293224 324654 293236
rect 477494 293224 477500 293236
rect 477552 293224 477558 293276
rect 112438 292000 112444 292052
rect 112496 292040 112502 292052
rect 251174 292040 251180 292052
rect 112496 292012 251180 292040
rect 112496 292000 112502 292012
rect 251174 292000 251180 292012
rect 251232 292000 251238 292052
rect 312078 292000 312084 292052
rect 312136 292040 312142 292052
rect 409874 292040 409880 292052
rect 312136 292012 409880 292040
rect 312136 292000 312142 292012
rect 409874 292000 409880 292012
rect 409932 292000 409938 292052
rect 92474 291932 92480 291984
rect 92532 291972 92538 291984
rect 250162 291972 250168 291984
rect 92532 291944 250168 291972
rect 92532 291932 92538 291944
rect 250162 291932 250168 291944
rect 250220 291932 250226 291984
rect 312170 291932 312176 291984
rect 312228 291972 312234 291984
rect 414014 291972 414020 291984
rect 312228 291944 414020 291972
rect 312228 291932 312234 291944
rect 414014 291932 414020 291944
rect 414072 291932 414078 291984
rect 88334 291864 88340 291916
rect 88392 291904 88398 291916
rect 249794 291904 249800 291916
rect 88392 291876 249800 291904
rect 88392 291864 88398 291876
rect 249794 291864 249800 291876
rect 249852 291864 249858 291916
rect 314838 291864 314844 291916
rect 314896 291904 314902 291916
rect 423674 291904 423680 291916
rect 314896 291876 423680 291904
rect 314896 291864 314902 291876
rect 423674 291864 423680 291876
rect 423732 291864 423738 291916
rect 85574 291796 85580 291848
rect 85632 291836 85638 291848
rect 248782 291836 248788 291848
rect 85632 291808 248788 291836
rect 85632 291796 85638 291808
rect 248782 291796 248788 291808
rect 248840 291796 248846 291848
rect 316310 291796 316316 291848
rect 316368 291836 316374 291848
rect 434714 291836 434720 291848
rect 316368 291808 434720 291836
rect 316368 291796 316374 291808
rect 434714 291796 434720 291808
rect 434772 291796 434778 291848
rect 104158 290640 104164 290692
rect 104216 290680 104222 290692
rect 247494 290680 247500 290692
rect 104216 290652 247500 290680
rect 104216 290640 104222 290652
rect 247494 290640 247500 290652
rect 247552 290640 247558 290692
rect 309410 290640 309416 290692
rect 309468 290680 309474 290692
rect 398834 290680 398840 290692
rect 309468 290652 398840 290680
rect 309468 290640 309474 290652
rect 398834 290640 398840 290652
rect 398892 290640 398898 290692
rect 77294 290572 77300 290624
rect 77352 290612 77358 290624
rect 247402 290612 247408 290624
rect 77352 290584 247408 290612
rect 77352 290572 77358 290584
rect 247402 290572 247408 290584
rect 247460 290572 247466 290624
rect 310698 290572 310704 290624
rect 310756 290612 310762 290624
rect 402974 290612 402980 290624
rect 310756 290584 402980 290612
rect 310756 290572 310762 290584
rect 402974 290572 402980 290584
rect 403032 290572 403038 290624
rect 74534 290504 74540 290556
rect 74592 290544 74598 290556
rect 246022 290544 246028 290556
rect 74592 290516 246028 290544
rect 74592 290504 74598 290516
rect 246022 290504 246028 290516
rect 246080 290504 246086 290556
rect 310790 290504 310796 290556
rect 310848 290544 310854 290556
rect 407206 290544 407212 290556
rect 310848 290516 407212 290544
rect 310848 290504 310854 290516
rect 407206 290504 407212 290516
rect 407264 290504 407270 290556
rect 70394 290436 70400 290488
rect 70452 290476 70458 290488
rect 246114 290476 246120 290488
rect 70452 290448 246120 290476
rect 70452 290436 70458 290448
rect 246114 290436 246120 290448
rect 246172 290436 246178 290488
rect 313642 290436 313648 290488
rect 313700 290476 313706 290488
rect 420914 290476 420920 290488
rect 313700 290448 420920 290476
rect 313700 290436 313706 290448
rect 420914 290436 420920 290448
rect 420972 290436 420978 290488
rect 122834 289280 122840 289332
rect 122892 289320 122898 289332
rect 255498 289320 255504 289332
rect 122892 289292 255504 289320
rect 122892 289280 122898 289292
rect 255498 289280 255504 289292
rect 255556 289280 255562 289332
rect 306650 289280 306656 289332
rect 306708 289320 306714 289332
rect 382366 289320 382372 289332
rect 306708 289292 382372 289320
rect 306708 289280 306714 289292
rect 382366 289280 382372 289292
rect 382424 289280 382430 289332
rect 118694 289212 118700 289264
rect 118752 289252 118758 289264
rect 255590 289252 255596 289264
rect 118752 289224 255596 289252
rect 118752 289212 118758 289224
rect 255590 289212 255596 289224
rect 255648 289212 255654 289264
rect 308030 289212 308036 289264
rect 308088 289252 308094 289264
rect 391934 289252 391940 289264
rect 308088 289224 391940 289252
rect 308088 289212 308094 289224
rect 391934 289212 391940 289224
rect 391992 289212 391998 289264
rect 115934 289144 115940 289196
rect 115992 289184 115998 289196
rect 254210 289184 254216 289196
rect 115992 289156 254216 289184
rect 115992 289144 115998 289156
rect 254210 289144 254216 289156
rect 254268 289144 254274 289196
rect 309318 289144 309324 289196
rect 309376 289184 309382 289196
rect 396074 289184 396080 289196
rect 309376 289156 396080 289184
rect 309376 289144 309382 289156
rect 396074 289144 396080 289156
rect 396132 289144 396138 289196
rect 63494 289076 63500 289128
rect 63552 289116 63558 289128
rect 244642 289116 244648 289128
rect 63552 289088 244648 289116
rect 63552 289076 63558 289088
rect 244642 289076 244648 289088
rect 244700 289076 244706 289128
rect 323302 289076 323308 289128
rect 323360 289116 323366 289128
rect 470594 289116 470600 289128
rect 323360 289088 470600 289116
rect 323360 289076 323366 289088
rect 470594 289076 470600 289088
rect 470652 289076 470658 289128
rect 111794 287852 111800 287904
rect 111852 287892 111858 287904
rect 254118 287892 254124 287904
rect 111852 287864 254124 287892
rect 111852 287852 111858 287864
rect 254118 287852 254124 287864
rect 254176 287852 254182 287904
rect 303982 287852 303988 287904
rect 304040 287892 304046 287904
rect 371234 287892 371240 287904
rect 304040 287864 371240 287892
rect 304040 287852 304046 287864
rect 371234 287852 371240 287864
rect 371292 287852 371298 287904
rect 109034 287784 109040 287836
rect 109092 287824 109098 287836
rect 252830 287824 252836 287836
rect 109092 287796 252836 287824
rect 109092 287784 109098 287796
rect 252830 287784 252836 287796
rect 252888 287784 252894 287836
rect 305270 287784 305276 287836
rect 305328 287824 305334 287836
rect 373994 287824 374000 287836
rect 305328 287796 374000 287824
rect 305328 287784 305334 287796
rect 373994 287784 374000 287796
rect 374052 287784 374058 287836
rect 104894 287716 104900 287768
rect 104952 287756 104958 287768
rect 252738 287756 252744 287768
rect 104952 287728 252744 287756
rect 104952 287716 104958 287728
rect 252738 287716 252744 287728
rect 252796 287716 252802 287768
rect 305178 287716 305184 287768
rect 305236 287756 305242 287768
rect 378134 287756 378140 287768
rect 305236 287728 378140 287756
rect 305236 287716 305242 287728
rect 378134 287716 378140 287728
rect 378192 287716 378198 287768
rect 52454 287648 52460 287700
rect 52512 287688 52518 287700
rect 241974 287688 241980 287700
rect 52512 287660 241980 287688
rect 52512 287648 52518 287660
rect 241974 287648 241980 287660
rect 242032 287648 242038 287700
rect 319254 287648 319260 287700
rect 319312 287688 319318 287700
rect 445754 287688 445760 287700
rect 319312 287660 445760 287688
rect 319312 287648 319318 287660
rect 445754 287648 445760 287660
rect 445812 287648 445818 287700
rect 102226 286492 102232 286544
rect 102284 286532 102290 286544
rect 251542 286532 251548 286544
rect 102284 286504 251548 286532
rect 102284 286492 102290 286504
rect 251542 286492 251548 286504
rect 251600 286492 251606 286544
rect 319162 286492 319168 286544
rect 319220 286532 319226 286544
rect 447134 286532 447140 286544
rect 319220 286504 447140 286532
rect 319220 286492 319226 286504
rect 447134 286492 447140 286504
rect 447192 286492 447198 286544
rect 97994 286424 98000 286476
rect 98052 286464 98058 286476
rect 251450 286464 251456 286476
rect 98052 286436 251456 286464
rect 98052 286424 98058 286436
rect 251450 286424 251456 286436
rect 251508 286424 251514 286476
rect 344002 286424 344008 286476
rect 344060 286464 344066 286476
rect 542998 286464 543004 286476
rect 344060 286436 543004 286464
rect 344060 286424 344066 286436
rect 542998 286424 543004 286436
rect 543056 286424 543062 286476
rect 91094 286356 91100 286408
rect 91152 286396 91158 286408
rect 250070 286396 250076 286408
rect 91152 286368 250076 286396
rect 91152 286356 91158 286368
rect 250070 286356 250076 286368
rect 250128 286356 250134 286408
rect 345198 286356 345204 286408
rect 345256 286396 345262 286408
rect 552658 286396 552664 286408
rect 345256 286368 552664 286396
rect 345256 286356 345262 286368
rect 552658 286356 552664 286368
rect 552716 286356 552722 286408
rect 49694 286288 49700 286340
rect 49752 286328 49758 286340
rect 241882 286328 241888 286340
rect 49752 286300 241888 286328
rect 49752 286288 49758 286300
rect 241882 286288 241888 286300
rect 241940 286288 241946 286340
rect 343910 286288 343916 286340
rect 343968 286328 343974 286340
rect 569954 286328 569960 286340
rect 343968 286300 569960 286328
rect 343968 286288 343974 286300
rect 569954 286288 569960 286300
rect 570012 286288 570018 286340
rect 114554 285200 114560 285252
rect 114612 285240 114618 285252
rect 254026 285240 254032 285252
rect 114612 285212 254032 285240
rect 114612 285200 114618 285212
rect 254026 285200 254032 285212
rect 254084 285200 254090 285252
rect 93854 285132 93860 285184
rect 93912 285172 93918 285184
rect 249978 285172 249984 285184
rect 93912 285144 249984 285172
rect 93912 285132 93918 285144
rect 249978 285132 249984 285144
rect 250036 285132 250042 285184
rect 327442 285132 327448 285184
rect 327500 285172 327506 285184
rect 485774 285172 485780 285184
rect 327500 285144 485780 285172
rect 327500 285132 327506 285144
rect 485774 285132 485780 285144
rect 485832 285132 485838 285184
rect 86954 285064 86960 285116
rect 87012 285104 87018 285116
rect 248690 285104 248696 285116
rect 87012 285076 248696 285104
rect 87012 285064 87018 285076
rect 248690 285064 248696 285076
rect 248748 285064 248754 285116
rect 341150 285064 341156 285116
rect 341208 285104 341214 285116
rect 538858 285104 538864 285116
rect 341208 285076 538864 285104
rect 341208 285064 341214 285076
rect 538858 285064 538864 285076
rect 538916 285064 538922 285116
rect 77386 284996 77392 285048
rect 77444 285036 77450 285048
rect 247310 285036 247316 285048
rect 77444 285008 247316 285036
rect 77444 284996 77450 285008
rect 247310 284996 247316 285008
rect 247368 284996 247374 285048
rect 342438 284996 342444 285048
rect 342496 285036 342502 285048
rect 563054 285036 563060 285048
rect 342496 285008 563060 285036
rect 342496 284996 342502 285008
rect 563054 284996 563060 285008
rect 563112 284996 563118 285048
rect 38654 284928 38660 284980
rect 38712 284968 38718 284980
rect 239122 284968 239128 284980
rect 38712 284940 239128 284968
rect 38712 284928 38718 284940
rect 239122 284928 239128 284940
rect 239180 284928 239186 284980
rect 342530 284928 342536 284980
rect 342588 284968 342594 284980
rect 565814 284968 565820 284980
rect 342588 284940 565820 284968
rect 342588 284928 342594 284940
rect 565814 284928 565820 284940
rect 565872 284928 565878 284980
rect 110506 283840 110512 283892
rect 110564 283880 110570 283892
rect 254394 283880 254400 283892
rect 110564 283852 254400 283880
rect 110564 283840 110570 283852
rect 254394 283840 254400 283852
rect 254452 283840 254458 283892
rect 107654 283772 107660 283824
rect 107712 283812 107718 283824
rect 252646 283812 252652 283824
rect 107712 283784 252652 283812
rect 107712 283772 107718 283784
rect 252646 283772 252652 283784
rect 252704 283772 252710 283824
rect 316218 283772 316224 283824
rect 316276 283812 316282 283824
rect 431954 283812 431960 283824
rect 316276 283784 431960 283812
rect 316276 283772 316282 283784
rect 431954 283772 431960 283784
rect 432012 283772 432018 283824
rect 100754 283704 100760 283756
rect 100812 283744 100818 283756
rect 251358 283744 251364 283756
rect 100812 283716 251364 283744
rect 100812 283704 100818 283716
rect 251358 283704 251364 283716
rect 251416 283704 251422 283756
rect 335630 283704 335636 283756
rect 335688 283744 335694 283756
rect 531406 283744 531412 283756
rect 335688 283716 531412 283744
rect 335688 283704 335694 283716
rect 531406 283704 531412 283716
rect 531464 283704 531470 283756
rect 73154 283636 73160 283688
rect 73212 283676 73218 283688
rect 245930 283676 245936 283688
rect 73212 283648 245936 283676
rect 73212 283636 73218 283648
rect 245930 283636 245936 283648
rect 245988 283636 245994 283688
rect 339678 283636 339684 283688
rect 339736 283676 339742 283688
rect 547874 283676 547880 283688
rect 339736 283648 547880 283676
rect 339736 283636 339742 283648
rect 547874 283636 547880 283648
rect 547932 283636 547938 283688
rect 43530 283568 43536 283620
rect 43588 283608 43594 283620
rect 240502 283608 240508 283620
rect 43588 283580 240508 283608
rect 43588 283568 43594 283580
rect 240502 283568 240508 283580
rect 240560 283568 240566 283620
rect 339770 283568 339776 283620
rect 339828 283608 339834 283620
rect 552014 283608 552020 283620
rect 339828 283580 552020 283608
rect 339828 283568 339834 283580
rect 552014 283568 552020 283580
rect 552072 283568 552078 283620
rect 160094 282412 160100 282464
rect 160152 282452 160158 282464
rect 264054 282452 264060 282464
rect 160152 282424 264060 282452
rect 160152 282412 160158 282424
rect 264054 282412 264060 282424
rect 264112 282412 264118 282464
rect 103514 282344 103520 282396
rect 103572 282384 103578 282396
rect 253014 282384 253020 282396
rect 103572 282356 253020 282384
rect 103572 282344 103578 282356
rect 253014 282344 253020 282356
rect 253072 282344 253078 282396
rect 313550 282344 313556 282396
rect 313608 282384 313614 282396
rect 416774 282384 416780 282396
rect 313608 282356 416780 282384
rect 313608 282344 313614 282356
rect 416774 282344 416780 282356
rect 416832 282344 416838 282396
rect 96614 282276 96620 282328
rect 96672 282316 96678 282328
rect 251266 282316 251272 282328
rect 96672 282288 251272 282316
rect 96672 282276 96678 282288
rect 251266 282276 251272 282288
rect 251324 282276 251330 282328
rect 333054 282276 333060 282328
rect 333112 282316 333118 282328
rect 516134 282316 516140 282328
rect 333112 282288 516140 282316
rect 333112 282276 333118 282288
rect 516134 282276 516140 282288
rect 516192 282276 516198 282328
rect 93946 282208 93952 282260
rect 94004 282248 94010 282260
rect 249886 282248 249892 282260
rect 94004 282220 249892 282248
rect 94004 282208 94010 282220
rect 249886 282208 249892 282220
rect 249944 282208 249950 282260
rect 334434 282208 334440 282260
rect 334492 282248 334498 282260
rect 520274 282248 520280 282260
rect 334492 282220 520280 282248
rect 334492 282208 334498 282220
rect 520274 282208 520280 282220
rect 520332 282208 520338 282260
rect 69014 282140 69020 282192
rect 69072 282180 69078 282192
rect 245838 282180 245844 282192
rect 69072 282152 245844 282180
rect 69072 282140 69078 282152
rect 245838 282140 245844 282152
rect 245896 282140 245902 282192
rect 335538 282140 335544 282192
rect 335596 282180 335602 282192
rect 527174 282180 527180 282192
rect 335596 282152 527180 282180
rect 335596 282140 335602 282152
rect 527174 282140 527180 282152
rect 527232 282140 527238 282192
rect 201494 281052 201500 281104
rect 201552 281092 201558 281104
rect 272242 281092 272248 281104
rect 201552 281064 272248 281092
rect 201552 281052 201558 281064
rect 272242 281052 272248 281064
rect 272300 281052 272306 281104
rect 155954 280984 155960 281036
rect 156012 281024 156018 281036
rect 262490 281024 262496 281036
rect 156012 280996 262496 281024
rect 156012 280984 156018 280996
rect 262490 280984 262496 280996
rect 262548 280984 262554 281036
rect 328822 280984 328828 281036
rect 328880 281024 328886 281036
rect 498194 281024 498200 281036
rect 328880 280996 498200 281024
rect 328880 280984 328886 280996
rect 498194 280984 498200 280996
rect 498252 280984 498258 281036
rect 151814 280916 151820 280968
rect 151872 280956 151878 280968
rect 262582 280956 262588 280968
rect 151872 280928 262588 280956
rect 151872 280916 151878 280928
rect 262582 280916 262588 280928
rect 262640 280916 262646 280968
rect 331398 280916 331404 280968
rect 331456 280956 331462 280968
rect 506566 280956 506572 280968
rect 331456 280928 506572 280956
rect 331456 280916 331462 280928
rect 506566 280916 506572 280928
rect 506624 280916 506630 280968
rect 66254 280848 66260 280900
rect 66312 280888 66318 280900
rect 244550 280888 244556 280900
rect 66312 280860 244556 280888
rect 66312 280848 66318 280860
rect 244550 280848 244556 280860
rect 244608 280848 244614 280900
rect 331490 280848 331496 280900
rect 331548 280888 331554 280900
rect 509234 280888 509240 280900
rect 331548 280860 509240 280888
rect 331548 280848 331554 280860
rect 509234 280848 509240 280860
rect 509292 280848 509298 280900
rect 31754 280780 31760 280832
rect 31812 280820 31818 280832
rect 237742 280820 237748 280832
rect 31812 280792 237748 280820
rect 31812 280780 31818 280792
rect 237742 280780 237748 280792
rect 237800 280780 237806 280832
rect 341058 280780 341064 280832
rect 341116 280820 341122 280832
rect 556246 280820 556252 280832
rect 341116 280792 556252 280820
rect 341116 280780 341122 280792
rect 556246 280780 556252 280792
rect 556304 280780 556310 280832
rect 198734 279760 198740 279812
rect 198792 279800 198798 279812
rect 270862 279800 270868 279812
rect 198792 279772 270868 279800
rect 198792 279760 198798 279772
rect 270862 279760 270868 279772
rect 270920 279760 270926 279812
rect 196618 279692 196624 279744
rect 196676 279732 196682 279744
rect 270954 279732 270960 279744
rect 196676 279704 270960 279732
rect 196676 279692 196682 279704
rect 270954 279692 270960 279704
rect 271012 279692 271018 279744
rect 191834 279624 191840 279676
rect 191892 279664 191898 279676
rect 269482 279664 269488 279676
rect 191892 279636 269488 279664
rect 191892 279624 191898 279636
rect 269482 279624 269488 279636
rect 269540 279624 269546 279676
rect 325970 279624 325976 279676
rect 326028 279664 326034 279676
rect 484394 279664 484400 279676
rect 326028 279636 484400 279664
rect 326028 279624 326034 279636
rect 484394 279624 484400 279636
rect 484452 279624 484458 279676
rect 149054 279556 149060 279608
rect 149112 279596 149118 279608
rect 261294 279596 261300 279608
rect 149112 279568 261300 279596
rect 149112 279556 149118 279568
rect 261294 279556 261300 279568
rect 261352 279556 261358 279608
rect 327350 279556 327356 279608
rect 327408 279596 327414 279608
rect 491294 279596 491300 279608
rect 327408 279568 491300 279596
rect 327408 279556 327414 279568
rect 491294 279556 491300 279568
rect 491352 279556 491358 279608
rect 89714 279488 89720 279540
rect 89772 279528 89778 279540
rect 250254 279528 250260 279540
rect 89772 279500 250260 279528
rect 89772 279488 89778 279500
rect 250254 279488 250260 279500
rect 250312 279488 250318 279540
rect 328730 279488 328736 279540
rect 328788 279528 328794 279540
rect 495434 279528 495440 279540
rect 328788 279500 495440 279528
rect 328788 279488 328794 279500
rect 495434 279488 495440 279500
rect 495492 279488 495498 279540
rect 26878 279420 26884 279472
rect 26936 279460 26942 279472
rect 236270 279460 236276 279472
rect 26936 279432 236276 279460
rect 26936 279420 26942 279432
rect 236270 279420 236276 279432
rect 236328 279420 236334 279472
rect 338482 279420 338488 279472
rect 338540 279460 338546 279472
rect 545114 279460 545120 279472
rect 338540 279432 545120 279460
rect 338540 279420 338546 279432
rect 545114 279420 545120 279432
rect 545172 279420 545178 279472
rect 187694 278264 187700 278316
rect 187752 278304 187758 278316
rect 269390 278304 269396 278316
rect 187752 278276 269396 278304
rect 187752 278264 187758 278276
rect 269390 278264 269396 278276
rect 269448 278264 269454 278316
rect 184934 278196 184940 278248
rect 184992 278236 184998 278248
rect 268194 278236 268200 278248
rect 184992 278208 268200 278236
rect 184992 278196 184998 278208
rect 268194 278196 268200 278208
rect 268252 278196 268258 278248
rect 320542 278196 320548 278248
rect 320600 278236 320606 278248
rect 455414 278236 455420 278248
rect 320600 278208 455420 278236
rect 320600 278196 320606 278208
rect 455414 278196 455420 278208
rect 455472 278196 455478 278248
rect 180794 278128 180800 278180
rect 180852 278168 180858 278180
rect 268102 278168 268108 278180
rect 180852 278140 268108 278168
rect 180852 278128 180858 278140
rect 268102 278128 268108 278140
rect 268160 278128 268166 278180
rect 321646 278128 321652 278180
rect 321704 278168 321710 278180
rect 462314 278168 462320 278180
rect 321704 278140 462320 278168
rect 321704 278128 321710 278140
rect 462314 278128 462320 278140
rect 462372 278128 462378 278180
rect 144914 278060 144920 278112
rect 144972 278100 144978 278112
rect 261202 278100 261208 278112
rect 144972 278072 261208 278100
rect 144972 278060 144978 278072
rect 261202 278060 261208 278072
rect 261260 278060 261266 278112
rect 325878 278060 325884 278112
rect 325936 278100 325942 278112
rect 481726 278100 481732 278112
rect 325936 278072 481732 278100
rect 325936 278060 325942 278072
rect 481726 278060 481732 278072
rect 481784 278060 481790 278112
rect 62114 277992 62120 278044
rect 62172 278032 62178 278044
rect 244458 278032 244464 278044
rect 62172 278004 244464 278032
rect 62172 277992 62178 278004
rect 244458 277992 244464 278004
rect 244516 277992 244522 278044
rect 327258 277992 327264 278044
rect 327316 278032 327322 278044
rect 488534 278032 488540 278044
rect 327316 278004 488540 278032
rect 327316 277992 327322 278004
rect 488534 277992 488540 278004
rect 488592 277992 488598 278044
rect 176654 276904 176660 276956
rect 176712 276944 176718 276956
rect 266630 276944 266636 276956
rect 176712 276916 266636 276944
rect 176712 276904 176718 276916
rect 266630 276904 266636 276916
rect 266688 276904 266694 276956
rect 173894 276836 173900 276888
rect 173952 276876 173958 276888
rect 266722 276876 266728 276888
rect 173952 276848 266728 276876
rect 173952 276836 173958 276848
rect 266722 276836 266728 276848
rect 266780 276836 266786 276888
rect 316126 276836 316132 276888
rect 316184 276876 316190 276888
rect 433334 276876 433340 276888
rect 316184 276848 433340 276876
rect 316184 276836 316190 276848
rect 433334 276836 433340 276848
rect 433392 276836 433398 276888
rect 169754 276768 169760 276820
rect 169812 276808 169818 276820
rect 265434 276808 265440 276820
rect 169812 276780 265440 276808
rect 169812 276768 169818 276780
rect 265434 276768 265440 276780
rect 265492 276768 265498 276820
rect 317782 276768 317788 276820
rect 317840 276808 317846 276820
rect 437474 276808 437480 276820
rect 317840 276780 437480 276808
rect 317840 276768 317846 276780
rect 437474 276768 437480 276780
rect 437532 276768 437538 276820
rect 142154 276700 142160 276752
rect 142212 276740 142218 276752
rect 259914 276740 259920 276752
rect 142212 276712 259920 276740
rect 142212 276700 142218 276712
rect 259914 276700 259920 276712
rect 259972 276700 259978 276752
rect 320450 276700 320456 276752
rect 320508 276740 320514 276752
rect 451274 276740 451280 276752
rect 320508 276712 451280 276740
rect 320508 276700 320514 276712
rect 451274 276700 451280 276712
rect 451332 276700 451338 276752
rect 61378 276632 61384 276684
rect 61436 276672 61442 276684
rect 243354 276672 243360 276684
rect 61436 276644 243360 276672
rect 61436 276632 61442 276644
rect 243354 276632 243360 276644
rect 243412 276632 243418 276684
rect 332962 276632 332968 276684
rect 333020 276672 333026 276684
rect 513374 276672 513380 276684
rect 333020 276644 513380 276672
rect 333020 276632 333026 276644
rect 513374 276632 513380 276644
rect 513432 276632 513438 276684
rect 166994 275408 167000 275460
rect 167052 275448 167058 275460
rect 265342 275448 265348 275460
rect 167052 275420 265348 275448
rect 167052 275408 167058 275420
rect 265342 275408 265348 275420
rect 265400 275408 265406 275460
rect 313366 275408 313372 275460
rect 313424 275448 313430 275460
rect 415486 275448 415492 275460
rect 313424 275420 415492 275448
rect 313424 275408 313430 275420
rect 415486 275408 415492 275420
rect 415544 275408 415550 275460
rect 162854 275340 162860 275392
rect 162912 275380 162918 275392
rect 263962 275380 263968 275392
rect 162912 275352 263968 275380
rect 162912 275340 162918 275352
rect 263962 275340 263968 275352
rect 264020 275340 264026 275392
rect 313458 275340 313464 275392
rect 313516 275380 313522 275392
rect 419534 275380 419540 275392
rect 313516 275352 419540 275380
rect 313516 275340 313522 275352
rect 419534 275340 419540 275352
rect 419592 275340 419598 275392
rect 57238 275272 57244 275324
rect 57296 275312 57302 275324
rect 243262 275312 243268 275324
rect 57296 275284 243268 275312
rect 57296 275272 57302 275284
rect 243262 275272 243268 275284
rect 243320 275272 243326 275324
rect 319070 275272 319076 275324
rect 319128 275312 319134 275324
rect 448514 275312 448520 275324
rect 319128 275284 448520 275312
rect 319128 275272 319134 275284
rect 448514 275272 448520 275284
rect 448572 275272 448578 275324
rect 211798 274252 211804 274304
rect 211856 274292 211862 274304
rect 272058 274292 272064 274304
rect 211856 274264 272064 274292
rect 211856 274252 211862 274264
rect 272058 274252 272064 274264
rect 272116 274252 272122 274304
rect 211154 274184 211160 274236
rect 211212 274224 211218 274236
rect 273622 274224 273628 274236
rect 211212 274196 273628 274224
rect 211212 274184 211218 274196
rect 273622 274184 273628 274196
rect 273680 274184 273686 274236
rect 206278 274116 206284 274168
rect 206336 274156 206342 274168
rect 272150 274156 272156 274168
rect 206336 274128 272156 274156
rect 206336 274116 206342 274128
rect 272150 274116 272156 274128
rect 272208 274116 272214 274168
rect 309226 274116 309232 274168
rect 309284 274156 309290 274168
rect 398926 274156 398932 274168
rect 309284 274128 398932 274156
rect 309284 274116 309290 274128
rect 398926 274116 398932 274128
rect 398984 274116 398990 274168
rect 158714 274048 158720 274100
rect 158772 274088 158778 274100
rect 262398 274088 262404 274100
rect 158772 274060 262404 274088
rect 158772 274048 158778 274060
rect 262398 274048 262404 274060
rect 262456 274048 262462 274100
rect 310606 274048 310612 274100
rect 310664 274088 310670 274100
rect 401594 274088 401600 274100
rect 310664 274060 401600 274088
rect 310664 274048 310670 274060
rect 401594 274048 401600 274060
rect 401652 274048 401658 274100
rect 138014 273980 138020 274032
rect 138072 274020 138078 274032
rect 259822 274020 259828 274032
rect 138072 273992 259828 274020
rect 138072 273980 138078 273992
rect 259822 273980 259828 273992
rect 259880 273980 259886 274032
rect 311986 273980 311992 274032
rect 312044 274020 312050 274032
rect 412634 274020 412640 274032
rect 312044 273992 412640 274020
rect 312044 273980 312050 273992
rect 412634 273980 412640 273992
rect 412692 273980 412698 274032
rect 36538 273912 36544 273964
rect 36596 273952 36602 273964
rect 239030 273952 239036 273964
rect 36596 273924 239036 273952
rect 36596 273912 36602 273924
rect 239030 273912 239036 273924
rect 239088 273912 239094 273964
rect 314746 273912 314752 273964
rect 314804 273952 314810 273964
rect 426434 273952 426440 273964
rect 314804 273924 426440 273952
rect 314804 273912 314810 273924
rect 426434 273912 426440 273924
rect 426492 273912 426498 273964
rect 367738 273164 367744 273216
rect 367796 273204 367802 273216
rect 580166 273204 580172 273216
rect 367796 273176 580172 273204
rect 367796 273164 367802 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 201586 272824 201592 272876
rect 201644 272864 201650 272876
rect 270678 272864 270684 272876
rect 201644 272836 270684 272864
rect 201644 272824 201650 272836
rect 270678 272824 270684 272836
rect 270736 272824 270742 272876
rect 197354 272756 197360 272808
rect 197412 272796 197418 272808
rect 270770 272796 270776 272808
rect 197412 272768 270776 272796
rect 197412 272756 197418 272768
rect 270770 272756 270776 272768
rect 270828 272756 270834 272808
rect 193214 272688 193220 272740
rect 193272 272728 193278 272740
rect 269298 272728 269304 272740
rect 193272 272700 269304 272728
rect 193272 272688 193278 272700
rect 269298 272688 269304 272700
rect 269356 272688 269362 272740
rect 154574 272620 154580 272672
rect 154632 272660 154638 272672
rect 262306 272660 262312 272672
rect 154632 272632 262312 272660
rect 154632 272620 154638 272632
rect 262306 272620 262312 272632
rect 262364 272620 262370 272672
rect 307938 272620 307944 272672
rect 307996 272660 308002 272672
rect 387794 272660 387800 272672
rect 307996 272632 387800 272660
rect 307996 272620 308002 272632
rect 387794 272620 387800 272632
rect 387852 272620 387858 272672
rect 131114 272552 131120 272604
rect 131172 272592 131178 272604
rect 258350 272592 258356 272604
rect 131172 272564 258356 272592
rect 131172 272552 131178 272564
rect 258350 272552 258356 272564
rect 258408 272552 258414 272604
rect 307846 272552 307852 272604
rect 307904 272592 307910 272604
rect 390646 272592 390652 272604
rect 307904 272564 390652 272592
rect 307904 272552 307910 272564
rect 390646 272552 390652 272564
rect 390704 272552 390710 272604
rect 30374 272484 30380 272536
rect 30432 272524 30438 272536
rect 237650 272524 237656 272536
rect 30432 272496 237656 272524
rect 30432 272484 30438 272496
rect 237650 272484 237656 272496
rect 237708 272484 237714 272536
rect 309134 272484 309140 272536
rect 309192 272524 309198 272536
rect 394694 272524 394700 272536
rect 309192 272496 394700 272524
rect 309192 272484 309198 272496
rect 394694 272484 394700 272496
rect 394752 272484 394758 272536
rect 188338 271464 188344 271516
rect 188396 271504 188402 271516
rect 268010 271504 268016 271516
rect 188396 271476 268016 271504
rect 188396 271464 188402 271476
rect 268010 271464 268016 271476
rect 268068 271464 268074 271516
rect 183554 271396 183560 271448
rect 183612 271436 183618 271448
rect 267918 271436 267924 271448
rect 183612 271408 267924 271436
rect 183612 271396 183618 271408
rect 267918 271396 267924 271408
rect 267976 271396 267982 271448
rect 179414 271328 179420 271380
rect 179472 271368 179478 271380
rect 266538 271368 266544 271380
rect 179472 271340 266544 271368
rect 179472 271328 179478 271340
rect 266538 271328 266544 271340
rect 266596 271328 266602 271380
rect 305086 271328 305092 271380
rect 305144 271368 305150 271380
rect 376754 271368 376760 271380
rect 305144 271340 376760 271368
rect 305144 271328 305150 271340
rect 376754 271328 376760 271340
rect 376812 271328 376818 271380
rect 143534 271260 143540 271312
rect 143592 271300 143598 271312
rect 259730 271300 259736 271312
rect 143592 271272 259736 271300
rect 143592 271260 143598 271272
rect 259730 271260 259736 271272
rect 259788 271260 259794 271312
rect 306466 271260 306472 271312
rect 306524 271300 306530 271312
rect 380894 271300 380900 271312
rect 306524 271272 380900 271300
rect 306524 271260 306530 271272
rect 380894 271260 380900 271272
rect 380952 271260 380958 271312
rect 85666 271192 85672 271244
rect 85724 271232 85730 271244
rect 248598 271232 248604 271244
rect 85724 271204 248604 271232
rect 85724 271192 85730 271204
rect 248598 271192 248604 271204
rect 248656 271192 248662 271244
rect 306558 271192 306564 271244
rect 306616 271232 306622 271244
rect 383654 271232 383660 271244
rect 306616 271204 383660 271232
rect 306616 271192 306622 271204
rect 383654 271192 383660 271204
rect 383712 271192 383718 271244
rect 27614 271124 27620 271176
rect 27672 271164 27678 271176
rect 237558 271164 237564 271176
rect 27672 271136 237564 271164
rect 27672 271124 27678 271136
rect 237558 271124 237564 271136
rect 237616 271124 237622 271176
rect 318978 271124 318984 271176
rect 319036 271164 319042 271176
rect 444374 271164 444380 271176
rect 319036 271136 444380 271164
rect 319036 271124 319042 271136
rect 444374 271124 444380 271136
rect 444432 271124 444438 271176
rect 178770 270104 178776 270156
rect 178828 270144 178834 270156
rect 266446 270144 266452 270156
rect 178828 270116 266452 270144
rect 178828 270104 178834 270116
rect 266446 270104 266452 270116
rect 266504 270104 266510 270156
rect 172514 270036 172520 270088
rect 172572 270076 172578 270088
rect 265250 270076 265256 270088
rect 172572 270048 265256 270076
rect 172572 270036 172578 270048
rect 265250 270036 265256 270048
rect 265308 270036 265314 270088
rect 168374 269968 168380 270020
rect 168432 270008 168438 270020
rect 265158 270008 265164 270020
rect 168432 269980 265164 270008
rect 168432 269968 168438 269980
rect 265158 269968 265164 269980
rect 265216 269968 265222 270020
rect 304994 269968 305000 270020
rect 305052 270008 305058 270020
rect 374086 270008 374092 270020
rect 305052 269980 374092 270008
rect 305052 269968 305058 269980
rect 374086 269968 374092 269980
rect 374144 269968 374150 270020
rect 140774 269900 140780 269952
rect 140832 269940 140838 269952
rect 259638 269940 259644 269952
rect 140832 269912 259644 269940
rect 140832 269900 140838 269912
rect 259638 269900 259644 269912
rect 259696 269900 259702 269952
rect 320358 269900 320364 269952
rect 320416 269940 320422 269952
rect 449894 269940 449900 269952
rect 320416 269912 449900 269940
rect 320416 269900 320422 269912
rect 449894 269900 449900 269912
rect 449952 269900 449958 269952
rect 82814 269832 82820 269884
rect 82872 269872 82878 269884
rect 248506 269872 248512 269884
rect 82872 269844 248512 269872
rect 82872 269832 82878 269844
rect 248506 269832 248512 269844
rect 248564 269832 248570 269884
rect 342346 269832 342352 269884
rect 342404 269872 342410 269884
rect 520918 269872 520924 269884
rect 342404 269844 520924 269872
rect 342404 269832 342410 269844
rect 520918 269832 520924 269844
rect 520976 269832 520982 269884
rect 13814 269764 13820 269816
rect 13872 269804 13878 269816
rect 235074 269804 235080 269816
rect 13872 269776 235080 269804
rect 13872 269764 13878 269776
rect 235074 269764 235080 269776
rect 235132 269764 235138 269816
rect 343818 269764 343824 269816
rect 343876 269804 343882 269816
rect 525058 269804 525064 269816
rect 343876 269776 525064 269804
rect 343876 269764 343882 269776
rect 525058 269764 525064 269776
rect 525116 269764 525122 269816
rect 165614 268608 165620 268660
rect 165672 268648 165678 268660
rect 263778 268648 263784 268660
rect 165672 268620 263784 268648
rect 165672 268608 165678 268620
rect 263778 268608 263784 268620
rect 263836 268608 263842 268660
rect 303706 268608 303712 268660
rect 303764 268648 303770 268660
rect 365714 268648 365720 268660
rect 303764 268620 365720 268648
rect 303764 268608 303770 268620
rect 365714 268608 365720 268620
rect 365772 268608 365778 268660
rect 161474 268540 161480 268592
rect 161532 268580 161538 268592
rect 263870 268580 263876 268592
rect 161532 268552 263876 268580
rect 161532 268540 161538 268552
rect 263870 268540 263876 268552
rect 263928 268540 263934 268592
rect 339494 268540 339500 268592
rect 339552 268580 339558 268592
rect 508498 268580 508504 268592
rect 339552 268552 508504 268580
rect 339552 268540 339558 268552
rect 508498 268540 508504 268552
rect 508556 268540 508562 268592
rect 157334 268472 157340 268524
rect 157392 268512 157398 268524
rect 262674 268512 262680 268524
rect 157392 268484 262680 268512
rect 157392 268472 157398 268484
rect 262674 268472 262680 268484
rect 262732 268472 262738 268524
rect 339586 268472 339592 268524
rect 339644 268512 339650 268524
rect 516778 268512 516784 268524
rect 339644 268484 516784 268512
rect 339644 268472 339650 268484
rect 516778 268472 516784 268484
rect 516836 268472 516842 268524
rect 136634 268404 136640 268456
rect 136692 268444 136698 268456
rect 258258 268444 258264 268456
rect 136692 268416 258264 268444
rect 136692 268404 136698 268416
rect 258258 268404 258264 268416
rect 258316 268404 258322 268456
rect 332870 268404 332876 268456
rect 332928 268444 332934 268456
rect 514846 268444 514852 268456
rect 332928 268416 514852 268444
rect 332928 268404 332934 268416
rect 514846 268404 514852 268416
rect 514904 268404 514910 268456
rect 52546 268336 52552 268388
rect 52604 268376 52610 268388
rect 241790 268376 241796 268388
rect 52604 268348 241796 268376
rect 52604 268336 52610 268348
rect 241790 268336 241796 268348
rect 241848 268336 241854 268388
rect 338390 268336 338396 268388
rect 338448 268376 338454 268388
rect 547966 268376 547972 268388
rect 338448 268348 547972 268376
rect 338448 268336 338454 268348
rect 547966 268336 547972 268348
rect 548024 268336 548030 268388
rect 3234 267656 3240 267708
rect 3292 267696 3298 267708
rect 228358 267696 228364 267708
rect 3292 267668 228364 267696
rect 3292 267656 3298 267668
rect 228358 267656 228364 267668
rect 228416 267656 228422 267708
rect 153194 267180 153200 267232
rect 153252 267220 153258 267232
rect 260098 267220 260104 267232
rect 153252 267192 260104 267220
rect 153252 267180 153258 267192
rect 260098 267180 260104 267192
rect 260156 267180 260162 267232
rect 335446 267180 335452 267232
rect 335504 267220 335510 267232
rect 496078 267220 496084 267232
rect 335504 267192 496084 267220
rect 335504 267180 335510 267192
rect 496078 267180 496084 267192
rect 496136 267180 496142 267232
rect 150434 267112 150440 267164
rect 150492 267152 150498 267164
rect 261110 267152 261116 267164
rect 150492 267124 261116 267152
rect 150492 267112 150498 267124
rect 261110 267112 261116 267124
rect 261168 267112 261174 267164
rect 336918 267112 336924 267164
rect 336976 267152 336982 267164
rect 502978 267152 502984 267164
rect 336976 267124 502984 267152
rect 336976 267112 336982 267124
rect 502978 267112 502984 267124
rect 503036 267112 503042 267164
rect 64874 267044 64880 267096
rect 64932 267084 64938 267096
rect 244366 267084 244372 267096
rect 64932 267056 244372 267084
rect 64932 267044 64938 267056
rect 244366 267044 244372 267056
rect 244424 267044 244430 267096
rect 334342 267044 334348 267096
rect 334400 267084 334406 267096
rect 523126 267084 523132 267096
rect 334400 267056 523132 267084
rect 334400 267044 334406 267056
rect 523126 267044 523132 267056
rect 523184 267044 523190 267096
rect 22094 266976 22100 267028
rect 22152 267016 22158 267028
rect 236178 267016 236184 267028
rect 22152 266988 236184 267016
rect 22152 266976 22158 266988
rect 236178 266976 236184 266988
rect 236236 266976 236242 267028
rect 337010 266976 337016 267028
rect 337068 267016 337074 267028
rect 539686 267016 539692 267028
rect 337068 266988 539692 267016
rect 337068 266976 337074 266988
rect 539686 266976 539692 266988
rect 539744 266976 539750 267028
rect 209774 265820 209780 265872
rect 209832 265860 209838 265872
rect 273438 265860 273444 265872
rect 209832 265832 273444 265860
rect 209832 265820 209838 265832
rect 273438 265820 273444 265832
rect 273496 265820 273502 265872
rect 311894 265820 311900 265872
rect 311952 265860 311958 265872
rect 408494 265860 408500 265872
rect 311952 265832 408500 265860
rect 311952 265820 311958 265832
rect 408494 265820 408500 265832
rect 408552 265820 408558 265872
rect 146294 265752 146300 265804
rect 146352 265792 146358 265804
rect 261018 265792 261024 265804
rect 146352 265764 261024 265792
rect 146352 265752 146358 265764
rect 261018 265752 261024 265764
rect 261076 265752 261082 265804
rect 332778 265752 332784 265804
rect 332836 265792 332842 265804
rect 440878 265792 440884 265804
rect 332836 265764 440884 265792
rect 332836 265752 332842 265764
rect 440878 265752 440884 265764
rect 440936 265752 440942 265804
rect 133874 265684 133880 265736
rect 133932 265724 133938 265736
rect 258166 265724 258172 265736
rect 133932 265696 258172 265724
rect 133932 265684 133938 265696
rect 258166 265684 258172 265696
rect 258224 265684 258230 265736
rect 334250 265684 334256 265736
rect 334308 265724 334314 265736
rect 446398 265724 446404 265736
rect 334308 265696 446404 265724
rect 334308 265684 334314 265696
rect 446398 265684 446404 265696
rect 446456 265684 446462 265736
rect 48314 265616 48320 265668
rect 48372 265656 48378 265668
rect 241698 265656 241704 265668
rect 48372 265628 241704 265656
rect 48372 265616 48378 265628
rect 241698 265616 241704 265628
rect 241756 265616 241762 265668
rect 334158 265616 334164 265668
rect 334216 265656 334222 265668
rect 525794 265656 525800 265668
rect 334216 265628 525800 265656
rect 334216 265616 334222 265628
rect 525794 265616 525800 265628
rect 525852 265616 525858 265668
rect 207014 264528 207020 264580
rect 207072 264568 207078 264580
rect 271966 264568 271972 264580
rect 207072 264540 271972 264568
rect 207072 264528 207078 264540
rect 271966 264528 271972 264540
rect 272024 264528 272030 264580
rect 195974 264460 195980 264512
rect 196032 264500 196038 264512
rect 270586 264500 270592 264512
rect 196032 264472 270592 264500
rect 196032 264460 196038 264472
rect 270586 264460 270592 264472
rect 270644 264460 270650 264512
rect 193306 264392 193312 264444
rect 193364 264432 193370 264444
rect 269206 264432 269212 264444
rect 193364 264404 269212 264432
rect 193364 264392 193370 264404
rect 269206 264392 269212 264404
rect 269264 264392 269270 264444
rect 332686 264392 332692 264444
rect 332744 264432 332750 264444
rect 432598 264432 432604 264444
rect 332744 264404 432604 264432
rect 332744 264392 332750 264404
rect 432598 264392 432604 264404
rect 432656 264392 432662 264444
rect 143626 264324 143632 264376
rect 143684 264364 143690 264376
rect 259546 264364 259552 264376
rect 143684 264336 259552 264364
rect 143684 264324 143690 264336
rect 259546 264324 259552 264336
rect 259604 264324 259610 264376
rect 317690 264324 317696 264376
rect 317748 264364 317754 264376
rect 440234 264364 440240 264376
rect 317748 264336 440240 264364
rect 317748 264324 317754 264336
rect 440234 264324 440240 264336
rect 440292 264324 440298 264376
rect 126974 264256 126980 264308
rect 127032 264296 127038 264308
rect 257062 264296 257068 264308
rect 127032 264268 257068 264296
rect 127032 264256 127038 264268
rect 257062 264256 257068 264268
rect 257120 264256 257126 264308
rect 331214 264256 331220 264308
rect 331272 264296 331278 264308
rect 507854 264296 507860 264308
rect 331272 264268 507860 264296
rect 331272 264256 331278 264268
rect 507854 264256 507860 264268
rect 507912 264256 507918 264308
rect 44174 264188 44180 264240
rect 44232 264228 44238 264240
rect 240410 264228 240416 264240
rect 44232 264200 240416 264228
rect 44232 264188 44238 264200
rect 240410 264188 240416 264200
rect 240468 264188 240474 264240
rect 331306 264188 331312 264240
rect 331364 264228 331370 264240
rect 511994 264228 512000 264240
rect 331364 264200 512000 264228
rect 331364 264188 331370 264200
rect 511994 264188 512000 264200
rect 512052 264188 512058 264240
rect 175274 263100 175280 263152
rect 175332 263140 175338 263152
rect 253290 263140 253296 263152
rect 175332 263112 253296 263140
rect 175332 263100 175338 263112
rect 253290 263100 253296 263112
rect 253348 263100 253354 263152
rect 185026 263032 185032 263084
rect 185084 263072 185090 263084
rect 267734 263072 267740 263084
rect 185084 263044 267740 263072
rect 185084 263032 185090 263044
rect 267734 263032 267740 263044
rect 267792 263032 267798 263084
rect 330018 263032 330024 263084
rect 330076 263072 330082 263084
rect 417418 263072 417424 263084
rect 330076 263044 417424 263072
rect 330076 263032 330082 263044
rect 417418 263032 417424 263044
rect 417476 263032 417482 263084
rect 182174 262964 182180 263016
rect 182232 263004 182238 263016
rect 267826 263004 267832 263016
rect 182232 262976 267832 263004
rect 182232 262964 182238 262976
rect 267826 262964 267832 262976
rect 267884 262964 267890 263016
rect 316034 262964 316040 263016
rect 316092 263004 316098 263016
rect 432046 263004 432052 263016
rect 316092 262976 432052 263004
rect 316092 262964 316098 262976
rect 432046 262964 432052 262976
rect 432104 262964 432110 263016
rect 139394 262896 139400 262948
rect 139452 262936 139458 262948
rect 259454 262936 259460 262948
rect 139452 262908 259460 262936
rect 139452 262896 139458 262908
rect 259454 262896 259460 262908
rect 259512 262896 259518 262948
rect 328638 262896 328644 262948
rect 328696 262936 328702 262948
rect 498286 262936 498292 262948
rect 328696 262908 498292 262936
rect 328696 262896 328702 262908
rect 498286 262896 498292 262908
rect 498344 262896 498350 262948
rect 40034 262828 40040 262880
rect 40092 262868 40098 262880
rect 240318 262868 240324 262880
rect 40092 262840 240324 262868
rect 40092 262828 40098 262840
rect 240318 262828 240324 262840
rect 240376 262828 240382 262880
rect 343726 262828 343732 262880
rect 343784 262868 343790 262880
rect 575474 262868 575480 262880
rect 343784 262840 575480 262868
rect 343784 262828 343790 262840
rect 575474 262828 575480 262840
rect 575532 262828 575538 262880
rect 207658 261808 207664 261860
rect 207716 261848 207722 261860
rect 266814 261848 266820 261860
rect 207716 261820 266820 261848
rect 207716 261808 207722 261820
rect 266814 261808 266820 261820
rect 266872 261808 266878 261860
rect 171134 261740 171140 261792
rect 171192 261780 171198 261792
rect 264974 261780 264980 261792
rect 171192 261752 264980 261780
rect 171192 261740 171198 261752
rect 264974 261740 264980 261752
rect 265032 261740 265038 261792
rect 168466 261672 168472 261724
rect 168524 261712 168530 261724
rect 265066 261712 265072 261724
rect 168524 261684 265072 261712
rect 168524 261672 168530 261684
rect 265066 261672 265072 261684
rect 265124 261672 265130 261724
rect 327074 261672 327080 261724
rect 327132 261712 327138 261724
rect 487154 261712 487160 261724
rect 327132 261684 487160 261712
rect 327132 261672 327138 261684
rect 487154 261672 487160 261684
rect 487212 261672 487218 261724
rect 164234 261604 164240 261656
rect 164292 261644 164298 261656
rect 263686 261644 263692 261656
rect 164292 261616 263692 261644
rect 164292 261604 164298 261616
rect 263686 261604 263692 261616
rect 263744 261604 263750 261656
rect 327166 261604 327172 261656
rect 327224 261644 327230 261656
rect 490006 261644 490012 261656
rect 327224 261616 490012 261644
rect 327224 261604 327230 261616
rect 490006 261604 490012 261616
rect 490064 261604 490070 261656
rect 128354 261536 128360 261588
rect 128412 261576 128418 261588
rect 256970 261576 256976 261588
rect 128412 261548 256976 261576
rect 128412 261536 128418 261548
rect 256970 261536 256976 261548
rect 257028 261536 257034 261588
rect 328546 261536 328552 261588
rect 328604 261576 328610 261588
rect 494054 261576 494060 261588
rect 328604 261548 494060 261576
rect 328604 261536 328610 261548
rect 494054 261536 494060 261548
rect 494112 261536 494118 261588
rect 35250 261468 35256 261520
rect 35308 261508 35314 261520
rect 238938 261508 238944 261520
rect 35308 261480 238944 261508
rect 35308 261468 35314 261480
rect 238938 261468 238944 261480
rect 238996 261468 239002 261520
rect 338298 261468 338304 261520
rect 338356 261508 338362 261520
rect 543734 261508 543740 261520
rect 338356 261480 543740 261508
rect 338356 261468 338362 261480
rect 543734 261468 543740 261480
rect 543792 261468 543798 261520
rect 160186 260312 160192 260364
rect 160244 260352 160250 260364
rect 263594 260352 263600 260364
rect 160244 260324 263600 260352
rect 160244 260312 160250 260324
rect 263594 260312 263600 260324
rect 263652 260312 263658 260364
rect 125594 260244 125600 260296
rect 125652 260284 125658 260296
rect 256878 260284 256884 260296
rect 125652 260256 256884 260284
rect 125652 260244 125658 260256
rect 256878 260244 256884 260256
rect 256936 260244 256942 260296
rect 60734 260176 60740 260228
rect 60792 260216 60798 260228
rect 244734 260216 244740 260228
rect 60792 260188 244740 260216
rect 60792 260176 60798 260188
rect 244734 260176 244740 260188
rect 244792 260176 244798 260228
rect 325786 260176 325792 260228
rect 325844 260216 325850 260228
rect 483014 260216 483020 260228
rect 325844 260188 483020 260216
rect 325844 260176 325850 260188
rect 483014 260176 483020 260188
rect 483072 260176 483078 260228
rect 8294 260108 8300 260160
rect 8352 260148 8358 260160
rect 233510 260148 233516 260160
rect 8352 260120 233516 260148
rect 8352 260108 8358 260120
rect 233510 260108 233516 260120
rect 233568 260108 233574 260160
rect 335354 260108 335360 260160
rect 335412 260148 335418 260160
rect 529934 260148 529940 260160
rect 335412 260120 529940 260148
rect 335412 260108 335418 260120
rect 529934 260108 529940 260120
rect 529992 260108 529998 260160
rect 51074 258884 51080 258936
rect 51132 258924 51138 258936
rect 241606 258924 241612 258936
rect 51132 258896 241612 258924
rect 51132 258884 51138 258896
rect 241606 258884 241612 258896
rect 241664 258884 241670 258936
rect 35894 258816 35900 258868
rect 35952 258856 35958 258868
rect 238846 258856 238852 258868
rect 35952 258828 238852 258856
rect 35952 258816 35958 258828
rect 238846 258816 238852 258828
rect 238904 258816 238910 258868
rect 3694 258748 3700 258800
rect 3752 258788 3758 258800
rect 231118 258788 231124 258800
rect 3752 258760 231124 258788
rect 3752 258748 3758 258760
rect 231118 258748 231124 258760
rect 231176 258748 231182 258800
rect 4798 258680 4804 258732
rect 4856 258720 4862 258732
rect 231854 258720 231860 258732
rect 4856 258692 231860 258720
rect 4856 258680 4862 258692
rect 231854 258680 231860 258692
rect 231912 258680 231918 258732
rect 217134 257320 217140 257372
rect 217192 257360 217198 257372
rect 345474 257360 345480 257372
rect 217192 257332 345480 257360
rect 217192 257320 217198 257332
rect 345474 257320 345480 257332
rect 345532 257320 345538 257372
rect 321554 256164 321560 256216
rect 321612 256204 321618 256216
rect 460934 256204 460940 256216
rect 321612 256176 460940 256204
rect 321612 256164 321618 256176
rect 460934 256164 460940 256176
rect 460992 256164 460998 256216
rect 24854 256096 24860 256148
rect 24912 256136 24918 256148
rect 236086 256136 236092 256148
rect 24912 256108 236092 256136
rect 24912 256096 24918 256108
rect 236086 256096 236092 256108
rect 236144 256096 236150 256148
rect 323210 256096 323216 256148
rect 323268 256136 323274 256148
rect 465074 256136 465080 256148
rect 323268 256108 465080 256136
rect 323268 256096 323274 256108
rect 465074 256096 465080 256108
rect 465132 256096 465138 256148
rect 17218 256028 17224 256080
rect 17276 256068 17282 256080
rect 234982 256068 234988 256080
rect 17276 256040 234988 256068
rect 17276 256028 17282 256040
rect 234982 256028 234988 256040
rect 235040 256028 235046 256080
rect 324406 256028 324412 256080
rect 324464 256068 324470 256080
rect 474734 256068 474740 256080
rect 324464 256040 474740 256068
rect 324464 256028 324470 256040
rect 474734 256028 474740 256040
rect 474792 256028 474798 256080
rect 7558 255960 7564 256012
rect 7616 256000 7622 256012
rect 233418 256000 233424 256012
rect 7616 255972 233424 256000
rect 7616 255960 7622 255972
rect 233418 255960 233424 255972
rect 233476 255960 233482 256012
rect 325694 255960 325700 256012
rect 325752 256000 325758 256012
rect 478874 256000 478880 256012
rect 325752 255972 478880 256000
rect 325752 255960 325758 255972
rect 478874 255960 478880 255972
rect 478932 255960 478938 256012
rect 116578 254804 116584 254856
rect 116636 254844 116642 254856
rect 240594 254844 240600 254856
rect 116636 254816 240600 254844
rect 116636 254804 116642 254816
rect 240594 254804 240600 254816
rect 240652 254804 240658 254856
rect 79318 254736 79324 254788
rect 79376 254776 79382 254788
rect 243078 254776 243084 254788
rect 79376 254748 243084 254776
rect 79376 254736 79382 254748
rect 243078 254736 243084 254748
rect 243136 254736 243142 254788
rect 302418 254736 302424 254788
rect 302476 254776 302482 254788
rect 361574 254776 361580 254788
rect 302476 254748 361580 254776
rect 302476 254736 302482 254748
rect 361574 254736 361580 254748
rect 361632 254736 361638 254788
rect 56594 254668 56600 254720
rect 56652 254708 56658 254720
rect 243170 254708 243176 254720
rect 56652 254680 243176 254708
rect 56652 254668 56658 254680
rect 243170 254668 243176 254680
rect 243228 254668 243234 254720
rect 313274 254668 313280 254720
rect 313332 254708 313338 254720
rect 385678 254708 385684 254720
rect 313332 254680 385684 254708
rect 313332 254668 313338 254680
rect 385678 254668 385684 254680
rect 385736 254668 385742 254720
rect 44266 254600 44272 254652
rect 44324 254640 44330 254652
rect 240226 254640 240232 254652
rect 44324 254612 240232 254640
rect 44324 254600 44330 254612
rect 240226 254600 240232 254612
rect 240284 254600 240290 254652
rect 318886 254600 318892 254652
rect 318944 254640 318950 254652
rect 442994 254640 443000 254652
rect 318944 254612 443000 254640
rect 318944 254600 318950 254612
rect 442994 254600 443000 254612
rect 443052 254600 443058 254652
rect 39298 254532 39304 254584
rect 39356 254572 39362 254584
rect 239214 254572 239220 254584
rect 39356 254544 239220 254572
rect 39356 254532 39362 254544
rect 239214 254532 239220 254544
rect 239272 254532 239278 254584
rect 345382 254532 345388 254584
rect 345440 254572 345446 254584
rect 578234 254572 578240 254584
rect 345440 254544 578240 254572
rect 345440 254532 345446 254544
rect 578234 254532 578240 254544
rect 578292 254532 578298 254584
rect 2774 254328 2780 254380
rect 2832 254368 2838 254380
rect 4890 254368 4896 254380
rect 2832 254340 4896 254368
rect 2832 254328 2838 254340
rect 4890 254328 4896 254340
rect 4948 254328 4954 254380
rect 301222 253512 301228 253564
rect 301280 253552 301286 253564
rect 361666 253552 361672 253564
rect 301280 253524 361672 253552
rect 301280 253512 301286 253524
rect 361666 253512 361672 253524
rect 361724 253512 361730 253564
rect 84194 253444 84200 253496
rect 84252 253484 84258 253496
rect 248414 253484 248420 253496
rect 84252 253456 248420 253484
rect 84252 253444 84258 253456
rect 248414 253444 248420 253456
rect 248472 253444 248478 253496
rect 301314 253444 301320 253496
rect 301372 253484 301378 253496
rect 365806 253484 365812 253496
rect 301372 253456 365812 253484
rect 301372 253444 301378 253456
rect 365806 253444 365812 253456
rect 365864 253444 365870 253496
rect 80054 253376 80060 253428
rect 80112 253416 80118 253428
rect 247218 253416 247224 253428
rect 80112 253388 247224 253416
rect 80112 253376 80118 253388
rect 247218 253376 247224 253388
rect 247276 253376 247282 253428
rect 332594 253376 332600 253428
rect 332652 253416 332658 253428
rect 517514 253416 517520 253428
rect 332652 253388 517520 253416
rect 332652 253376 332658 253388
rect 517514 253376 517520 253388
rect 517572 253376 517578 253428
rect 17954 253308 17960 253360
rect 18012 253348 18018 253360
rect 234798 253348 234804 253360
rect 18012 253320 234804 253348
rect 18012 253308 18018 253320
rect 234798 253308 234804 253320
rect 234856 253308 234862 253360
rect 334066 253308 334072 253360
rect 334124 253348 334130 253360
rect 521654 253348 521660 253360
rect 334124 253320 521660 253348
rect 334124 253308 334130 253320
rect 521654 253308 521660 253320
rect 521712 253308 521718 253360
rect 12434 253240 12440 253292
rect 12492 253280 12498 253292
rect 234890 253280 234896 253292
rect 12492 253252 234896 253280
rect 12492 253240 12498 253252
rect 234890 253240 234896 253252
rect 234948 253240 234954 253292
rect 333974 253240 333980 253292
rect 334032 253280 334038 253292
rect 524414 253280 524420 253292
rect 334032 253252 524420 253280
rect 334032 253240 334038 253252
rect 524414 253240 524420 253252
rect 524472 253240 524478 253292
rect 9674 253172 9680 253224
rect 9732 253212 9738 253224
rect 233326 253212 233332 253224
rect 9732 253184 233332 253212
rect 9732 253172 9738 253184
rect 233326 253172 233332 253184
rect 233384 253172 233390 253224
rect 343634 253172 343640 253224
rect 343692 253212 343698 253224
rect 571334 253212 571340 253224
rect 343692 253184 571340 253212
rect 343692 253172 343698 253184
rect 571334 253172 571340 253184
rect 571392 253172 571398 253224
rect 121454 252084 121460 252136
rect 121512 252124 121518 252136
rect 255406 252124 255412 252136
rect 121512 252096 255412 252124
rect 121512 252084 121518 252096
rect 255406 252084 255412 252096
rect 255464 252084 255470 252136
rect 118786 252016 118792 252068
rect 118844 252056 118850 252068
rect 255774 252056 255780 252068
rect 118844 252028 255780 252056
rect 118844 252016 118850 252028
rect 255774 252016 255780 252028
rect 255832 252016 255838 252068
rect 318794 252016 318800 252068
rect 318852 252056 318858 252068
rect 448606 252056 448612 252068
rect 318852 252028 448612 252056
rect 318852 252016 318858 252028
rect 448606 252016 448612 252028
rect 448664 252016 448670 252068
rect 31018 251948 31024 252000
rect 31076 251988 31082 252000
rect 237466 251988 237472 252000
rect 31076 251960 237472 251988
rect 31076 251948 31082 251960
rect 237466 251948 237472 251960
rect 237524 251948 237530 252000
rect 320266 251948 320272 252000
rect 320324 251988 320330 252000
rect 452654 251988 452660 252000
rect 320324 251960 452660 251988
rect 320324 251948 320330 251960
rect 452654 251948 452660 251960
rect 452712 251948 452718 252000
rect 26234 251880 26240 251932
rect 26292 251920 26298 251932
rect 237834 251920 237840 251932
rect 26292 251892 237840 251920
rect 26292 251880 26298 251892
rect 237834 251880 237840 251892
rect 237892 251880 237898 251932
rect 320174 251880 320180 251932
rect 320232 251920 320238 251932
rect 456886 251920 456892 251932
rect 320232 251892 456892 251920
rect 320232 251880 320238 251892
rect 456886 251880 456892 251892
rect 456944 251880 456950 251932
rect 20714 251812 20720 251864
rect 20772 251852 20778 251864
rect 236362 251852 236368 251864
rect 20772 251824 236368 251852
rect 20772 251812 20778 251824
rect 236362 251812 236368 251824
rect 236420 251812 236426 251864
rect 323026 251812 323032 251864
rect 323084 251852 323090 251864
rect 466454 251852 466460 251864
rect 323084 251824 466460 251852
rect 323084 251812 323090 251824
rect 466454 251812 466460 251824
rect 466512 251812 466518 251864
rect 299750 251132 299756 251184
rect 299808 251172 299814 251184
rect 364702 251172 364708 251184
rect 299808 251144 364708 251172
rect 299808 251132 299814 251144
rect 364702 251132 364708 251144
rect 364760 251132 364766 251184
rect 299934 251064 299940 251116
rect 299992 251104 299998 251116
rect 366174 251104 366180 251116
rect 299992 251076 366180 251104
rect 299992 251064 299998 251076
rect 366174 251064 366180 251076
rect 366232 251064 366238 251116
rect 292942 250996 292948 251048
rect 293000 251036 293006 251048
rect 360194 251036 360200 251048
rect 293000 251008 360200 251036
rect 293000 250996 293006 251008
rect 360194 250996 360200 251008
rect 360252 250996 360258 251048
rect 298278 250928 298284 250980
rect 298336 250968 298342 250980
rect 365898 250968 365904 250980
rect 298336 250940 365904 250968
rect 298336 250928 298342 250940
rect 365898 250928 365904 250940
rect 365956 250928 365962 250980
rect 298370 250860 298376 250912
rect 298428 250900 298434 250912
rect 366082 250900 366088 250912
rect 298428 250872 366088 250900
rect 298428 250860 298434 250872
rect 366082 250860 366088 250872
rect 366140 250860 366146 250912
rect 297174 250792 297180 250844
rect 297232 250832 297238 250844
rect 366266 250832 366272 250844
rect 297232 250804 366272 250832
rect 297232 250792 297238 250804
rect 366266 250792 366272 250804
rect 366324 250792 366330 250844
rect 174538 250724 174544 250776
rect 174596 250764 174602 250776
rect 251634 250764 251640 250776
rect 174596 250736 251640 250764
rect 174596 250724 174602 250736
rect 251634 250724 251640 250736
rect 251692 250724 251698 250776
rect 294138 250724 294144 250776
rect 294196 250764 294202 250776
rect 363506 250764 363512 250776
rect 294196 250736 363512 250764
rect 294196 250724 294202 250736
rect 363506 250724 363512 250736
rect 363564 250724 363570 250776
rect 78674 250656 78680 250708
rect 78732 250696 78738 250708
rect 247126 250696 247132 250708
rect 78732 250668 247132 250696
rect 78732 250656 78738 250668
rect 247126 250656 247132 250668
rect 247184 250656 247190 250708
rect 294046 250656 294052 250708
rect 294104 250696 294110 250708
rect 365990 250696 365996 250708
rect 294104 250668 365996 250696
rect 294104 250656 294110 250668
rect 365990 250656 365996 250668
rect 366048 250656 366054 250708
rect 75914 250588 75920 250640
rect 75972 250628 75978 250640
rect 247034 250628 247040 250640
rect 75972 250600 247040 250628
rect 75972 250588 75978 250600
rect 247034 250588 247040 250600
rect 247092 250588 247098 250640
rect 291562 250588 291568 250640
rect 291620 250628 291626 250640
rect 368474 250628 368480 250640
rect 291620 250600 368480 250628
rect 291620 250588 291626 250600
rect 368474 250588 368480 250600
rect 368532 250588 368538 250640
rect 71774 250520 71780 250572
rect 71832 250560 71838 250572
rect 245746 250560 245752 250572
rect 71832 250532 245752 250560
rect 71832 250520 71838 250532
rect 245746 250520 245752 250532
rect 245804 250520 245810 250572
rect 306374 250520 306380 250572
rect 306432 250560 306438 250572
rect 385034 250560 385040 250572
rect 306432 250532 385040 250560
rect 306432 250520 306438 250532
rect 385034 250520 385040 250532
rect 385092 250520 385098 250572
rect 16574 250452 16580 250504
rect 16632 250492 16638 250504
rect 234706 250492 234712 250504
rect 16632 250464 234712 250492
rect 16632 250452 16638 250464
rect 234706 250452 234712 250464
rect 234764 250452 234770 250504
rect 307754 250452 307760 250504
rect 307812 250492 307818 250504
rect 389174 250492 389180 250504
rect 307812 250464 389180 250492
rect 307812 250452 307818 250464
rect 389174 250452 389180 250464
rect 389232 250452 389238 250504
rect 299842 250384 299848 250436
rect 299900 250424 299906 250436
rect 362954 250424 362960 250436
rect 299900 250396 362960 250424
rect 299900 250384 299906 250396
rect 362954 250384 362960 250396
rect 363012 250384 363018 250436
rect 295794 250316 295800 250368
rect 295852 250356 295858 250368
rect 358814 250356 358820 250368
rect 295852 250328 358820 250356
rect 295852 250316 295858 250328
rect 358814 250316 358820 250328
rect 358872 250316 358878 250368
rect 295702 250248 295708 250300
rect 295760 250288 295766 250300
rect 357434 250288 357440 250300
rect 295760 250260 357440 250288
rect 295760 250248 295766 250260
rect 357434 250248 357440 250260
rect 357492 250248 357498 250300
rect 209866 249228 209872 249280
rect 209924 249268 209930 249280
rect 273254 249268 273260 249280
rect 209924 249240 273260 249268
rect 209924 249228 209930 249240
rect 273254 249228 273260 249240
rect 273312 249228 273318 249280
rect 317506 249228 317512 249280
rect 317564 249268 317570 249280
rect 436094 249268 436100 249280
rect 317564 249240 436100 249268
rect 317564 249228 317570 249240
rect 436094 249228 436100 249240
rect 436152 249228 436158 249280
rect 205634 249160 205640 249212
rect 205692 249200 205698 249212
rect 272334 249200 272340 249212
rect 205692 249172 272340 249200
rect 205692 249160 205698 249172
rect 272334 249160 272340 249172
rect 272392 249160 272398 249212
rect 338114 249160 338120 249212
rect 338172 249200 338178 249212
rect 534718 249200 534724 249212
rect 338172 249172 534724 249200
rect 338172 249160 338178 249172
rect 534718 249160 534724 249172
rect 534776 249160 534782 249212
rect 135254 249092 135260 249144
rect 135312 249132 135318 249144
rect 258442 249132 258448 249144
rect 135312 249104 258448 249132
rect 135312 249092 135318 249104
rect 258442 249092 258448 249104
rect 258500 249092 258506 249144
rect 336826 249092 336832 249144
rect 336884 249132 336890 249144
rect 534074 249132 534080 249144
rect 336884 249104 534080 249132
rect 336884 249092 336890 249104
rect 534074 249092 534080 249104
rect 534132 249092 534138 249144
rect 13078 249024 13084 249076
rect 13136 249064 13142 249076
rect 234614 249064 234620 249076
rect 13136 249036 234620 249064
rect 13136 249024 13142 249036
rect 234614 249024 234620 249036
rect 234672 249024 234678 249076
rect 336734 249024 336740 249076
rect 336792 249064 336798 249076
rect 538214 249064 538220 249076
rect 336792 249036 538220 249064
rect 336792 249024 336798 249036
rect 538214 249024 538220 249036
rect 538272 249024 538278 249076
rect 295610 248344 295616 248396
rect 295668 248384 295674 248396
rect 361758 248384 361764 248396
rect 295668 248356 361764 248384
rect 295668 248344 295674 248356
rect 361758 248344 361764 248356
rect 361816 248344 361822 248396
rect 297082 248276 297088 248328
rect 297140 248316 297146 248328
rect 363414 248316 363420 248328
rect 297140 248288 363420 248316
rect 297140 248276 297146 248288
rect 363414 248276 363420 248288
rect 363472 248276 363478 248328
rect 298094 248208 298100 248260
rect 298152 248248 298158 248260
rect 364610 248248 364616 248260
rect 298152 248220 364616 248248
rect 298152 248208 298158 248220
rect 364610 248208 364616 248220
rect 364668 248208 364674 248260
rect 292666 248140 292672 248192
rect 292724 248180 292730 248192
rect 359182 248180 359188 248192
rect 292724 248152 359188 248180
rect 292724 248140 292730 248152
rect 359182 248140 359188 248152
rect 359240 248140 359246 248192
rect 296990 248072 296996 248124
rect 297048 248112 297054 248124
rect 364426 248112 364432 248124
rect 297048 248084 364432 248112
rect 297048 248072 297054 248084
rect 364426 248072 364432 248084
rect 364484 248072 364490 248124
rect 296806 248004 296812 248056
rect 296864 248044 296870 248056
rect 364518 248044 364524 248056
rect 296864 248016 364524 248044
rect 296864 248004 296870 248016
rect 364518 248004 364524 248016
rect 364576 248004 364582 248056
rect 151906 247936 151912 247988
rect 151964 247976 151970 247988
rect 260926 247976 260932 247988
rect 151964 247948 260932 247976
rect 151964 247936 151970 247948
rect 260926 247936 260932 247948
rect 260984 247936 260990 247988
rect 292758 247936 292764 247988
rect 292816 247976 292822 247988
rect 360746 247976 360752 247988
rect 292816 247948 360752 247976
rect 292816 247936 292822 247948
rect 360746 247936 360752 247948
rect 360804 247936 360810 247988
rect 147674 247868 147680 247920
rect 147732 247908 147738 247920
rect 260834 247908 260840 247920
rect 147732 247880 260840 247908
rect 147732 247868 147738 247880
rect 260834 247868 260840 247880
rect 260892 247868 260898 247920
rect 292850 247868 292856 247920
rect 292908 247908 292914 247920
rect 362218 247908 362224 247920
rect 292908 247880 362224 247908
rect 292908 247868 292914 247880
rect 362218 247868 362224 247880
rect 362276 247868 362282 247920
rect 127066 247800 127072 247852
rect 127124 247840 127130 247852
rect 256786 247840 256792 247852
rect 127124 247812 256792 247840
rect 127124 247800 127130 247812
rect 256786 247800 256792 247812
rect 256844 247800 256850 247852
rect 293954 247800 293960 247852
rect 294012 247840 294018 247852
rect 368658 247840 368664 247852
rect 294012 247812 368664 247840
rect 294012 247800 294018 247812
rect 368658 247800 368664 247812
rect 368716 247800 368722 247852
rect 69106 247732 69112 247784
rect 69164 247772 69170 247784
rect 245654 247772 245660 247784
rect 69164 247744 245660 247772
rect 69164 247732 69170 247744
rect 245654 247732 245660 247744
rect 245712 247732 245718 247784
rect 288802 247732 288808 247784
rect 288860 247772 288866 247784
rect 367094 247772 367100 247784
rect 288860 247744 367100 247772
rect 288860 247732 288866 247744
rect 367094 247732 367100 247744
rect 367152 247732 367158 247784
rect 2774 247664 2780 247716
rect 2832 247704 2838 247716
rect 232130 247704 232136 247716
rect 2832 247676 232136 247704
rect 2832 247664 2838 247676
rect 232130 247664 232136 247676
rect 232188 247664 232194 247716
rect 288710 247664 288716 247716
rect 288768 247704 288774 247716
rect 368566 247704 368572 247716
rect 288768 247676 368572 247704
rect 288768 247664 288774 247676
rect 368566 247664 368572 247676
rect 368624 247664 368630 247716
rect 298186 247596 298192 247648
rect 298244 247636 298250 247648
rect 364334 247636 364340 247648
rect 298244 247608 364340 247636
rect 298244 247596 298250 247608
rect 364334 247596 364340 247608
rect 364392 247596 364398 247648
rect 291470 247528 291476 247580
rect 291528 247568 291534 247580
rect 356698 247568 356704 247580
rect 291528 247540 356704 247568
rect 291528 247528 291534 247540
rect 356698 247528 356704 247540
rect 356756 247528 356762 247580
rect 299658 247460 299664 247512
rect 299716 247500 299722 247512
rect 364794 247500 364800 247512
rect 299716 247472 364800 247500
rect 299716 247460 299722 247472
rect 364794 247460 364800 247472
rect 364852 247460 364858 247512
rect 291378 246644 291384 246696
rect 291436 246684 291442 246696
rect 366358 246684 366364 246696
rect 291436 246656 366364 246684
rect 291436 246644 291442 246656
rect 366358 246644 366364 246656
rect 366416 246644 366422 246696
rect 192478 246576 192484 246628
rect 192536 246616 192542 246628
rect 269574 246616 269580 246628
rect 192536 246588 269580 246616
rect 192536 246576 192542 246588
rect 269574 246576 269580 246588
rect 269632 246576 269638 246628
rect 310514 246576 310520 246628
rect 310572 246616 310578 246628
rect 405734 246616 405740 246628
rect 310572 246588 405740 246616
rect 310572 246576 310578 246588
rect 405734 246576 405740 246588
rect 405792 246576 405798 246628
rect 129734 246508 129740 246560
rect 129792 246548 129798 246560
rect 257154 246548 257160 246560
rect 129792 246520 257160 246548
rect 129792 246508 129798 246520
rect 257154 246508 257160 246520
rect 257212 246508 257218 246560
rect 331858 246508 331864 246560
rect 331916 246548 331922 246560
rect 430574 246548 430580 246560
rect 331916 246520 430580 246548
rect 331916 246508 331922 246520
rect 430574 246508 430580 246520
rect 430632 246508 430638 246560
rect 57974 246440 57980 246492
rect 58032 246480 58038 246492
rect 242986 246480 242992 246492
rect 58032 246452 242992 246480
rect 58032 246440 58038 246452
rect 242986 246440 242992 246452
rect 243044 246440 243050 246492
rect 314654 246440 314660 246492
rect 314712 246480 314718 246492
rect 423766 246480 423772 246492
rect 314712 246452 423772 246480
rect 314712 246440 314718 246452
rect 423766 246440 423772 246452
rect 423824 246440 423830 246492
rect 53834 246372 53840 246424
rect 53892 246412 53898 246424
rect 242894 246412 242900 246424
rect 53892 246384 242900 246412
rect 53892 246372 53898 246384
rect 242894 246372 242900 246384
rect 242952 246372 242958 246424
rect 317414 246372 317420 246424
rect 317472 246412 317478 246424
rect 440326 246412 440332 246424
rect 317472 246384 440332 246412
rect 317472 246372 317478 246384
rect 440326 246372 440332 246384
rect 440384 246372 440390 246424
rect 48958 246304 48964 246356
rect 49016 246344 49022 246356
rect 241514 246344 241520 246356
rect 49016 246316 241520 246344
rect 49016 246304 49022 246316
rect 241514 246304 241520 246316
rect 241572 246304 241578 246356
rect 328454 246304 328460 246356
rect 328512 246344 328518 246356
rect 496814 246344 496820 246356
rect 328512 246316 496820 246344
rect 328512 246304 328518 246316
rect 496814 246304 496820 246316
rect 496872 246304 496878 246356
rect 300946 245556 300952 245608
rect 301004 245596 301010 245608
rect 357434 245596 357440 245608
rect 301004 245568 357440 245596
rect 301004 245556 301010 245568
rect 357434 245556 357440 245568
rect 357492 245556 357498 245608
rect 357250 245488 357256 245540
rect 357308 245528 357314 245540
rect 369854 245528 369860 245540
rect 357308 245500 369860 245528
rect 357308 245488 357314 245500
rect 369854 245488 369860 245500
rect 369912 245488 369918 245540
rect 301038 245420 301044 245472
rect 301096 245460 301102 245472
rect 362126 245460 362132 245472
rect 301096 245432 362132 245460
rect 301096 245420 301102 245432
rect 362126 245420 362132 245432
rect 362184 245420 362190 245472
rect 299566 245352 299572 245404
rect 299624 245392 299630 245404
rect 363322 245392 363328 245404
rect 299624 245364 363328 245392
rect 299624 245352 299630 245364
rect 363322 245352 363328 245364
rect 363380 245352 363386 245404
rect 214834 245284 214840 245336
rect 214892 245324 214898 245336
rect 288618 245324 288624 245336
rect 214892 245296 288624 245324
rect 214892 245284 214898 245296
rect 288618 245284 288624 245296
rect 288676 245284 288682 245336
rect 295334 245284 295340 245336
rect 295392 245324 295398 245336
rect 360654 245324 360660 245336
rect 295392 245296 360660 245324
rect 295392 245284 295398 245296
rect 360654 245284 360660 245296
rect 360712 245284 360718 245336
rect 212994 245216 213000 245268
rect 213052 245256 213058 245268
rect 288526 245256 288532 245268
rect 213052 245228 288532 245256
rect 213052 245216 213058 245228
rect 288526 245216 288532 245228
rect 288584 245216 288590 245268
rect 292574 245216 292580 245268
rect 292632 245256 292638 245268
rect 357986 245256 357992 245268
rect 292632 245228 357992 245256
rect 292632 245216 292638 245228
rect 357986 245216 357992 245228
rect 358044 245216 358050 245268
rect 358078 245216 358084 245268
rect 358136 245256 358142 245268
rect 369946 245256 369952 245268
rect 358136 245228 369952 245256
rect 358136 245216 358142 245228
rect 369946 245216 369952 245228
rect 370004 245216 370010 245268
rect 135346 245148 135352 245200
rect 135404 245188 135410 245200
rect 253198 245188 253204 245200
rect 135404 245160 253204 245188
rect 135404 245148 135410 245160
rect 253198 245148 253204 245160
rect 253256 245148 253262 245200
rect 291286 245148 291292 245200
rect 291344 245188 291350 245200
rect 367186 245188 367192 245200
rect 291344 245160 367192 245188
rect 291344 245148 291350 245160
rect 367186 245148 367192 245160
rect 367244 245148 367250 245200
rect 132494 245080 132500 245132
rect 132552 245120 132558 245132
rect 257338 245120 257344 245132
rect 132552 245092 257344 245120
rect 132552 245080 132558 245092
rect 257338 245080 257344 245092
rect 257396 245080 257402 245132
rect 329834 245080 329840 245132
rect 329892 245120 329898 245132
rect 502334 245120 502340 245132
rect 329892 245092 502340 245120
rect 329892 245080 329898 245092
rect 502334 245080 502340 245092
rect 502392 245080 502398 245132
rect 6914 245012 6920 245064
rect 6972 245052 6978 245064
rect 233234 245052 233240 245064
rect 6972 245024 233240 245052
rect 6972 245012 6978 245024
rect 233234 245012 233240 245024
rect 233292 245012 233298 245064
rect 340966 245012 340972 245064
rect 341024 245052 341030 245064
rect 557534 245052 557540 245064
rect 341024 245024 557540 245052
rect 341024 245012 341030 245024
rect 557534 245012 557540 245024
rect 557592 245012 557598 245064
rect 4890 244944 4896 244996
rect 4948 244984 4954 244996
rect 232038 244984 232044 244996
rect 4948 244956 232044 244984
rect 4948 244944 4954 244956
rect 232038 244944 232044 244956
rect 232096 244944 232102 244996
rect 340874 244944 340880 244996
rect 340932 244984 340938 244996
rect 561674 244984 561680 244996
rect 340932 244956 561680 244984
rect 340932 244944 340938 244956
rect 561674 244944 561680 244956
rect 561732 244944 561738 244996
rect 2866 244876 2872 244928
rect 2924 244916 2930 244928
rect 231946 244916 231952 244928
rect 2924 244888 231952 244916
rect 2924 244876 2930 244888
rect 231946 244876 231952 244888
rect 232004 244876 232010 244928
rect 342254 244876 342260 244928
rect 342312 244916 342318 244928
rect 564526 244916 564532 244928
rect 342312 244888 564532 244916
rect 342312 244876 342318 244888
rect 564526 244876 564532 244888
rect 564584 244876 564590 244928
rect 357066 244808 357072 244860
rect 357124 244848 357130 244860
rect 364886 244848 364892 244860
rect 357124 244820 364892 244848
rect 357124 244808 357130 244820
rect 364886 244808 364892 244820
rect 364944 244808 364950 244860
rect 356974 244604 356980 244656
rect 357032 244644 357038 244656
rect 363690 244644 363696 244656
rect 357032 244616 363696 244644
rect 357032 244604 357038 244616
rect 363690 244604 363696 244616
rect 363748 244604 363754 244656
rect 357158 244468 357164 244520
rect 357216 244508 357222 244520
rect 362310 244508 362316 244520
rect 357216 244480 362316 244508
rect 357216 244468 357222 244480
rect 362310 244468 362316 244480
rect 362368 244468 362374 244520
rect 355318 244060 355324 244112
rect 355376 244100 355382 244112
rect 362402 244100 362408 244112
rect 355376 244072 362408 244100
rect 355376 244060 355382 244072
rect 362402 244060 362408 244072
rect 362460 244060 362466 244112
rect 355410 243992 355416 244044
rect 355468 244032 355474 244044
rect 359274 244032 359280 244044
rect 355468 244004 359280 244032
rect 355468 243992 355474 244004
rect 359274 243992 359280 244004
rect 359332 243992 359338 244044
rect 219158 243720 219164 243772
rect 219216 243760 219222 243772
rect 287330 243760 287336 243772
rect 219216 243732 287336 243760
rect 219216 243720 219222 243732
rect 287330 243720 287336 243732
rect 287388 243720 287394 243772
rect 289998 243720 290004 243772
rect 290056 243760 290062 243772
rect 358078 243760 358084 243772
rect 290056 243732 358084 243760
rect 290056 243720 290062 243732
rect 358078 243720 358084 243732
rect 358136 243720 358142 243772
rect 217226 243652 217232 243704
rect 217284 243692 217290 243704
rect 286042 243692 286048 243704
rect 217284 243664 286048 243692
rect 217284 243652 217290 243664
rect 286042 243652 286048 243664
rect 286100 243652 286106 243704
rect 289814 243652 289820 243704
rect 289872 243692 289878 243704
rect 360838 243692 360844 243704
rect 289872 243664 360844 243692
rect 289872 243652 289878 243664
rect 360838 243652 360844 243664
rect 360896 243652 360902 243704
rect 219250 243584 219256 243636
rect 219308 243624 219314 243636
rect 288894 243624 288900 243636
rect 219308 243596 288900 243624
rect 219308 243584 219314 243596
rect 288894 243584 288900 243596
rect 288952 243584 288958 243636
rect 289906 243584 289912 243636
rect 289964 243624 289970 243636
rect 363598 243624 363604 243636
rect 289964 243596 363604 243624
rect 289964 243584 289970 243596
rect 363598 243584 363604 243596
rect 363656 243584 363662 243636
rect 215754 243516 215760 243568
rect 215812 243556 215818 243568
rect 287422 243556 287428 243568
rect 215812 243528 287428 243556
rect 215812 243516 215818 243528
rect 287422 243516 287428 243528
rect 287480 243516 287486 243568
rect 291194 243516 291200 243568
rect 291252 243556 291258 243568
rect 364978 243556 364984 243568
rect 291252 243528 364984 243556
rect 291252 243516 291258 243528
rect 364978 243516 364984 243528
rect 365036 243516 365042 243568
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 210418 215268 210424 215280
rect 3384 215240 210424 215268
rect 3384 215228 3390 215240
rect 210418 215228 210424 215240
rect 210476 215228 210482 215280
rect 214374 195236 214380 195288
rect 214432 195276 214438 195288
rect 217318 195276 217324 195288
rect 214432 195248 217324 195276
rect 214432 195236 214438 195248
rect 217318 195236 217324 195248
rect 217376 195236 217382 195288
rect 215754 193128 215760 193180
rect 215812 193168 215818 193180
rect 217410 193168 217416 193180
rect 215812 193140 217416 193168
rect 215812 193128 215818 193140
rect 217410 193128 217416 193140
rect 217468 193128 217474 193180
rect 210510 193060 210516 193112
rect 210568 193100 210574 193112
rect 216674 193100 216680 193112
rect 210568 193072 216680 193100
rect 210568 193060 210574 193072
rect 216674 193060 216680 193072
rect 216732 193060 216738 193112
rect 215846 189252 215852 189304
rect 215904 189292 215910 189304
rect 218606 189292 218612 189304
rect 215904 189264 218612 189292
rect 215904 189252 215910 189264
rect 218606 189252 218612 189264
rect 218664 189252 218670 189304
rect 210602 188980 210608 189032
rect 210660 189020 210666 189032
rect 216674 189020 216680 189032
rect 210660 188992 216680 189020
rect 210660 188980 210666 188992
rect 216674 188980 216680 188992
rect 216732 188980 216738 189032
rect 212994 169532 213000 169584
rect 213052 169572 213058 169584
rect 217502 169572 217508 169584
rect 213052 169544 217508 169572
rect 213052 169532 213058 169544
rect 217502 169532 217508 169544
rect 217560 169532 217566 169584
rect 351914 159672 351920 159724
rect 351972 159712 351978 159724
rect 357894 159712 357900 159724
rect 351972 159684 357900 159712
rect 351972 159672 351978 159684
rect 357894 159672 357900 159684
rect 357952 159672 357958 159724
rect 213086 159604 213092 159656
rect 213144 159644 213150 159656
rect 256694 159644 256700 159656
rect 213144 159616 256700 159644
rect 213144 159604 213150 159616
rect 256694 159604 256700 159616
rect 256752 159604 256758 159656
rect 325878 159604 325884 159656
rect 325936 159644 325942 159656
rect 357802 159644 357808 159656
rect 325936 159616 357808 159644
rect 325936 159604 325942 159616
rect 357802 159604 357808 159616
rect 357860 159604 357866 159656
rect 217870 159536 217876 159588
rect 217928 159576 217934 159588
rect 263594 159576 263600 159588
rect 217928 159548 263600 159576
rect 217928 159536 217934 159548
rect 263594 159536 263600 159548
rect 263652 159536 263658 159588
rect 313274 159536 313280 159588
rect 313332 159576 313338 159588
rect 356790 159576 356796 159588
rect 313332 159548 356796 159576
rect 313332 159536 313338 159548
rect 356790 159536 356796 159548
rect 356848 159536 356854 159588
rect 214466 159468 214472 159520
rect 214524 159508 214530 159520
rect 260834 159508 260840 159520
rect 214524 159480 260840 159508
rect 214524 159468 214530 159480
rect 260834 159468 260840 159480
rect 260892 159468 260898 159520
rect 310974 159468 310980 159520
rect 311032 159508 311038 159520
rect 358998 159508 359004 159520
rect 311032 159480 359004 159508
rect 311032 159468 311038 159480
rect 358998 159468 359004 159480
rect 359056 159468 359062 159520
rect 217778 159400 217784 159452
rect 217836 159440 217842 159452
rect 264974 159440 264980 159452
rect 217836 159412 264980 159440
rect 217836 159400 217842 159412
rect 264974 159400 264980 159412
rect 265032 159400 265038 159452
rect 291102 159400 291108 159452
rect 291160 159440 291166 159452
rect 359090 159440 359096 159452
rect 291160 159412 359096 159440
rect 291160 159400 291166 159412
rect 359090 159400 359096 159412
rect 359148 159400 359154 159452
rect 216122 159332 216128 159384
rect 216180 159372 216186 159384
rect 284386 159372 284392 159384
rect 216180 159344 284392 159372
rect 216180 159332 216186 159344
rect 284386 159332 284392 159344
rect 284444 159332 284450 159384
rect 285674 159332 285680 159384
rect 285732 159372 285738 159384
rect 360562 159372 360568 159384
rect 285732 159344 360568 159372
rect 285732 159332 285738 159344
rect 360562 159332 360568 159344
rect 360620 159332 360626 159384
rect 363230 159236 363236 159248
rect 355060 159208 363236 159236
rect 279234 159128 279240 159180
rect 279292 159168 279298 159180
rect 355060 159168 355088 159208
rect 363230 159196 363236 159208
rect 363288 159196 363294 159248
rect 363138 159168 363144 159180
rect 279292 159140 355088 159168
rect 355152 159140 363144 159168
rect 279292 159128 279298 159140
rect 278130 159060 278136 159112
rect 278188 159100 278194 159112
rect 355152 159100 355180 159140
rect 363138 159128 363144 159140
rect 363196 159128 363202 159180
rect 278188 159072 355180 159100
rect 278188 159060 278194 159072
rect 355226 159060 355232 159112
rect 355284 159100 355290 159112
rect 361942 159100 361948 159112
rect 355284 159072 361948 159100
rect 355284 159060 355290 159072
rect 361942 159060 361948 159072
rect 362000 159060 362006 159112
rect 277026 158992 277032 159044
rect 277084 159032 277090 159044
rect 362034 159032 362040 159044
rect 277084 159004 362040 159032
rect 277084 158992 277090 159004
rect 362034 158992 362040 159004
rect 362092 158992 362098 159044
rect 273346 158924 273352 158976
rect 273404 158964 273410 158976
rect 360470 158964 360476 158976
rect 273404 158936 360476 158964
rect 273404 158924 273410 158936
rect 360470 158924 360476 158936
rect 360528 158924 360534 158976
rect 275830 158856 275836 158908
rect 275888 158896 275894 158908
rect 355226 158896 355232 158908
rect 275888 158868 355232 158896
rect 275888 158856 275894 158868
rect 355226 158856 355232 158868
rect 355284 158856 355290 158908
rect 361022 158896 361028 158908
rect 355336 158868 361028 158896
rect 274450 158788 274456 158840
rect 274508 158828 274514 158840
rect 355336 158828 355364 158868
rect 361022 158856 361028 158868
rect 361080 158856 361086 158908
rect 359366 158828 359372 158840
rect 274508 158800 355364 158828
rect 355428 158800 359372 158828
rect 274508 158788 274514 158800
rect 211890 158720 211896 158772
rect 211948 158760 211954 158772
rect 239582 158760 239588 158772
rect 211948 158732 239588 158760
rect 211948 158720 211954 158732
rect 239582 158720 239588 158732
rect 239640 158720 239646 158772
rect 261110 158720 261116 158772
rect 261168 158760 261174 158772
rect 355428 158760 355456 158800
rect 359366 158788 359372 158800
rect 359424 158788 359430 158840
rect 357618 158760 357624 158772
rect 261168 158732 355456 158760
rect 356164 158732 357624 158760
rect 261168 158720 261174 158732
rect 213362 158652 213368 158704
rect 213420 158692 213426 158704
rect 238110 158692 238116 158704
rect 213420 158664 238116 158692
rect 213420 158652 213426 158664
rect 238110 158652 238116 158664
rect 238168 158652 238174 158704
rect 269942 158652 269948 158704
rect 270000 158692 270006 158704
rect 291102 158692 291108 158704
rect 270000 158664 291108 158692
rect 270000 158652 270006 158664
rect 291102 158652 291108 158664
rect 291160 158652 291166 158704
rect 295978 158652 295984 158704
rect 296036 158692 296042 158704
rect 356164 158692 356192 158732
rect 357618 158720 357624 158732
rect 357676 158720 357682 158772
rect 296036 158664 356192 158692
rect 296036 158652 296042 158664
rect 214558 158584 214564 158636
rect 214616 158624 214622 158636
rect 233234 158624 233240 158636
rect 214616 158596 233240 158624
rect 214616 158584 214622 158596
rect 233234 158584 233240 158596
rect 233292 158584 233298 158636
rect 315850 158584 315856 158636
rect 315908 158624 315914 158636
rect 361850 158624 361856 158636
rect 315908 158596 361856 158624
rect 315908 158584 315914 158596
rect 361850 158584 361856 158596
rect 361908 158584 361914 158636
rect 218974 158516 218980 158568
rect 219032 158556 219038 158568
rect 238754 158556 238760 158568
rect 219032 158528 238760 158556
rect 219032 158516 219038 158528
rect 238754 158516 238760 158528
rect 238812 158516 238818 158568
rect 272242 158516 272248 158568
rect 272300 158556 272306 158568
rect 285674 158556 285680 158568
rect 272300 158528 285680 158556
rect 272300 158516 272306 158528
rect 285674 158516 285680 158528
rect 285732 158516 285738 158568
rect 293586 158516 293592 158568
rect 293644 158556 293650 158568
rect 351914 158556 351920 158568
rect 293644 158528 351920 158556
rect 293644 158516 293650 158528
rect 351914 158516 351920 158528
rect 351972 158516 351978 158568
rect 211982 158448 211988 158500
rect 212040 158488 212046 158500
rect 237374 158488 237380 158500
rect 212040 158460 237380 158488
rect 212040 158448 212046 158460
rect 237374 158448 237380 158460
rect 237432 158448 237438 158500
rect 298554 158448 298560 158500
rect 298612 158488 298618 158500
rect 358354 158488 358360 158500
rect 298612 158460 358360 158488
rect 298612 158448 298618 158460
rect 358354 158448 358360 158460
rect 358412 158448 358418 158500
rect 216398 158380 216404 158432
rect 216456 158420 216462 158432
rect 242986 158420 242992 158432
rect 216456 158392 242992 158420
rect 216456 158380 216462 158392
rect 242986 158380 242992 158392
rect 243044 158380 243050 158432
rect 300946 158380 300952 158432
rect 301004 158420 301010 158432
rect 358906 158420 358912 158432
rect 301004 158392 358912 158420
rect 301004 158380 301010 158392
rect 358906 158380 358912 158392
rect 358964 158380 358970 158432
rect 213270 158312 213276 158364
rect 213328 158352 213334 158364
rect 241514 158352 241520 158364
rect 213328 158324 241520 158352
rect 213328 158312 213334 158324
rect 241514 158312 241520 158324
rect 241572 158312 241578 158364
rect 303522 158312 303528 158364
rect 303580 158352 303586 158364
rect 358170 158352 358176 158364
rect 303580 158324 358176 158352
rect 303580 158312 303586 158324
rect 358170 158312 358176 158324
rect 358228 158312 358234 158364
rect 216490 158244 216496 158296
rect 216548 158284 216554 158296
rect 245654 158284 245660 158296
rect 216548 158256 245660 158284
rect 216548 158244 216554 158256
rect 245654 158244 245660 158256
rect 245712 158244 245718 158296
rect 306098 158244 306104 158296
rect 306156 158284 306162 158296
rect 358262 158284 358268 158296
rect 306156 158256 358268 158284
rect 306156 158244 306162 158256
rect 358262 158244 358268 158256
rect 358320 158244 358326 158296
rect 214650 158176 214656 158228
rect 214708 158216 214714 158228
rect 247034 158216 247040 158228
rect 214708 158188 247040 158216
rect 214708 158176 214714 158188
rect 247034 158176 247040 158188
rect 247092 158176 247098 158228
rect 308674 158176 308680 158228
rect 308732 158216 308738 158228
rect 360378 158216 360384 158228
rect 308732 158188 360384 158216
rect 308732 158176 308738 158188
rect 360378 158176 360384 158188
rect 360436 158176 360442 158228
rect 215938 158108 215944 158160
rect 215996 158148 216002 158160
rect 248414 158148 248420 158160
rect 215996 158120 248420 158148
rect 215996 158108 216002 158120
rect 248414 158108 248420 158120
rect 248472 158108 248478 158160
rect 268746 158108 268752 158160
rect 268804 158148 268810 158160
rect 310974 158148 310980 158160
rect 268804 158120 310980 158148
rect 268804 158108 268810 158120
rect 310974 158108 310980 158120
rect 311032 158108 311038 158160
rect 311066 158108 311072 158160
rect 311124 158148 311130 158160
rect 360286 158148 360292 158160
rect 311124 158120 360292 158148
rect 311124 158108 311130 158120
rect 360286 158108 360292 158120
rect 360344 158108 360350 158160
rect 216306 158040 216312 158092
rect 216364 158080 216370 158092
rect 249794 158080 249800 158092
rect 216364 158052 249800 158080
rect 216364 158040 216370 158052
rect 249794 158040 249800 158052
rect 249852 158040 249858 158092
rect 288250 158040 288256 158092
rect 288308 158080 288314 158092
rect 313274 158080 313280 158092
rect 288308 158052 313280 158080
rect 288308 158040 288314 158052
rect 313274 158040 313280 158052
rect 313332 158040 313338 158092
rect 313458 158040 313464 158092
rect 313516 158080 313522 158092
rect 359642 158080 359648 158092
rect 313516 158052 359648 158080
rect 313516 158040 313522 158052
rect 359642 158040 359648 158052
rect 359700 158040 359706 158092
rect 218698 157972 218704 158024
rect 218756 158012 218762 158024
rect 252554 158012 252560 158024
rect 218756 157984 252560 158012
rect 218756 157972 218762 157984
rect 252554 157972 252560 157984
rect 252612 157972 252618 158024
rect 318610 157972 318616 158024
rect 318668 158012 318674 158024
rect 359550 158012 359556 158024
rect 318668 157984 359556 158012
rect 318668 157972 318674 157984
rect 359550 157972 359556 157984
rect 359608 157972 359614 158024
rect 212074 157904 212080 157956
rect 212132 157944 212138 157956
rect 230474 157944 230480 157956
rect 212132 157916 230480 157944
rect 212132 157904 212138 157916
rect 230474 157904 230480 157916
rect 230532 157904 230538 157956
rect 323394 157904 323400 157956
rect 323452 157944 323458 157956
rect 363046 157944 363052 157956
rect 323452 157916 363052 157944
rect 323452 157904 323458 157916
rect 363046 157904 363052 157916
rect 363104 157904 363110 157956
rect 216214 157836 216220 157888
rect 216272 157876 216278 157888
rect 229094 157876 229100 157888
rect 216272 157848 229100 157876
rect 216272 157836 216278 157848
rect 229094 157836 229100 157848
rect 229152 157836 229158 157888
rect 321002 157836 321008 157888
rect 321060 157876 321066 157888
rect 359458 157876 359464 157888
rect 321060 157848 359464 157876
rect 321060 157836 321066 157848
rect 359458 157836 359464 157848
rect 359516 157836 359522 157888
rect 219066 157768 219072 157820
rect 219124 157808 219130 157820
rect 231854 157808 231860 157820
rect 219124 157780 231860 157808
rect 219124 157768 219130 157780
rect 231854 157768 231860 157780
rect 231912 157768 231918 157820
rect 265434 157768 265440 157820
rect 265492 157808 265498 157820
rect 325878 157808 325884 157820
rect 265492 157780 325884 157808
rect 265492 157768 265498 157780
rect 325878 157768 325884 157780
rect 325936 157768 325942 157820
rect 325970 157768 325976 157820
rect 326028 157808 326034 157820
rect 360930 157808 360936 157820
rect 326028 157780 360936 157808
rect 326028 157768 326034 157780
rect 360930 157768 360936 157780
rect 360988 157768 360994 157820
rect 242434 157292 242440 157344
rect 242492 157332 242498 157344
rect 372706 157332 372712 157344
rect 242492 157304 372712 157332
rect 242492 157292 242498 157304
rect 372706 157292 372712 157304
rect 372764 157292 372770 157344
rect 244642 157224 244648 157276
rect 244700 157264 244706 157276
rect 370038 157264 370044 157276
rect 244700 157236 370044 157264
rect 244700 157224 244706 157236
rect 370038 157224 370044 157236
rect 370096 157224 370102 157276
rect 248322 157156 248328 157208
rect 248380 157196 248386 157208
rect 369302 157196 369308 157208
rect 248380 157168 369308 157196
rect 248380 157156 248386 157168
rect 369302 157156 369308 157168
rect 369360 157156 369366 157208
rect 245562 157088 245568 157140
rect 245620 157128 245626 157140
rect 363782 157128 363788 157140
rect 245620 157100 363788 157128
rect 245620 157088 245626 157100
rect 363782 157088 363788 157100
rect 363840 157088 363846 157140
rect 252370 157020 252376 157072
rect 252428 157060 252434 157072
rect 369210 157060 369216 157072
rect 252428 157032 369216 157060
rect 252428 157020 252434 157032
rect 369210 157020 369216 157032
rect 369268 157020 369274 157072
rect 255866 156952 255872 157004
rect 255924 156992 255930 157004
rect 367278 156992 367284 157004
rect 255924 156964 367284 156992
rect 255924 156952 255930 156964
rect 367278 156952 367284 156964
rect 367336 156952 367342 157004
rect 257246 156884 257252 156936
rect 257304 156924 257310 156936
rect 367370 156924 367376 156936
rect 257304 156896 367376 156924
rect 257304 156884 257310 156896
rect 367370 156884 367376 156896
rect 367428 156884 367434 156936
rect 261754 156816 261760 156868
rect 261812 156856 261818 156868
rect 370130 156856 370136 156868
rect 261812 156828 370136 156856
rect 261812 156816 261818 156828
rect 370130 156816 370136 156828
rect 370188 156816 370194 156868
rect 265986 156748 265992 156800
rect 266044 156788 266050 156800
rect 372890 156788 372896 156800
rect 266044 156760 372896 156788
rect 266044 156748 266050 156760
rect 372890 156748 372896 156760
rect 372948 156748 372954 156800
rect 266538 156680 266544 156732
rect 266596 156720 266602 156732
rect 368842 156720 368848 156732
rect 266596 156692 368848 156720
rect 266596 156680 266602 156692
rect 368842 156680 368848 156692
rect 368900 156680 368906 156732
rect 270954 156612 270960 156664
rect 271012 156652 271018 156664
rect 372798 156652 372804 156664
rect 271012 156624 372804 156652
rect 271012 156612 271018 156624
rect 372798 156612 372804 156624
rect 372856 156612 372862 156664
rect 276106 156544 276112 156596
rect 276164 156584 276170 156596
rect 371786 156584 371792 156596
rect 276164 156556 371792 156584
rect 276164 156544 276170 156556
rect 371786 156544 371792 156556
rect 371844 156544 371850 156596
rect 281074 156476 281080 156528
rect 281132 156516 281138 156528
rect 371878 156516 371884 156528
rect 281132 156488 371884 156516
rect 281132 156476 281138 156488
rect 371878 156476 371884 156488
rect 371936 156476 371942 156528
rect 217962 156408 217968 156460
rect 218020 156448 218026 156460
rect 285674 156448 285680 156460
rect 218020 156420 285680 156448
rect 218020 156408 218026 156420
rect 285674 156408 285680 156420
rect 285732 156408 285738 156460
rect 291010 156408 291016 156460
rect 291068 156448 291074 156460
rect 371694 156448 371700 156460
rect 291068 156420 371700 156448
rect 291068 156408 291074 156420
rect 371694 156408 371700 156420
rect 371752 156408 371758 156460
rect 241422 155864 241428 155916
rect 241480 155904 241486 155916
rect 374178 155904 374184 155916
rect 241480 155876 374184 155904
rect 241480 155864 241486 155876
rect 374178 155864 374184 155876
rect 374236 155864 374242 155916
rect 246666 155796 246672 155848
rect 246724 155836 246730 155848
rect 370222 155836 370228 155848
rect 246724 155808 370228 155836
rect 246724 155796 246730 155808
rect 370222 155796 370228 155808
rect 370280 155796 370286 155848
rect 251082 155728 251088 155780
rect 251140 155768 251146 155780
rect 371970 155768 371976 155780
rect 251140 155740 371976 155768
rect 251140 155728 251146 155740
rect 371970 155728 371976 155740
rect 372028 155728 372034 155780
rect 247954 155660 247960 155712
rect 248012 155700 248018 155712
rect 368934 155700 368940 155712
rect 248012 155672 368940 155700
rect 248012 155660 248018 155672
rect 368934 155660 368940 155672
rect 368992 155660 368998 155712
rect 248690 155592 248696 155644
rect 248748 155632 248754 155644
rect 370314 155632 370320 155644
rect 248748 155604 370320 155632
rect 248748 155592 248754 155604
rect 370314 155592 370320 155604
rect 370372 155592 370378 155644
rect 250438 155524 250444 155576
rect 250496 155564 250502 155576
rect 369026 155564 369032 155576
rect 250496 155536 369032 155564
rect 250496 155524 250502 155536
rect 369026 155524 369032 155536
rect 369084 155524 369090 155576
rect 252462 155456 252468 155508
rect 252520 155496 252526 155508
rect 370406 155496 370412 155508
rect 252520 155468 370412 155496
rect 252520 155456 252526 155468
rect 370406 155456 370412 155468
rect 370464 155456 370470 155508
rect 218790 155388 218796 155440
rect 218848 155428 218854 155440
rect 251174 155428 251180 155440
rect 218848 155400 251180 155428
rect 218848 155388 218854 155400
rect 251174 155388 251180 155400
rect 251232 155388 251238 155440
rect 253474 155388 253480 155440
rect 253532 155428 253538 155440
rect 365070 155428 365076 155440
rect 253532 155400 365076 155428
rect 253532 155388 253538 155400
rect 365070 155388 365076 155400
rect 365128 155388 365134 155440
rect 210786 155320 210792 155372
rect 210844 155360 210850 155372
rect 267734 155360 267740 155372
rect 210844 155332 267740 155360
rect 210844 155320 210850 155332
rect 267734 155320 267740 155332
rect 267792 155320 267798 155372
rect 268378 155320 268384 155372
rect 268436 155360 268442 155372
rect 374270 155360 374276 155372
rect 268436 155332 374276 155360
rect 268436 155320 268442 155332
rect 374270 155320 374276 155332
rect 374328 155320 374334 155372
rect 212166 155252 212172 155304
rect 212224 155292 212230 155304
rect 271874 155292 271880 155304
rect 212224 155264 271880 155292
rect 212224 155252 212230 155264
rect 271874 155252 271880 155264
rect 271932 155252 271938 155304
rect 273714 155252 273720 155304
rect 273772 155292 273778 155304
rect 371510 155292 371516 155304
rect 273772 155264 371516 155292
rect 273772 155252 273778 155264
rect 371510 155252 371516 155264
rect 371568 155252 371574 155304
rect 210694 155184 210700 155236
rect 210752 155224 210758 155236
rect 270494 155224 270500 155236
rect 210752 155196 270500 155224
rect 210752 155184 210758 155196
rect 270494 155184 270500 155196
rect 270552 155184 270558 155236
rect 271322 155184 271328 155236
rect 271380 155224 271386 155236
rect 368750 155224 368756 155236
rect 271380 155196 368756 155224
rect 271380 155184 271386 155196
rect 368750 155184 368756 155196
rect 368808 155184 368814 155236
rect 216030 155116 216036 155168
rect 216088 155156 216094 155168
rect 277394 155156 277400 155168
rect 216088 155128 277400 155156
rect 216088 155116 216094 155128
rect 277394 155116 277400 155128
rect 277452 155116 277458 155168
rect 278498 155116 278504 155168
rect 278556 155156 278562 155168
rect 371418 155156 371424 155168
rect 278556 155128 371424 155156
rect 278556 155116 278562 155128
rect 371418 155116 371424 155128
rect 371476 155116 371482 155168
rect 214742 155048 214748 155100
rect 214800 155088 214806 155100
rect 282914 155088 282920 155100
rect 214800 155060 282920 155088
rect 214800 155048 214806 155060
rect 282914 155048 282920 155060
rect 282972 155048 282978 155100
rect 283650 155048 283656 155100
rect 283708 155088 283714 155100
rect 371326 155088 371332 155100
rect 283708 155060 371332 155088
rect 283708 155048 283714 155060
rect 371326 155048 371332 155060
rect 371384 155048 371390 155100
rect 217226 154980 217232 155032
rect 217284 155020 217290 155032
rect 278774 155020 278780 155032
rect 217284 154992 278780 155020
rect 217284 154980 217290 154992
rect 278774 154980 278780 154992
rect 278832 154980 278838 155032
rect 256234 154504 256240 154556
rect 256292 154544 256298 154556
rect 367646 154544 367652 154556
rect 256292 154516 367652 154544
rect 256292 154504 256298 154516
rect 367646 154504 367652 154516
rect 367704 154504 367710 154556
rect 263686 154436 263692 154488
rect 263744 154476 263750 154488
rect 371602 154476 371608 154488
rect 263744 154448 371608 154476
rect 263744 154436 263750 154448
rect 371602 154436 371608 154448
rect 371660 154436 371666 154488
rect 286042 154368 286048 154420
rect 286100 154408 286106 154420
rect 370590 154408 370596 154420
rect 286100 154380 370596 154408
rect 286100 154368 286106 154380
rect 370590 154368 370596 154380
rect 370648 154368 370654 154420
rect 218606 152600 218612 152652
rect 218664 152640 218670 152652
rect 276106 152640 276112 152652
rect 218664 152612 276112 152640
rect 218664 152600 218670 152612
rect 276106 152600 276112 152612
rect 276164 152600 276170 152652
rect 212258 152532 212264 152584
rect 212316 152572 212322 152584
rect 273254 152572 273260 152584
rect 212316 152544 273260 152572
rect 212316 152532 212322 152544
rect 273254 152532 273260 152544
rect 273312 152532 273318 152584
rect 213454 152464 213460 152516
rect 213512 152504 213518 152516
rect 288434 152504 288440 152516
rect 213512 152476 288440 152504
rect 213512 152464 213518 152476
rect 288434 152464 288440 152476
rect 288492 152464 288498 152516
rect 3510 150356 3516 150408
rect 3568 150396 3574 150408
rect 43438 150396 43444 150408
rect 3568 150368 43444 150396
rect 3568 150356 3574 150368
rect 43438 150356 43444 150368
rect 43496 150356 43502 150408
rect 3510 137912 3516 137964
rect 3568 137952 3574 137964
rect 180058 137952 180064 137964
rect 3568 137924 180064 137952
rect 3568 137912 3574 137924
rect 180058 137912 180064 137924
rect 180116 137912 180122 137964
rect 143534 11704 143540 11756
rect 143592 11744 143598 11756
rect 144730 11744 144736 11756
rect 143592 11716 144736 11744
rect 143592 11704 143598 11716
rect 144730 11704 144736 11716
rect 144788 11704 144794 11756
rect 168374 11704 168380 11756
rect 168432 11744 168438 11756
rect 169570 11744 169576 11756
rect 168432 11716 169576 11744
rect 168432 11704 168438 11716
rect 169570 11704 169576 11716
rect 169628 11704 169634 11756
rect 201494 11704 201500 11756
rect 201552 11744 201558 11756
rect 202690 11744 202696 11756
rect 201552 11716 202696 11744
rect 201552 11704 201558 11716
rect 202690 11704 202696 11716
rect 202748 11704 202754 11756
rect 234614 11704 234620 11756
rect 234672 11744 234678 11756
rect 235810 11744 235816 11756
rect 234672 11716 235816 11744
rect 234672 11704 234678 11716
rect 235810 11704 235816 11716
rect 235868 11704 235874 11756
rect 151722 9596 151728 9648
rect 151780 9636 151786 9648
rect 153010 9636 153016 9648
rect 151780 9608 153016 9636
rect 151780 9596 151786 9608
rect 153010 9596 153016 9608
rect 153068 9596 153074 9648
rect 209682 9596 209688 9648
rect 209740 9636 209746 9648
rect 210970 9636 210976 9648
rect 209740 9608 210976 9636
rect 209740 9596 209746 9608
rect 210970 9596 210976 9608
rect 211028 9596 211034 9648
rect 300762 9596 300768 9648
rect 300820 9636 300826 9648
rect 360838 9636 360844 9648
rect 300820 9608 360844 9636
rect 300820 9596 300826 9608
rect 360838 9596 360844 9608
rect 360896 9596 360902 9648
rect 301958 9528 301964 9580
rect 302016 9568 302022 9580
rect 362402 9568 362408 9580
rect 302016 9540 362408 9568
rect 302016 9528 302022 9540
rect 362402 9528 362408 9540
rect 362460 9528 362466 9580
rect 309042 9460 309048 9512
rect 309100 9500 309106 9512
rect 369854 9500 369860 9512
rect 309100 9472 369860 9500
rect 309100 9460 309106 9472
rect 369854 9460 369860 9472
rect 369912 9460 369918 9512
rect 306742 9392 306748 9444
rect 306800 9432 306806 9444
rect 368474 9432 368480 9444
rect 306800 9404 368480 9432
rect 306800 9392 306806 9404
rect 368474 9392 368480 9404
rect 368532 9392 368538 9444
rect 305546 9324 305552 9376
rect 305604 9364 305610 9376
rect 367186 9364 367192 9376
rect 305604 9336 367192 9364
rect 305604 9324 305610 9336
rect 367186 9324 367192 9336
rect 367244 9324 367250 9376
rect 304350 9256 304356 9308
rect 304408 9296 304414 9308
rect 366358 9296 366364 9308
rect 304408 9268 366364 9296
rect 304408 9256 304414 9268
rect 366358 9256 366364 9268
rect 366416 9256 366422 9308
rect 303154 9188 303160 9240
rect 303212 9228 303218 9240
rect 364978 9228 364984 9240
rect 303212 9200 364984 9228
rect 303212 9188 303218 9200
rect 364978 9188 364984 9200
rect 365036 9188 365042 9240
rect 296070 9120 296076 9172
rect 296128 9160 296134 9172
rect 358078 9160 358084 9172
rect 296128 9132 358084 9160
rect 296128 9120 296134 9132
rect 358078 9120 358084 9132
rect 358136 9120 358142 9172
rect 299658 9052 299664 9104
rect 299716 9092 299722 9104
rect 362310 9092 362316 9104
rect 299716 9064 362316 9092
rect 299716 9052 299722 9064
rect 362310 9052 362316 9064
rect 362368 9052 362374 9104
rect 294874 8984 294880 9036
rect 294932 9024 294938 9036
rect 369946 9024 369952 9036
rect 294932 8996 369952 9024
rect 294932 8984 294938 8996
rect 369946 8984 369952 8996
rect 370004 8984 370010 9036
rect 293678 8916 293684 8968
rect 293736 8956 293742 8968
rect 368566 8956 368572 8968
rect 293736 8928 368572 8956
rect 293736 8916 293742 8928
rect 368566 8916 368572 8928
rect 368624 8916 368630 8968
rect 298462 8848 298468 8900
rect 298520 8888 298526 8900
rect 359274 8888 359280 8900
rect 298520 8860 359280 8888
rect 298520 8848 298526 8860
rect 359274 8848 359280 8860
rect 359332 8848 359338 8900
rect 312630 8780 312636 8832
rect 312688 8820 312694 8832
rect 360746 8820 360752 8832
rect 312688 8792 360752 8820
rect 312688 8780 312694 8792
rect 360746 8780 360752 8792
rect 360804 8780 360810 8832
rect 316218 8712 316224 8764
rect 316276 8752 316282 8764
rect 363506 8752 363512 8764
rect 316276 8724 363512 8752
rect 316276 8712 316282 8724
rect 363506 8712 363512 8724
rect 363564 8712 363570 8764
rect 330386 6808 330392 6860
rect 330444 6848 330450 6860
rect 363414 6848 363420 6860
rect 330444 6820 363420 6848
rect 330444 6808 330450 6820
rect 363414 6808 363420 6820
rect 363472 6808 363478 6860
rect 333882 6740 333888 6792
rect 333940 6780 333946 6792
rect 366266 6780 366272 6792
rect 333940 6752 366272 6780
rect 333940 6740 333946 6752
rect 366266 6740 366272 6752
rect 366324 6740 366330 6792
rect 323302 6672 323308 6724
rect 323360 6712 323366 6724
rect 357526 6712 357532 6724
rect 323360 6684 357532 6712
rect 323360 6672 323366 6684
rect 357526 6672 357532 6684
rect 357584 6672 357590 6724
rect 313826 6604 313832 6656
rect 313884 6644 313890 6656
rect 360194 6644 360200 6656
rect 313884 6616 360200 6644
rect 313884 6604 313890 6616
rect 360194 6604 360200 6616
rect 360252 6604 360258 6656
rect 319714 6536 319720 6588
rect 319772 6576 319778 6588
rect 365990 6576 365996 6588
rect 319772 6548 365996 6576
rect 319772 6536 319778 6548
rect 365990 6536 365996 6548
rect 366048 6536 366054 6588
rect 318518 6468 318524 6520
rect 318576 6508 318582 6520
rect 364886 6508 364892 6520
rect 318576 6480 364892 6508
rect 318576 6468 318582 6480
rect 364886 6468 364892 6480
rect 364944 6468 364950 6520
rect 317322 6400 317328 6452
rect 317380 6440 317386 6452
rect 363690 6440 363696 6452
rect 317380 6412 363696 6440
rect 317380 6400 317386 6412
rect 363690 6400 363696 6412
rect 363748 6400 363754 6452
rect 315022 6332 315028 6384
rect 315080 6372 315086 6384
rect 362218 6372 362224 6384
rect 315080 6344 362224 6372
rect 315080 6332 315086 6344
rect 362218 6332 362224 6344
rect 362276 6332 362282 6384
rect 311434 6264 311440 6316
rect 311492 6304 311498 6316
rect 359182 6304 359188 6316
rect 311492 6276 359188 6304
rect 311492 6264 311498 6276
rect 359182 6264 359188 6276
rect 359240 6264 359246 6316
rect 310238 6196 310244 6248
rect 310296 6236 310302 6248
rect 357986 6236 357992 6248
rect 310296 6208 357992 6236
rect 310296 6196 310302 6208
rect 357986 6196 357992 6208
rect 358044 6196 358050 6248
rect 292574 6128 292580 6180
rect 292632 6168 292638 6180
rect 367094 6168 367100 6180
rect 292632 6140 367100 6168
rect 292632 6128 292638 6140
rect 367094 6128 367100 6140
rect 367152 6128 367158 6180
rect 326798 6060 326804 6112
rect 326856 6100 326862 6112
rect 358814 6100 358820 6112
rect 326856 6072 358820 6100
rect 326856 6060 326862 6072
rect 358814 6060 358820 6072
rect 358872 6060 358878 6112
rect 337470 5992 337476 6044
rect 337528 6032 337534 6044
rect 366082 6032 366088 6044
rect 337528 6004 366088 6032
rect 337528 5992 337534 6004
rect 366082 5992 366088 6004
rect 366140 5992 366146 6044
rect 340966 5924 340972 5976
rect 341024 5964 341030 5976
rect 365898 5964 365904 5976
rect 341024 5936 365904 5964
rect 341024 5924 341030 5936
rect 365898 5924 365904 5936
rect 365956 5924 365962 5976
rect 220556 4168 220860 4196
rect 6454 4088 6460 4140
rect 6512 4128 6518 4140
rect 7558 4128 7564 4140
rect 6512 4100 7564 4128
rect 6512 4088 6518 4100
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 15930 4088 15936 4140
rect 15988 4128 15994 4140
rect 17218 4128 17224 4140
rect 15988 4100 17224 4128
rect 15988 4088 15994 4100
rect 17218 4088 17224 4100
rect 17276 4088 17282 4140
rect 24210 4088 24216 4140
rect 24268 4128 24274 4140
rect 26878 4128 26884 4140
rect 24268 4100 26884 4128
rect 24268 4088 24274 4100
rect 26878 4088 26884 4100
rect 26936 4088 26942 4140
rect 213638 4088 213644 4140
rect 213696 4128 213702 4140
rect 220446 4128 220452 4140
rect 213696 4100 220452 4128
rect 213696 4088 213702 4100
rect 220446 4088 220452 4100
rect 220504 4088 220510 4140
rect 34790 4020 34796 4072
rect 34848 4060 34854 4072
rect 36538 4060 36544 4072
rect 34848 4032 36544 4060
rect 34848 4020 34854 4032
rect 36538 4020 36544 4032
rect 36596 4020 36602 4072
rect 213730 4020 213736 4072
rect 213788 4060 213794 4072
rect 220556 4060 220584 4168
rect 220832 4128 220860 4168
rect 258258 4128 258264 4140
rect 220832 4100 258264 4128
rect 258258 4088 258264 4100
rect 258316 4088 258322 4140
rect 355226 4088 355232 4140
rect 355284 4128 355290 4140
rect 365806 4128 365812 4140
rect 355284 4100 365812 4128
rect 355284 4088 355290 4100
rect 365806 4088 365812 4100
rect 365864 4088 365870 4140
rect 213788 4032 220584 4060
rect 213788 4020 213794 4032
rect 220814 4020 220820 4072
rect 220872 4060 220878 4072
rect 260650 4060 260656 4072
rect 220872 4032 260656 4060
rect 220872 4020 220878 4032
rect 260650 4020 260656 4032
rect 260708 4020 260714 4072
rect 350442 4020 350448 4072
rect 350500 4060 350506 4072
rect 362954 4060 362960 4072
rect 350500 4032 362960 4060
rect 350500 4020 350506 4032
rect 362954 4020 362960 4032
rect 363012 4020 363018 4072
rect 219342 3952 219348 4004
rect 219400 3992 219406 4004
rect 266538 3992 266544 4004
rect 219400 3964 266544 3992
rect 219400 3952 219406 3964
rect 266538 3952 266544 3964
rect 266596 3952 266602 4004
rect 349246 3952 349252 4004
rect 349304 3992 349310 4004
rect 363322 3992 363328 4004
rect 349304 3964 363328 3992
rect 349304 3952 349310 3964
rect 363322 3952 363328 3964
rect 363380 3952 363386 4004
rect 214926 3884 214932 3936
rect 214984 3924 214990 3936
rect 262950 3924 262956 3936
rect 214984 3896 262956 3924
rect 214984 3884 214990 3896
rect 262950 3884 262956 3896
rect 263008 3884 263014 3936
rect 343358 3884 343364 3936
rect 343416 3924 343422 3936
rect 364334 3924 364340 3936
rect 343416 3896 364340 3924
rect 343416 3884 343422 3896
rect 364334 3884 364340 3896
rect 364392 3884 364398 3936
rect 503070 3884 503076 3936
rect 503128 3924 503134 3936
rect 537202 3924 537208 3936
rect 503128 3896 537208 3924
rect 503128 3884 503134 3896
rect 537202 3884 537208 3896
rect 537260 3884 537266 3936
rect 217318 3816 217324 3868
rect 217376 3856 217382 3868
rect 276014 3856 276020 3868
rect 217376 3828 276020 3856
rect 217376 3816 217382 3828
rect 276014 3816 276020 3828
rect 276072 3816 276078 3868
rect 339862 3816 339868 3868
rect 339920 3856 339926 3868
rect 364610 3856 364616 3868
rect 339920 3828 364616 3856
rect 339920 3816 339926 3828
rect 364610 3816 364616 3828
rect 364668 3816 364674 3868
rect 496078 3816 496084 3868
rect 496136 3856 496142 3868
rect 533706 3856 533712 3868
rect 496136 3828 533712 3856
rect 496136 3816 496142 3828
rect 533706 3816 533712 3828
rect 533764 3816 533770 3868
rect 538858 3816 538864 3868
rect 538916 3856 538922 3868
rect 559742 3856 559748 3868
rect 538916 3828 559748 3856
rect 538916 3816 538922 3828
rect 559742 3816 559748 3828
rect 559800 3816 559806 3868
rect 219158 3748 219164 3800
rect 219216 3788 219222 3800
rect 280706 3788 280712 3800
rect 219216 3760 280712 3788
rect 219216 3748 219222 3760
rect 280706 3748 280712 3760
rect 280764 3748 280770 3800
rect 336274 3748 336280 3800
rect 336332 3788 336338 3800
rect 364518 3788 364524 3800
rect 336332 3760 364524 3788
rect 336332 3748 336338 3760
rect 364518 3748 364524 3760
rect 364576 3748 364582 3800
rect 516778 3748 516784 3800
rect 516836 3788 516842 3800
rect 516836 3760 552704 3788
rect 516836 3748 516842 3760
rect 43070 3680 43076 3732
rect 43128 3720 43134 3732
rect 50338 3720 50344 3732
rect 43128 3692 50344 3720
rect 43128 3680 43134 3692
rect 50338 3680 50344 3692
rect 50396 3680 50402 3732
rect 217410 3680 217416 3732
rect 217468 3720 217474 3732
rect 284294 3720 284300 3732
rect 217468 3692 284300 3720
rect 217468 3680 217474 3692
rect 284294 3680 284300 3692
rect 284352 3680 284358 3732
rect 332686 3680 332692 3732
rect 332744 3720 332750 3732
rect 364426 3720 364432 3732
rect 332744 3692 364432 3720
rect 332744 3680 332750 3692
rect 364426 3680 364432 3692
rect 364484 3680 364490 3732
rect 508498 3680 508504 3732
rect 508556 3720 508562 3732
rect 551462 3720 551468 3732
rect 508556 3692 551468 3720
rect 508556 3680 508562 3692
rect 551462 3680 551468 3692
rect 551520 3680 551526 3732
rect 11146 3612 11152 3664
rect 11204 3652 11210 3664
rect 35158 3652 35164 3664
rect 11204 3624 16574 3652
rect 11204 3612 11210 3624
rect 12342 3544 12348 3596
rect 12400 3584 12406 3596
rect 13078 3584 13084 3596
rect 12400 3556 13084 3584
rect 12400 3544 12406 3556
rect 13078 3544 13084 3556
rect 13136 3544 13142 3596
rect 16546 3584 16574 3624
rect 26206 3624 35164 3652
rect 26206 3584 26234 3624
rect 35158 3612 35164 3624
rect 35216 3612 35222 3664
rect 35986 3612 35992 3664
rect 36044 3652 36050 3664
rect 46198 3652 46204 3664
rect 36044 3624 46204 3652
rect 36044 3612 36050 3624
rect 46198 3612 46204 3624
rect 46256 3612 46262 3664
rect 46658 3612 46664 3664
rect 46716 3652 46722 3664
rect 46716 3624 55214 3652
rect 46716 3612 46722 3624
rect 16546 3556 26234 3584
rect 30098 3544 30104 3596
rect 30156 3584 30162 3596
rect 31018 3584 31024 3596
rect 30156 3556 31024 3584
rect 30156 3544 30162 3556
rect 31018 3544 31024 3556
rect 31076 3544 31082 3596
rect 33594 3544 33600 3596
rect 33652 3584 33658 3596
rect 35250 3584 35256 3596
rect 33652 3556 35256 3584
rect 33652 3544 33658 3556
rect 35250 3544 35256 3556
rect 35308 3544 35314 3596
rect 52454 3544 52460 3596
rect 52512 3584 52518 3596
rect 53374 3584 53380 3596
rect 52512 3556 53380 3584
rect 52512 3544 52518 3556
rect 53374 3544 53380 3556
rect 53432 3544 53438 3596
rect 55186 3584 55214 3624
rect 60826 3612 60832 3664
rect 60884 3652 60890 3664
rect 79318 3652 79324 3664
rect 60884 3624 79324 3652
rect 60884 3612 60890 3624
rect 79318 3612 79324 3624
rect 79376 3612 79382 3664
rect 96246 3612 96252 3664
rect 96304 3652 96310 3664
rect 112438 3652 112444 3664
rect 96304 3624 112444 3652
rect 96304 3612 96310 3624
rect 112438 3612 112444 3624
rect 112496 3612 112502 3664
rect 114002 3612 114008 3664
rect 114060 3652 114066 3664
rect 182818 3652 182824 3664
rect 114060 3624 182824 3652
rect 114060 3612 114066 3624
rect 182818 3612 182824 3624
rect 182876 3612 182882 3664
rect 189718 3652 189724 3664
rect 184216 3624 189724 3652
rect 116578 3584 116584 3596
rect 55186 3556 116584 3584
rect 116578 3544 116584 3556
rect 116636 3544 116642 3596
rect 118694 3544 118700 3596
rect 118752 3584 118758 3596
rect 119890 3584 119896 3596
rect 118752 3556 119896 3584
rect 118752 3544 118758 3556
rect 119890 3544 119896 3556
rect 119948 3544 119954 3596
rect 121086 3544 121092 3596
rect 121144 3584 121150 3596
rect 184216 3584 184244 3624
rect 189718 3612 189724 3624
rect 189776 3612 189782 3664
rect 213822 3612 213828 3664
rect 213880 3652 213886 3664
rect 281902 3652 281908 3664
rect 213880 3624 281908 3652
rect 213880 3612 213886 3624
rect 281902 3612 281908 3624
rect 281960 3612 281966 3664
rect 329190 3612 329196 3664
rect 329248 3652 329254 3664
rect 361758 3652 361764 3664
rect 329248 3624 361764 3652
rect 329248 3612 329254 3624
rect 361758 3612 361764 3624
rect 361816 3612 361822 3664
rect 446398 3612 446404 3664
rect 446456 3652 446462 3664
rect 523034 3652 523040 3664
rect 446456 3624 523040 3652
rect 446456 3612 446462 3624
rect 523034 3612 523040 3624
rect 523092 3612 523098 3664
rect 542998 3612 543004 3664
rect 543056 3652 543062 3664
rect 552566 3652 552572 3664
rect 543056 3624 552572 3652
rect 543056 3612 543062 3624
rect 552566 3612 552572 3624
rect 552624 3612 552630 3664
rect 121144 3556 184244 3584
rect 121144 3544 121150 3556
rect 187326 3544 187332 3596
rect 187384 3584 187390 3596
rect 188338 3584 188344 3596
rect 187384 3556 188344 3584
rect 187384 3544 187390 3556
rect 188338 3544 188344 3556
rect 188396 3544 188402 3596
rect 193214 3544 193220 3596
rect 193272 3584 193278 3596
rect 194410 3584 194416 3596
rect 193272 3556 194416 3584
rect 193272 3544 193278 3556
rect 194410 3544 194416 3556
rect 194468 3544 194474 3596
rect 195606 3544 195612 3596
rect 195664 3584 195670 3596
rect 196618 3584 196624 3596
rect 195664 3556 196624 3584
rect 195664 3544 195670 3556
rect 196618 3544 196624 3556
rect 196676 3544 196682 3596
rect 208578 3544 208584 3596
rect 208636 3584 208642 3596
rect 211798 3584 211804 3596
rect 208636 3556 211804 3584
rect 208636 3544 208642 3556
rect 211798 3544 211804 3556
rect 211856 3544 211862 3596
rect 219250 3544 219256 3596
rect 219308 3584 219314 3596
rect 287790 3584 287796 3596
rect 219308 3556 287796 3584
rect 219308 3544 219314 3556
rect 287790 3544 287796 3556
rect 287848 3544 287854 3596
rect 327994 3544 328000 3596
rect 328052 3584 328058 3596
rect 360654 3584 360660 3596
rect 328052 3556 360660 3584
rect 328052 3544 328058 3556
rect 360654 3544 360660 3556
rect 360712 3544 360718 3596
rect 385678 3544 385684 3596
rect 385736 3544 385742 3596
rect 398834 3544 398840 3596
rect 398892 3584 398898 3596
rect 400122 3584 400128 3596
rect 398892 3556 400128 3584
rect 398892 3544 398898 3556
rect 400122 3544 400128 3556
rect 400180 3544 400186 3596
rect 426158 3584 426164 3596
rect 412606 3556 426164 3584
rect 566 3476 572 3528
rect 624 3516 630 3528
rect 4798 3516 4804 3528
rect 624 3488 4804 3516
rect 624 3476 630 3488
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 5258 3476 5264 3528
rect 5316 3516 5322 3528
rect 75178 3516 75184 3528
rect 5316 3488 75184 3516
rect 5316 3476 5322 3488
rect 75178 3476 75184 3488
rect 75236 3476 75242 3528
rect 77294 3476 77300 3528
rect 77352 3516 77358 3528
rect 78214 3516 78220 3528
rect 77352 3488 78220 3516
rect 77352 3476 77358 3488
rect 78214 3476 78220 3488
rect 78272 3476 78278 3528
rect 82078 3476 82084 3528
rect 82136 3516 82142 3528
rect 104158 3516 104164 3528
rect 82136 3488 104164 3516
rect 82136 3476 82142 3488
rect 104158 3476 104164 3488
rect 104216 3476 104222 3528
rect 106918 3476 106924 3528
rect 106976 3516 106982 3528
rect 106976 3488 174952 3516
rect 106976 3476 106982 3488
rect 2774 3408 2780 3460
rect 2832 3448 2838 3460
rect 3694 3448 3700 3460
rect 2832 3420 3700 3448
rect 2832 3408 2838 3420
rect 3694 3408 3700 3420
rect 3752 3408 3758 3460
rect 20622 3408 20628 3460
rect 20680 3448 20686 3460
rect 68278 3448 68284 3460
rect 20680 3420 68284 3448
rect 20680 3408 20686 3420
rect 68278 3408 68284 3420
rect 68336 3408 68342 3460
rect 69014 3408 69020 3460
rect 69072 3448 69078 3460
rect 69934 3448 69940 3460
rect 69072 3420 69940 3448
rect 69072 3408 69078 3420
rect 69934 3408 69940 3420
rect 69992 3408 69998 3460
rect 93854 3408 93860 3460
rect 93912 3448 93918 3460
rect 94774 3448 94780 3460
rect 93912 3420 94780 3448
rect 93912 3408 93918 3420
rect 94774 3408 94780 3420
rect 94832 3408 94838 3460
rect 102134 3408 102140 3460
rect 102192 3448 102198 3460
rect 103330 3448 103336 3460
rect 102192 3420 103336 3448
rect 102192 3408 102198 3420
rect 103330 3408 103336 3420
rect 103388 3408 103394 3460
rect 174538 3448 174544 3460
rect 103486 3420 174544 3448
rect 28902 3340 28908 3392
rect 28960 3380 28966 3392
rect 32398 3380 32404 3392
rect 28960 3352 32404 3380
rect 28960 3340 28966 3352
rect 32398 3340 32404 3352
rect 32456 3340 32462 3392
rect 56042 3340 56048 3392
rect 56100 3380 56106 3392
rect 57238 3380 57244 3392
rect 56100 3352 57244 3380
rect 56100 3340 56106 3352
rect 57238 3340 57244 3352
rect 57296 3340 57302 3392
rect 59630 3340 59636 3392
rect 59688 3380 59694 3392
rect 61378 3380 61384 3392
rect 59688 3352 61384 3380
rect 59688 3340 59694 3352
rect 61378 3340 61384 3352
rect 61436 3340 61442 3392
rect 99834 3340 99840 3392
rect 99892 3380 99898 3392
rect 103486 3380 103514 3420
rect 174538 3408 174544 3420
rect 174596 3408 174602 3460
rect 174924 3448 174952 3488
rect 176654 3476 176660 3528
rect 176712 3516 176718 3528
rect 177850 3516 177856 3528
rect 176712 3488 177856 3516
rect 176712 3476 176718 3488
rect 177850 3476 177856 3488
rect 177908 3476 177914 3528
rect 190822 3476 190828 3528
rect 190880 3516 190886 3528
rect 192478 3516 192484 3528
rect 190880 3488 192484 3516
rect 190880 3476 190886 3488
rect 192478 3476 192484 3488
rect 192536 3476 192542 3528
rect 205082 3476 205088 3528
rect 205140 3516 205146 3528
rect 206278 3516 206284 3528
rect 205140 3488 206284 3516
rect 205140 3476 205146 3488
rect 206278 3476 206284 3488
rect 206336 3476 206342 3528
rect 217502 3476 217508 3528
rect 217560 3516 217566 3528
rect 291378 3516 291384 3528
rect 217560 3488 291384 3516
rect 217560 3476 217566 3488
rect 291378 3476 291384 3488
rect 291436 3476 291442 3528
rect 307938 3476 307944 3528
rect 307996 3516 308002 3528
rect 356698 3516 356704 3528
rect 307996 3488 356704 3516
rect 307996 3476 308002 3488
rect 356698 3476 356704 3488
rect 356756 3476 356762 3528
rect 365714 3476 365720 3528
rect 365772 3516 365778 3528
rect 367002 3516 367008 3528
rect 365772 3488 367008 3516
rect 365772 3476 365778 3488
rect 367002 3476 367008 3488
rect 367060 3476 367066 3528
rect 373994 3476 374000 3528
rect 374052 3516 374058 3528
rect 375282 3516 375288 3528
rect 374052 3488 375288 3516
rect 374052 3476 374058 3488
rect 375282 3476 375288 3488
rect 375340 3476 375346 3528
rect 382274 3476 382280 3528
rect 382332 3516 382338 3528
rect 383562 3516 383568 3528
rect 382332 3488 383568 3516
rect 382332 3476 382338 3488
rect 383562 3476 383568 3488
rect 383620 3476 383626 3528
rect 178678 3448 178684 3460
rect 174924 3420 178684 3448
rect 178678 3408 178684 3420
rect 178736 3408 178742 3460
rect 179046 3408 179052 3460
rect 179104 3448 179110 3460
rect 207658 3448 207664 3460
rect 179104 3420 207664 3448
rect 179104 3408 179110 3420
rect 207658 3408 207664 3420
rect 207716 3408 207722 3460
rect 214834 3408 214840 3460
rect 214892 3448 214898 3460
rect 290182 3448 290188 3460
rect 214892 3420 290188 3448
rect 214892 3408 214898 3420
rect 290182 3408 290188 3420
rect 290240 3408 290246 3460
rect 297266 3408 297272 3460
rect 297324 3448 297330 3460
rect 363598 3448 363604 3460
rect 297324 3420 363604 3448
rect 297324 3408 297330 3420
rect 363598 3408 363604 3420
rect 363656 3408 363662 3460
rect 385696 3448 385724 3544
rect 390646 3476 390652 3528
rect 390704 3516 390710 3528
rect 391842 3516 391848 3528
rect 390704 3488 391848 3516
rect 390704 3476 390710 3488
rect 391842 3476 391848 3488
rect 391900 3476 391906 3528
rect 392670 3476 392676 3528
rect 392728 3516 392734 3528
rect 412606 3516 412634 3556
rect 426158 3544 426164 3556
rect 426216 3544 426222 3596
rect 432598 3544 432604 3596
rect 432656 3584 432662 3596
rect 432656 3556 433380 3584
rect 432656 3544 432662 3556
rect 392728 3488 412634 3516
rect 392728 3476 392734 3488
rect 415486 3476 415492 3528
rect 415544 3516 415550 3528
rect 416682 3516 416688 3528
rect 415544 3488 416688 3516
rect 415544 3476 415550 3488
rect 416682 3476 416688 3488
rect 416740 3476 416746 3528
rect 423674 3476 423680 3528
rect 423732 3516 423738 3528
rect 424962 3516 424968 3528
rect 423732 3488 424968 3516
rect 423732 3476 423738 3488
rect 424962 3476 424968 3488
rect 425020 3476 425026 3528
rect 432046 3476 432052 3528
rect 432104 3516 432110 3528
rect 433242 3516 433248 3528
rect 432104 3488 433248 3516
rect 432104 3476 432110 3488
rect 433242 3476 433248 3488
rect 433300 3476 433306 3528
rect 433352 3516 433380 3556
rect 440878 3544 440884 3596
rect 440936 3584 440942 3596
rect 519538 3584 519544 3596
rect 440936 3556 519544 3584
rect 440936 3544 440942 3556
rect 519538 3544 519544 3556
rect 519596 3544 519602 3596
rect 525058 3544 525064 3596
rect 525116 3544 525122 3596
rect 531314 3544 531320 3596
rect 531372 3584 531378 3596
rect 532142 3584 532148 3596
rect 531372 3556 532148 3584
rect 531372 3544 531378 3556
rect 532142 3544 532148 3556
rect 532200 3544 532206 3596
rect 534718 3544 534724 3596
rect 534776 3584 534782 3596
rect 541986 3584 541992 3596
rect 534776 3556 541992 3584
rect 534776 3544 534782 3556
rect 541986 3544 541992 3556
rect 542044 3544 542050 3596
rect 547874 3544 547880 3596
rect 547932 3584 547938 3596
rect 548702 3584 548708 3596
rect 547932 3556 548708 3584
rect 547932 3544 547938 3556
rect 548702 3544 548708 3556
rect 548760 3544 548766 3596
rect 552676 3584 552704 3760
rect 552750 3748 552756 3800
rect 552808 3788 552814 3800
rect 552808 3760 557534 3788
rect 552808 3748 552814 3760
rect 554038 3680 554044 3732
rect 554096 3720 554102 3732
rect 557506 3720 557534 3760
rect 558178 3748 558184 3800
rect 558236 3788 558242 3800
rect 583386 3788 583392 3800
rect 558236 3760 583392 3788
rect 558236 3748 558242 3760
rect 583386 3748 583392 3760
rect 583444 3748 583450 3800
rect 577406 3720 577412 3732
rect 554096 3692 557120 3720
rect 557506 3692 577412 3720
rect 554096 3680 554102 3692
rect 554958 3584 554964 3596
rect 552676 3556 554964 3584
rect 554958 3544 554964 3556
rect 555016 3544 555022 3596
rect 556154 3544 556160 3596
rect 556212 3584 556218 3596
rect 556982 3584 556988 3596
rect 556212 3556 556988 3584
rect 556212 3544 556218 3556
rect 556982 3544 556988 3556
rect 557040 3544 557046 3596
rect 557092 3584 557120 3692
rect 577406 3680 577412 3692
rect 577464 3680 577470 3732
rect 557166 3612 557172 3664
rect 557224 3652 557230 3664
rect 573910 3652 573916 3664
rect 557224 3624 573916 3652
rect 557224 3612 557230 3624
rect 573910 3612 573916 3624
rect 573968 3612 573974 3664
rect 582190 3584 582196 3596
rect 557092 3556 582196 3584
rect 582190 3544 582196 3556
rect 582248 3544 582254 3596
rect 515950 3516 515956 3528
rect 433352 3488 515956 3516
rect 515950 3476 515956 3488
rect 516008 3476 516014 3528
rect 525076 3516 525104 3544
rect 572714 3516 572720 3528
rect 525076 3488 572720 3516
rect 572714 3476 572720 3488
rect 572772 3476 572778 3528
rect 385696 3420 415532 3448
rect 415504 3392 415532 3420
rect 417510 3408 417516 3460
rect 417568 3448 417574 3460
rect 505370 3448 505376 3460
rect 417568 3420 505376 3448
rect 417568 3408 417574 3420
rect 505370 3408 505376 3420
rect 505428 3408 505434 3460
rect 506474 3408 506480 3460
rect 506532 3448 506538 3460
rect 507302 3448 507308 3460
rect 506532 3420 507308 3448
rect 506532 3408 506538 3420
rect 507302 3408 507308 3420
rect 507360 3408 507366 3460
rect 520918 3408 520924 3460
rect 520976 3448 520982 3460
rect 569126 3448 569132 3460
rect 520976 3420 569132 3448
rect 520976 3408 520982 3420
rect 569126 3408 569132 3420
rect 569184 3408 569190 3460
rect 99892 3352 103514 3380
rect 99892 3340 99898 3352
rect 212442 3340 212448 3392
rect 212500 3380 212506 3392
rect 245194 3380 245200 3392
rect 212500 3352 245200 3380
rect 212500 3340 212506 3352
rect 245194 3340 245200 3352
rect 245252 3340 245258 3392
rect 251174 3340 251180 3392
rect 251232 3380 251238 3392
rect 252370 3380 252376 3392
rect 251232 3352 252376 3380
rect 251232 3340 251238 3352
rect 252370 3340 252376 3352
rect 252428 3340 252434 3392
rect 352834 3340 352840 3392
rect 352892 3380 352898 3392
rect 363874 3380 363880 3392
rect 352892 3352 363880 3380
rect 352892 3340 352898 3352
rect 363874 3340 363880 3352
rect 363932 3340 363938 3392
rect 415486 3340 415492 3392
rect 415544 3340 415550 3392
rect 440326 3340 440332 3392
rect 440384 3380 440390 3392
rect 441522 3380 441528 3392
rect 440384 3352 441528 3380
rect 440384 3340 440390 3352
rect 441522 3340 441528 3352
rect 441580 3340 441586 3392
rect 448606 3340 448612 3392
rect 448664 3380 448670 3392
rect 449802 3380 449808 3392
rect 448664 3352 449808 3380
rect 448664 3340 448670 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 456794 3340 456800 3392
rect 456852 3380 456858 3392
rect 458082 3380 458088 3392
rect 456852 3352 458088 3380
rect 456852 3340 456858 3352
rect 458082 3340 458088 3352
rect 458140 3340 458146 3392
rect 473354 3340 473360 3392
rect 473412 3380 473418 3392
rect 474182 3380 474188 3392
rect 473412 3352 474188 3380
rect 473412 3340 473418 3352
rect 474182 3340 474188 3352
rect 474240 3340 474246 3392
rect 481634 3340 481640 3392
rect 481692 3380 481698 3392
rect 482462 3380 482468 3392
rect 481692 3352 482468 3380
rect 481692 3340 481698 3352
rect 482462 3340 482468 3352
rect 482520 3340 482526 3392
rect 498194 3340 498200 3392
rect 498252 3380 498258 3392
rect 499022 3380 499028 3392
rect 498252 3352 499028 3380
rect 498252 3340 498258 3352
rect 499022 3340 499028 3352
rect 499080 3340 499086 3392
rect 552566 3340 552572 3392
rect 552624 3380 552630 3392
rect 557166 3380 557172 3392
rect 552624 3352 557172 3380
rect 552624 3340 552630 3352
rect 557166 3340 557172 3352
rect 557224 3340 557230 3392
rect 215202 3272 215208 3324
rect 215260 3312 215266 3324
rect 242894 3312 242900 3324
rect 215260 3284 242900 3312
rect 215260 3272 215266 3284
rect 242894 3272 242900 3284
rect 242952 3272 242958 3324
rect 354030 3272 354036 3324
rect 354088 3312 354094 3324
rect 361022 3312 361028 3324
rect 354088 3284 361028 3312
rect 354088 3272 354094 3284
rect 361022 3272 361028 3284
rect 361080 3272 361086 3324
rect 47854 3204 47860 3256
rect 47912 3244 47918 3256
rect 48958 3244 48964 3256
rect 47912 3216 48964 3244
rect 47912 3204 47918 3216
rect 48958 3204 48964 3216
rect 49016 3204 49022 3256
rect 215018 3204 215024 3256
rect 215076 3244 215082 3256
rect 240502 3244 240508 3256
rect 215076 3216 240508 3244
rect 215076 3204 215082 3216
rect 240502 3204 240508 3216
rect 240560 3204 240566 3256
rect 1670 3136 1676 3188
rect 1728 3176 1734 3188
rect 4890 3176 4896 3188
rect 1728 3148 4896 3176
rect 1728 3136 1734 3148
rect 4890 3136 4896 3148
rect 4948 3136 4954 3188
rect 38378 3136 38384 3188
rect 38436 3176 38442 3188
rect 39298 3176 39304 3188
rect 38436 3148 39304 3176
rect 38436 3136 38442 3148
rect 39298 3136 39304 3148
rect 39356 3136 39362 3188
rect 176654 3000 176660 3052
rect 176712 3040 176718 3052
rect 178770 3040 178776 3052
rect 176712 3012 178776 3040
rect 176712 3000 176718 3012
rect 178770 3000 178776 3012
rect 178828 3000 178834 3052
rect 356330 3000 356336 3052
rect 356388 3040 356394 3052
rect 362126 3040 362132 3052
rect 356388 3012 362132 3040
rect 356388 3000 356394 3012
rect 362126 3000 362132 3012
rect 362184 3000 362190 3052
rect 19426 2932 19432 2984
rect 19484 2972 19490 2984
rect 25498 2972 25504 2984
rect 19484 2944 25504 2972
rect 19484 2932 19490 2944
rect 25498 2932 25504 2944
rect 25556 2932 25562 2984
rect 41874 2864 41880 2916
rect 41932 2904 41938 2916
rect 43530 2904 43536 2916
rect 41932 2876 43536 2904
rect 41932 2864 41938 2876
rect 43530 2864 43536 2876
rect 43588 2864 43594 2916
rect 407114 2184 407120 2236
rect 407172 2224 407178 2236
rect 408402 2224 408408 2236
rect 407172 2196 408408 2224
rect 407172 2184 407178 2196
rect 408402 2184 408408 2196
rect 408460 2184 408466 2236
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 348792 700476 348844 700528
rect 358912 700476 358964 700528
rect 300124 700408 300176 700460
rect 357532 700408 357584 700460
rect 283840 700340 283892 700392
rect 358820 700340 358872 700392
rect 359464 700340 359516 700392
rect 397460 700340 397512 700392
rect 267648 700272 267700 700324
rect 357440 700272 357492 700324
rect 358084 700272 358136 700324
rect 559656 700272 559708 700324
rect 360844 699660 360896 699712
rect 364984 699660 365036 699712
rect 359556 696940 359608 696992
rect 580172 696940 580224 696992
rect 2780 683680 2832 683732
rect 4804 683680 4856 683732
rect 358176 670692 358228 670744
rect 580172 670692 580224 670744
rect 3516 656888 3568 656940
rect 178684 656888 178736 656940
rect 2780 632068 2832 632120
rect 4896 632068 4948 632120
rect 362224 630640 362276 630692
rect 580172 630640 580224 630692
rect 359648 616836 359700 616888
rect 580172 616836 580224 616888
rect 3332 605820 3384 605872
rect 203524 605820 203576 605872
rect 362316 590656 362368 590708
rect 579620 590656 579672 590708
rect 2780 579912 2832 579964
rect 4988 579912 5040 579964
rect 3056 565836 3108 565888
rect 31024 565836 31076 565888
rect 217968 565088 218020 565140
rect 234620 565088 234672 565140
rect 331220 565088 331272 565140
rect 359004 565088 359056 565140
rect 371884 563048 371936 563100
rect 580172 563048 580224 563100
rect 2780 553664 2832 553716
rect 5080 553664 5132 553716
rect 358268 536800 358320 536852
rect 580172 536800 580224 536852
rect 3332 527756 3384 527808
rect 8944 527756 8996 527808
rect 358360 484372 358412 484424
rect 580172 484372 580224 484424
rect 217416 478864 217468 478916
rect 220084 478864 220136 478916
rect 311900 478184 311952 478236
rect 358912 478184 358964 478236
rect 3700 478116 3752 478168
rect 354680 478116 354732 478168
rect 280252 476688 280304 476740
rect 302240 476688 302292 476740
rect 241612 476620 241664 476672
rect 252560 476620 252612 476672
rect 255412 476620 255464 476672
rect 264980 476620 265032 476672
rect 281540 476620 281592 476672
rect 305000 476620 305052 476672
rect 259552 476552 259604 476604
rect 270500 476552 270552 476604
rect 283104 476552 283156 476604
rect 307760 476552 307812 476604
rect 238760 476484 238812 476536
rect 244280 476484 244332 476536
rect 236092 476416 236144 476468
rect 247040 476416 247092 476468
rect 238852 476348 238904 476400
rect 249800 476484 249852 476536
rect 252652 476484 252704 476536
rect 263600 476484 263652 476536
rect 265072 476484 265124 476536
rect 280160 476484 280212 476536
rect 284300 476484 284352 476536
rect 310520 476484 310572 476536
rect 251180 476416 251232 476468
rect 260840 476416 260892 476468
rect 258172 476348 258224 476400
rect 268016 476416 268068 476468
rect 285680 476416 285732 476468
rect 313280 476416 313332 476468
rect 234712 476280 234764 476332
rect 242900 476280 242952 476332
rect 245752 476280 245804 476332
rect 255320 476280 255372 476332
rect 241520 476212 241572 476264
rect 244280 476212 244332 476264
rect 248420 476212 248472 476264
rect 242808 476144 242860 476196
rect 244924 476144 244976 476196
rect 252376 476144 252428 476196
rect 256700 476144 256752 476196
rect 260932 476280 260984 476332
rect 273260 476348 273312 476400
rect 287244 476348 287296 476400
rect 314660 476348 314712 476400
rect 263692 476280 263744 476332
rect 277860 476280 277912 476332
rect 288532 476280 288584 476332
rect 317420 476280 317472 476332
rect 262404 476212 262456 476264
rect 276020 476212 276072 476264
rect 292764 476212 292816 476264
rect 322940 476212 322992 476264
rect 258264 476144 258316 476196
rect 267740 476144 267792 476196
rect 282920 476144 282972 476196
rect 290004 476144 290056 476196
rect 320180 476144 320232 476196
rect 234620 476076 234672 476128
rect 235908 476076 235960 476128
rect 241428 476076 241480 476128
rect 242900 476076 242952 476128
rect 244280 476076 244332 476128
rect 245660 476076 245712 476128
rect 251088 476076 251140 476128
rect 252560 476076 252612 476128
rect 263508 476076 263560 476128
rect 267004 476076 267056 476128
rect 280068 476076 280120 476128
rect 282184 476076 282236 476128
rect 293960 476076 294012 476128
rect 325792 476076 325844 476128
rect 219072 475396 219124 475448
rect 249892 475396 249944 475448
rect 217600 475328 217652 475380
rect 253940 475328 253992 475380
rect 3332 474716 3384 474768
rect 333980 474716 334032 474768
rect 217508 473968 217560 474020
rect 251272 473968 251324 474020
rect 219164 472608 219216 472660
rect 247132 472608 247184 472660
rect 3424 462340 3476 462392
rect 335360 462340 335412 462392
rect 271972 461660 272024 461712
rect 289912 461660 289964 461712
rect 273260 461592 273312 461644
rect 292672 461592 292724 461644
rect 274548 460300 274600 460352
rect 285128 460300 285180 460352
rect 273168 460232 273220 460284
rect 283012 460232 283064 460284
rect 270592 460164 270644 460216
rect 287152 460164 287204 460216
rect 266268 458940 266320 458992
rect 274640 458940 274692 458992
rect 267556 458872 267608 458924
rect 276020 458872 276072 458924
rect 271788 458804 271840 458856
rect 282092 458804 282144 458856
rect 269028 457716 269080 457768
rect 279056 457716 279108 457768
rect 270408 457648 270460 457700
rect 280528 457648 280580 457700
rect 275192 457580 275244 457632
rect 295340 457580 295392 457632
rect 276572 457512 276624 457564
rect 298100 457512 298152 457564
rect 217876 457444 217928 457496
rect 256792 457444 256844 457496
rect 267648 457444 267700 457496
rect 277400 457444 277452 457496
rect 277952 457444 278004 457496
rect 300860 457444 300912 457496
rect 300860 456220 300912 456272
rect 362224 456220 362276 456272
rect 219256 456152 219308 456204
rect 240968 456152 241020 456204
rect 278688 456152 278740 456204
rect 291384 456152 291436 456204
rect 303160 456152 303212 456204
rect 580264 456152 580316 456204
rect 219348 456084 219400 456136
rect 244372 456084 244424 456136
rect 269212 456084 269264 456136
rect 285772 456084 285824 456136
rect 298376 456084 298428 456136
rect 580448 456084 580500 456136
rect 3608 456016 3660 456068
rect 333520 456016 333572 456068
rect 218060 454928 218112 454980
rect 317420 454928 317472 454980
rect 31024 454860 31076 454912
rect 331220 454860 331272 454912
rect 337384 454860 337436 454912
rect 359464 454860 359516 454912
rect 3332 454792 3384 454844
rect 325700 454792 325752 454844
rect 325792 454792 325844 454844
rect 362316 454792 362368 454844
rect 3516 454724 3568 454776
rect 328736 454724 328788 454776
rect 329840 454724 329892 454776
rect 359556 454724 359608 454776
rect 5080 454656 5132 454708
rect 354772 454656 354824 454708
rect 323400 453636 323452 453688
rect 358268 453636 358320 453688
rect 321008 453568 321060 453620
rect 358360 453568 358412 453620
rect 310888 453500 310940 453552
rect 360844 453500 360896 453552
rect 203524 453432 203576 453484
rect 353760 453432 353812 453484
rect 178684 453364 178736 453416
rect 353392 453364 353444 453416
rect 6920 453296 6972 453348
rect 351368 453296 351420 453348
rect 303896 452208 303948 452260
rect 358084 452208 358136 452260
rect 308496 452140 308548 452192
rect 429200 452140 429252 452192
rect 306380 452072 306432 452124
rect 494060 452072 494112 452124
rect 71780 452004 71832 452056
rect 349252 452004 349304 452056
rect 8944 451936 8996 451988
rect 331864 451936 331916 451988
rect 4988 451868 5040 451920
rect 329932 451868 329984 451920
rect 301964 450780 302016 450832
rect 358176 450780 358228 450832
rect 299664 450712 299716 450764
rect 359648 450712 359700 450764
rect 217692 450644 217744 450696
rect 234252 450644 234304 450696
rect 297272 450644 297324 450696
rect 371884 450644 371936 450696
rect 4804 450576 4856 450628
rect 325332 450576 325384 450628
rect 4896 450508 4948 450560
rect 327632 450508 327684 450560
rect 335452 450508 335504 450560
rect 462320 450508 462372 450560
rect 310520 449488 310572 449540
rect 412640 449488 412692 449540
rect 153200 449420 153252 449472
rect 319904 449420 319956 449472
rect 308220 449352 308272 449404
rect 477500 449352 477552 449404
rect 88340 449284 88392 449336
rect 322204 449284 322256 449336
rect 305828 449216 305880 449268
rect 542360 449216 542412 449268
rect 23480 449148 23532 449200
rect 324504 449148 324556 449200
rect 201500 448128 201552 448180
rect 344744 448128 344796 448180
rect 169760 448060 169812 448112
rect 318340 448060 318392 448112
rect 136640 447992 136692 448044
rect 347044 447992 347096 448044
rect 104900 447924 104952 447976
rect 320640 447924 320692 447976
rect 333060 447924 333112 447976
rect 527180 447924 527232 447976
rect 40040 447856 40092 447908
rect 322940 447856 322992 447908
rect 328460 447856 328512 447908
rect 580356 447856 580408 447908
rect 2872 447788 2924 447840
rect 356428 447788 356480 447840
rect 244280 447244 244332 447296
rect 244924 447244 244976 447296
rect 249800 447244 249852 447296
rect 250260 447244 250312 447296
rect 283012 447244 283064 447296
rect 283748 447244 283800 447296
rect 325700 447244 325752 447296
rect 326620 447244 326672 447296
rect 329840 447244 329892 447296
rect 330484 447244 330536 447296
rect 354680 447244 354732 447296
rect 355324 447244 355376 447296
rect 245016 447040 245068 447092
rect 246764 447040 246816 447092
rect 252468 447040 252520 447092
rect 255320 447040 255372 447092
rect 262864 447040 262916 447092
rect 270040 447040 270092 447092
rect 253848 446972 253900 447024
rect 259184 446972 259236 447024
rect 259368 446972 259420 447024
rect 265440 446972 265492 447024
rect 255228 446904 255280 446956
rect 260380 446904 260432 446956
rect 261484 446904 261536 446956
rect 268476 446972 268528 447024
rect 217968 446836 218020 446888
rect 315948 446836 316000 446888
rect 210424 446768 210476 446820
rect 345940 446768 345992 446820
rect 267004 446632 267056 446684
rect 271604 446632 271656 446684
rect 282184 446632 282236 446684
rect 293408 446632 293460 446684
rect 340052 446632 340104 446684
rect 359004 446632 359056 446684
rect 256608 446564 256660 446616
rect 262312 446564 262364 446616
rect 276664 446564 276716 446616
rect 288716 446564 288768 446616
rect 307392 446564 307444 446616
rect 340880 446564 340932 446616
rect 342444 446564 342496 446616
rect 357440 446564 357492 446616
rect 220084 446496 220136 446548
rect 232780 446496 232832 446548
rect 260748 446496 260800 446548
rect 267004 446496 267056 446548
rect 275284 446496 275336 446548
rect 287152 446496 287204 446548
rect 315212 446496 315264 446548
rect 358820 446496 358872 446548
rect 217784 446428 217836 446480
rect 233516 446428 233568 446480
rect 257988 446428 258040 446480
rect 263876 446428 263928 446480
rect 264888 446428 264940 446480
rect 273168 446428 273220 446480
rect 278044 446428 278096 446480
rect 290280 446428 290332 446480
rect 313648 446428 313700 446480
rect 357532 446428 357584 446480
rect 256700 446360 256752 446412
rect 257252 446360 257304 446412
rect 309784 446360 309836 446412
rect 346308 446360 346360 446412
rect 318708 446292 318760 446344
rect 357992 446292 358044 446344
rect 314384 446224 314436 446276
rect 364984 446224 365036 446276
rect 288348 446156 288400 446208
rect 359556 446156 359608 446208
rect 232320 446088 232372 446140
rect 338488 446088 338540 446140
rect 233792 446020 233844 446072
rect 343180 446020 343232 446072
rect 343272 446020 343324 446072
rect 357164 446020 357216 446072
rect 231124 445952 231176 446004
rect 347872 445952 347924 446004
rect 232228 445884 232280 445936
rect 352564 445884 352616 445936
rect 233884 445816 233936 445868
rect 360292 445816 360344 445868
rect 305092 445748 305144 445800
rect 338764 445748 338816 445800
rect 351920 445748 351972 445800
rect 358728 445748 358780 445800
rect 4896 445136 4948 445188
rect 345572 445136 345624 445188
rect 346308 445136 346360 445188
rect 580632 445136 580684 445188
rect 40684 445068 40736 445120
rect 337016 445068 337068 445120
rect 340880 445068 340932 445120
rect 580540 445068 580592 445120
rect 3884 445000 3936 445052
rect 318708 445000 318760 445052
rect 338764 445000 338816 445052
rect 580448 445000 580500 445052
rect 312084 444932 312136 444984
rect 367744 444932 367796 444984
rect 231216 444864 231268 444916
rect 340880 444864 340932 444916
rect 228364 444796 228416 444848
rect 344008 444796 344060 444848
rect 218428 444728 218480 444780
rect 348608 444728 348660 444780
rect 174544 444660 174596 444712
rect 341616 444660 341668 444712
rect 106924 444592 106976 444644
rect 339316 444592 339368 444644
rect 316776 444524 316828 444576
rect 365076 444524 365128 444576
rect 43444 444456 43496 444508
rect 350172 444456 350224 444508
rect 319076 444388 319128 444440
rect 365168 444388 365220 444440
rect 3792 443912 3844 443964
rect 233792 443912 233844 443964
rect 3516 443844 3568 443896
rect 233884 443844 233936 443896
rect 3608 443776 3660 443828
rect 288348 444048 288400 444100
rect 3976 443708 4028 443760
rect 343272 443708 343324 443760
rect 3700 443640 3752 443692
rect 351920 443640 351972 443692
rect 320824 443572 320876 443624
rect 298192 443436 298244 443488
rect 180064 443096 180116 443148
rect 303160 443436 303212 443488
rect 320824 443436 320876 443488
rect 360844 443436 360896 443488
rect 580356 443028 580408 443080
rect 580264 442960 580316 443012
rect 3424 433984 3476 434036
rect 232228 433984 232280 434036
rect 365168 431876 365220 431928
rect 580172 431876 580224 431928
rect 3332 423580 3384 423632
rect 40684 423580 40736 423632
rect 3332 411204 3384 411256
rect 232228 411204 232280 411256
rect 365076 379448 365128 379500
rect 579620 379448 579672 379500
rect 3332 372512 3384 372564
rect 106924 372512 106976 372564
rect 3332 358708 3384 358760
rect 231216 358708 231268 358760
rect 364984 325592 365036 325644
rect 579988 325592 580040 325644
rect 3332 320084 3384 320136
rect 174544 320084 174596 320136
rect 305000 310496 305052 310548
rect 305184 310496 305236 310548
rect 309416 310496 309468 310548
rect 309784 310496 309836 310548
rect 310796 310496 310848 310548
rect 311164 310496 311216 310548
rect 312176 310496 312228 310548
rect 312544 310496 312596 310548
rect 215208 309068 215260 309120
rect 279700 309068 279752 309120
rect 323768 309068 323820 309120
rect 359004 309068 359056 309120
rect 216496 309000 216548 309052
rect 280436 309000 280488 309052
rect 324504 309000 324556 309052
rect 361488 309000 361540 309052
rect 189724 308932 189776 308984
rect 255964 308932 256016 308984
rect 316408 308932 316460 308984
rect 326344 308932 326396 308984
rect 331128 308932 331180 308984
rect 331496 308932 331548 308984
rect 354220 308932 354272 308984
rect 367284 308932 367336 308984
rect 182824 308864 182876 308916
rect 254584 308864 254636 308916
rect 294972 308864 295024 308916
rect 356888 308864 356940 308916
rect 356980 308864 357032 308916
rect 369124 308864 369176 308916
rect 213828 308796 213880 308848
rect 287336 308796 287388 308848
rect 294236 308796 294288 308848
rect 356152 308796 356204 308848
rect 178684 308728 178736 308780
rect 253204 308728 253256 308780
rect 294512 308728 294564 308780
rect 357072 308728 357124 308780
rect 68284 308660 68336 308712
rect 236368 308660 236420 308712
rect 50344 308592 50396 308644
rect 240784 308592 240836 308644
rect 253388 308592 253440 308644
rect 266636 308660 266688 308712
rect 291292 308660 291344 308712
rect 355324 308660 355376 308712
rect 356520 308660 356572 308712
rect 292672 308592 292724 308644
rect 357256 308592 357308 308644
rect 46204 308524 46256 308576
rect 239404 308524 239456 308576
rect 248604 308524 248656 308576
rect 249156 308524 249208 308576
rect 290556 308524 290608 308576
rect 355416 308524 355468 308576
rect 358360 308524 358412 308576
rect 368848 308524 368900 308576
rect 370136 308524 370188 308576
rect 32404 308456 32456 308508
rect 233056 308456 233108 308508
rect 233332 308456 233384 308508
rect 234160 308456 234212 308508
rect 247224 308456 247276 308508
rect 247960 308456 248012 308508
rect 248420 308456 248472 308508
rect 248788 308456 248840 308508
rect 252744 308456 252796 308508
rect 253020 308456 253072 308508
rect 271880 308456 271932 308508
rect 272156 308456 272208 308508
rect 290832 308456 290884 308508
rect 357164 308456 357216 308508
rect 25504 308388 25556 308440
rect 231768 308388 231820 308440
rect 231952 308388 232004 308440
rect 232780 308388 232832 308440
rect 233240 308388 233292 308440
rect 233700 308388 233752 308440
rect 247132 308388 247184 308440
rect 247868 308388 247920 308440
rect 248696 308388 248748 308440
rect 249524 308388 249576 308440
rect 249892 308388 249944 308440
rect 250536 308388 250588 308440
rect 251548 308388 251600 308440
rect 252284 308388 252336 308440
rect 252652 308388 252704 308440
rect 253296 308388 253348 308440
rect 264980 308388 265032 308440
rect 265348 308388 265400 308440
rect 266452 308388 266504 308440
rect 266820 308388 266872 308440
rect 269212 308388 269264 308440
rect 270040 308388 270092 308440
rect 270684 308388 270736 308440
rect 271512 308388 271564 308440
rect 271972 308388 272024 308440
rect 272800 308388 272852 308440
rect 218980 308320 219032 308372
rect 279056 308320 279108 308372
rect 219072 308252 219124 308304
rect 277676 308252 277728 308304
rect 218888 308184 218940 308236
rect 244372 308116 244424 308168
rect 244740 308116 244792 308168
rect 245936 308116 245988 308168
rect 246580 308116 246632 308168
rect 249984 308116 250036 308168
rect 250260 308116 250312 308168
rect 252836 308116 252888 308168
rect 253664 308116 253716 308168
rect 231768 308048 231820 308100
rect 236184 308048 236236 308100
rect 244556 308048 244608 308100
rect 245200 308048 245252 308100
rect 246028 308048 246080 308100
rect 246948 308048 247000 308100
rect 263508 308184 263560 308236
rect 264060 308184 264112 308236
rect 266544 308184 266596 308236
rect 267372 308184 267424 308236
rect 268016 308184 268068 308236
rect 268752 308184 268804 308236
rect 269304 308184 269356 308236
rect 270132 308184 270184 308236
rect 270500 308184 270552 308236
rect 270960 308184 271012 308236
rect 289912 308184 289964 308236
rect 357808 308388 357860 308440
rect 358820 308388 358872 308440
rect 370504 308388 370556 308440
rect 356152 308320 356204 308372
rect 356980 308320 357032 308372
rect 358268 308320 358320 308372
rect 360016 308320 360068 308372
rect 355600 308252 355652 308304
rect 367928 308252 367980 308304
rect 355140 308184 355192 308236
rect 367560 308184 367612 308236
rect 263692 308116 263744 308168
rect 264336 308116 264388 308168
rect 265256 308116 265308 308168
rect 265992 308116 266044 308168
rect 276296 308116 276348 308168
rect 359648 308116 359700 308168
rect 362316 308116 362368 308168
rect 270500 308048 270552 308100
rect 271420 308048 271472 308100
rect 326344 308048 326396 308100
rect 331772 308048 331824 308100
rect 351000 308048 351052 308100
rect 359464 308048 359516 308100
rect 360200 308048 360252 308100
rect 368756 308048 368808 308100
rect 233056 307980 233108 308032
rect 238024 307980 238076 308032
rect 244372 307980 244424 308032
rect 245108 307980 245160 308032
rect 249984 307980 250036 308032
rect 250904 307980 250956 308032
rect 263784 307980 263836 308032
rect 264704 307980 264756 308032
rect 267740 307980 267792 308032
rect 268108 307980 268160 308032
rect 356060 307980 356112 308032
rect 366456 307980 366508 308032
rect 256792 307912 256844 307964
rect 257344 307912 257396 307964
rect 354680 307912 354732 307964
rect 253204 307844 253256 307896
rect 259000 307844 259052 307896
rect 360108 307912 360160 307964
rect 362776 307912 362828 307964
rect 257344 307776 257396 307828
rect 258264 307776 258316 307828
rect 260288 307776 260340 307828
rect 262404 307776 262456 307828
rect 358176 307776 358228 307828
rect 359556 307776 359608 307828
rect 360936 307844 360988 307896
rect 363696 307844 363748 307896
rect 361028 307776 361080 307828
rect 361580 307776 361632 307828
rect 367376 307776 367428 307828
rect 251364 307640 251416 307692
rect 251916 307640 251968 307692
rect 267740 307640 267792 307692
rect 268660 307640 268712 307692
rect 359832 307640 359884 307692
rect 361396 307640 361448 307692
rect 266636 307504 266688 307556
rect 266912 307504 266964 307556
rect 264980 307232 265032 307284
rect 265900 307232 265952 307284
rect 202880 307164 202932 307216
rect 271880 307164 271932 307216
rect 314844 307164 314896 307216
rect 422300 307164 422352 307216
rect 189080 307096 189132 307148
rect 269488 307096 269540 307148
rect 269580 307096 269632 307148
rect 272064 307096 272116 307148
rect 272248 307096 272300 307148
rect 321928 307096 321980 307148
rect 458180 307096 458232 307148
rect 67640 307028 67692 307080
rect 245568 307028 245620 307080
rect 245752 306960 245804 307012
rect 246488 306960 246540 307012
rect 254308 306960 254360 307012
rect 254492 306960 254544 307012
rect 261024 306960 261076 307012
rect 272064 306960 272116 307012
rect 272892 306960 272944 307012
rect 300860 306960 300912 307012
rect 301136 306960 301188 307012
rect 317788 306960 317840 307012
rect 326068 306960 326120 307012
rect 480260 307028 480312 307080
rect 336832 306960 336884 307012
rect 337016 306960 337068 307012
rect 269580 306892 269632 306944
rect 261024 306756 261076 306808
rect 317788 306756 317840 306808
rect 243268 306688 243320 306740
rect 299572 306552 299624 306604
rect 300216 306552 300268 306604
rect 328644 306552 328696 306604
rect 329012 306552 329064 306604
rect 332692 306552 332744 306604
rect 332876 306552 332928 306604
rect 236092 306484 236144 306536
rect 237288 306484 237340 306536
rect 243268 306484 243320 306536
rect 234804 306416 234856 306468
rect 235908 306416 235960 306468
rect 236184 306416 236236 306468
rect 236828 306416 236880 306468
rect 237564 306416 237616 306468
rect 237840 306416 237892 306468
rect 240232 306416 240284 306468
rect 241060 306416 241112 306468
rect 243084 306416 243136 306468
rect 244188 306416 244240 306468
rect 254032 306416 254084 306468
rect 254676 306416 254728 306468
rect 255412 306416 255464 306468
rect 256056 306416 256108 306468
rect 256976 306416 257028 306468
rect 257436 306416 257488 306468
rect 259460 306416 259512 306468
rect 259828 306416 259880 306468
rect 260840 306416 260892 306468
rect 261208 306416 261260 306468
rect 234712 306348 234764 306400
rect 235540 306348 235592 306400
rect 236276 306348 236328 306400
rect 236920 306348 236972 306400
rect 237472 306348 237524 306400
rect 238208 306348 238260 306400
rect 238852 306348 238904 306400
rect 239588 306348 239640 306400
rect 240416 306348 240468 306400
rect 240968 306348 241020 306400
rect 241612 306348 241664 306400
rect 242348 306348 242400 306400
rect 242992 306348 243044 306400
rect 243728 306348 243780 306400
rect 254216 306348 254268 306400
rect 255044 306348 255096 306400
rect 255504 306348 255556 306400
rect 255780 306348 255832 306400
rect 257160 306348 257212 306400
rect 257804 306348 257856 306400
rect 261116 306348 261168 306400
rect 261576 306348 261628 306400
rect 262404 306348 262456 306400
rect 263324 306348 263376 306400
rect 216404 306280 216456 306332
rect 279976 306484 280028 306536
rect 288532 306484 288584 306536
rect 273076 306416 273128 306468
rect 273352 306348 273404 306400
rect 273812 306348 273864 306400
rect 273536 306280 273588 306332
rect 274180 306280 274232 306332
rect 280988 306416 281040 306468
rect 285956 306416 286008 306468
rect 288808 306416 288860 306468
rect 284300 306348 284352 306400
rect 285496 306348 285548 306400
rect 281816 306280 281868 306332
rect 284668 306280 284720 306332
rect 285128 306280 285180 306332
rect 286048 306280 286100 306332
rect 286876 306280 286928 306332
rect 218704 306212 218756 306264
rect 273076 306212 273128 306264
rect 284392 306212 284444 306264
rect 284576 306212 284628 306264
rect 285772 306212 285824 306264
rect 286140 306212 286192 306264
rect 288624 306212 288676 306264
rect 296812 306484 296864 306536
rect 297180 306484 297232 306536
rect 292948 306416 293000 306468
rect 327080 306416 327132 306468
rect 327448 306416 327500 306468
rect 289820 306348 289872 306400
rect 291016 306348 291068 306400
rect 292672 306348 292724 306400
rect 298100 306348 298152 306400
rect 298652 306348 298704 306400
rect 302424 306348 302476 306400
rect 302884 306348 302936 306400
rect 305092 306348 305144 306400
rect 306012 306348 306064 306400
rect 307852 306348 307904 306400
rect 308772 306348 308824 306400
rect 316132 306348 316184 306400
rect 316960 306348 317012 306400
rect 321652 306348 321704 306400
rect 322480 306348 322532 306400
rect 324320 306348 324372 306400
rect 325240 306348 325292 306400
rect 328460 306348 328512 306400
rect 329288 306348 329340 306400
rect 329932 306348 329984 306400
rect 330208 306348 330260 306400
rect 331588 306348 331640 306400
rect 331956 306348 332008 306400
rect 289912 306280 289964 306332
rect 290188 306280 290240 306332
rect 291292 306280 291344 306332
rect 291936 306280 291988 306332
rect 293960 306280 294012 306332
rect 295156 306280 295208 306332
rect 298284 306280 298336 306332
rect 298744 306280 298796 306332
rect 299572 306280 299624 306332
rect 300492 306280 300544 306332
rect 300952 306280 301004 306332
rect 301964 306280 302016 306332
rect 302608 306280 302660 306332
rect 303252 306280 303304 306332
rect 305184 306280 305236 306332
rect 306104 306280 306156 306332
rect 306380 306280 306432 306332
rect 307484 306280 307536 306332
rect 307760 306280 307812 306332
rect 308312 306280 308364 306332
rect 309232 306280 309284 306332
rect 310152 306280 310204 306332
rect 310520 306280 310572 306332
rect 311532 306280 311584 306332
rect 311992 306280 312044 306332
rect 312912 306280 312964 306332
rect 314752 306280 314804 306332
rect 315580 306280 315632 306332
rect 316040 306280 316092 306332
rect 316868 306280 316920 306332
rect 317696 306280 317748 306332
rect 318248 306280 318300 306332
rect 318800 306280 318852 306332
rect 320088 306280 320140 306332
rect 320180 306280 320232 306332
rect 321468 306280 321520 306332
rect 321560 306280 321612 306332
rect 322388 306280 322440 306332
rect 323032 306280 323084 306332
rect 323400 306280 323452 306332
rect 324412 306280 324464 306332
rect 325148 306280 325200 306332
rect 325792 306280 325844 306332
rect 326620 306280 326672 306332
rect 327172 306280 327224 306332
rect 328000 306280 328052 306332
rect 328644 306280 328696 306332
rect 329380 306280 329432 306332
rect 329840 306280 329892 306332
rect 330300 306280 330352 306332
rect 331496 306280 331548 306332
rect 331864 306280 331916 306332
rect 335636 306280 335688 306332
rect 336004 306280 336056 306332
rect 337108 306280 337160 306332
rect 337476 306280 337528 306332
rect 341156 306280 341208 306332
rect 341524 306280 341576 306332
rect 342720 306484 342772 306536
rect 342628 306416 342680 306468
rect 343640 306416 343692 306468
rect 344008 306416 344060 306468
rect 357716 306416 357768 306468
rect 357992 306416 358044 306468
rect 358360 306416 358412 306468
rect 360016 306416 360068 306468
rect 360292 306416 360344 306468
rect 360752 306416 360804 306468
rect 288900 306212 288952 306264
rect 291476 306212 291528 306264
rect 292396 306212 292448 306264
rect 292856 306212 292908 306264
rect 293776 306212 293828 306264
rect 296904 306212 296956 306264
rect 297548 306212 297600 306264
rect 298192 306212 298244 306264
rect 299204 306212 299256 306264
rect 302332 306212 302384 306264
rect 303344 306212 303396 306264
rect 303620 306212 303672 306264
rect 304080 306212 304132 306264
rect 321744 306212 321796 306264
rect 322020 306212 322072 306264
rect 323124 306212 323176 306264
rect 323860 306212 323912 306264
rect 325976 306212 326028 306264
rect 326988 306212 327040 306264
rect 327264 306212 327316 306264
rect 327540 306212 327592 306264
rect 328828 306212 328880 306264
rect 329748 306212 329800 306264
rect 331312 306212 331364 306264
rect 332324 306212 332376 306264
rect 332600 306212 332652 306264
rect 332968 306212 333020 306264
rect 340972 306212 341024 306264
rect 341340 306212 341392 306264
rect 342260 306212 342312 306264
rect 214564 306144 214616 306196
rect 277860 306144 277912 306196
rect 285864 306144 285916 306196
rect 286508 306144 286560 306196
rect 288716 306144 288768 306196
rect 289636 306144 289688 306196
rect 294052 306144 294104 306196
rect 294696 306144 294748 306196
rect 296812 306144 296864 306196
rect 297916 306144 297968 306196
rect 303988 306144 304040 306196
rect 304724 306144 304776 306196
rect 319168 306144 319220 306196
rect 319628 306144 319680 306196
rect 320548 306144 320600 306196
rect 321100 306144 321152 306196
rect 321836 306144 321888 306196
rect 322848 306144 322900 306196
rect 327356 306144 327408 306196
rect 328368 306144 328420 306196
rect 333980 306144 334032 306196
rect 334440 306144 334492 306196
rect 335360 306144 335412 306196
rect 335820 306144 335872 306196
rect 337016 306144 337068 306196
rect 337844 306144 337896 306196
rect 338212 306144 338264 306196
rect 338580 306144 338632 306196
rect 339500 306144 339552 306196
rect 339960 306144 340012 306196
rect 340880 306144 340932 306196
rect 341984 306144 342036 306196
rect 216312 306076 216364 306128
rect 281080 306076 281132 306128
rect 284392 306076 284444 306128
rect 285036 306076 285088 306128
rect 288532 306076 288584 306128
rect 289176 306076 289228 306128
rect 295340 306076 295392 306128
rect 295708 306076 295760 306128
rect 299848 306076 299900 306128
rect 300584 306076 300636 306128
rect 303804 306076 303856 306128
rect 304632 306076 304684 306128
rect 313464 306076 313516 306128
rect 314292 306076 314344 306128
rect 319076 306076 319128 306128
rect 319720 306076 319772 306128
rect 330024 306076 330076 306128
rect 330760 306076 330812 306128
rect 332600 306076 332652 306128
rect 333336 306076 333388 306128
rect 334164 306076 334216 306128
rect 335084 306076 335136 306128
rect 336740 306076 336792 306128
rect 337384 306076 337436 306128
rect 338396 306076 338448 306128
rect 339224 306076 339276 306128
rect 339592 306076 339644 306128
rect 340604 306076 340656 306128
rect 355876 306280 355928 306332
rect 360200 306348 360252 306400
rect 360476 306348 360528 306400
rect 361120 306348 361172 306400
rect 363052 306348 363104 306400
rect 363236 306348 363288 306400
rect 343732 306212 343784 306264
rect 344744 306212 344796 306264
rect 345020 306212 345072 306264
rect 345480 306212 345532 306264
rect 357624 306212 357676 306264
rect 358084 306212 358136 306264
rect 354956 306144 355008 306196
rect 371424 306280 371476 306332
rect 342812 306076 342864 306128
rect 357808 306076 357860 306128
rect 358084 306076 358136 306128
rect 359924 306212 359976 306264
rect 360200 306212 360252 306264
rect 371332 306212 371384 306264
rect 215024 306008 215076 306060
rect 279240 306008 279292 306060
rect 288808 306008 288860 306060
rect 289268 306008 289320 306060
rect 295616 306008 295668 306060
rect 296536 306008 296588 306060
rect 303620 306008 303672 306060
rect 304264 306008 304316 306060
rect 332784 306008 332836 306060
rect 333704 306008 333756 306060
rect 333980 306008 334032 306060
rect 334716 306008 334768 306060
rect 338212 306008 338264 306060
rect 338856 306008 338908 306060
rect 342352 306008 342404 306060
rect 343364 306008 343416 306060
rect 355508 306008 355560 306060
rect 214656 305940 214708 305992
rect 280620 305940 280672 305992
rect 295340 305940 295392 305992
rect 296168 305940 296220 305992
rect 354036 305940 354088 305992
rect 358360 305940 358412 305992
rect 369216 306144 369268 306196
rect 359924 306076 359976 306128
rect 371884 306076 371936 306128
rect 360016 306008 360068 306060
rect 371516 306008 371568 306060
rect 213736 305872 213788 305924
rect 282736 305872 282788 305924
rect 352840 305872 352892 305924
rect 358820 305940 358872 305992
rect 369032 305940 369084 305992
rect 358544 305872 358596 305924
rect 370412 305872 370464 305924
rect 214472 305804 214524 305856
rect 283472 305804 283524 305856
rect 354496 305804 354548 305856
rect 371792 305804 371844 305856
rect 216128 305736 216180 305788
rect 288072 305736 288124 305788
rect 350080 305736 350132 305788
rect 368940 305736 368992 305788
rect 214748 305668 214800 305720
rect 287612 305668 287664 305720
rect 352196 305668 352248 305720
rect 358544 305668 358596 305720
rect 358728 305668 358780 305720
rect 370320 305668 370372 305720
rect 217692 305600 217744 305652
rect 345664 305600 345716 305652
rect 346584 305600 346636 305652
rect 369308 305600 369360 305652
rect 215116 305532 215168 305584
rect 276480 305532 276532 305584
rect 348240 305532 348292 305584
rect 363788 305532 363840 305584
rect 216588 305464 216640 305516
rect 278596 305464 278648 305516
rect 357348 305464 357400 305516
rect 371700 305464 371752 305516
rect 216220 305396 216272 305448
rect 277216 305396 277268 305448
rect 351460 305396 351512 305448
rect 358820 305396 358872 305448
rect 359096 305396 359148 305448
rect 359740 305396 359792 305448
rect 234988 305328 235040 305380
rect 235448 305328 235500 305380
rect 237656 305328 237708 305380
rect 238300 305328 238352 305380
rect 239128 305328 239180 305380
rect 240048 305328 240100 305380
rect 241796 305328 241848 305380
rect 242440 305328 242492 305380
rect 253940 305328 253992 305380
rect 254308 305328 254360 305380
rect 255504 305328 255556 305380
rect 256424 305328 256476 305380
rect 258264 305328 258316 305380
rect 259184 305328 259236 305380
rect 259736 305328 259788 305380
rect 260564 305328 260616 305380
rect 260840 305328 260892 305380
rect 261300 305328 261352 305380
rect 262220 305328 262272 305380
rect 262588 305328 262640 305380
rect 353300 305328 353352 305380
rect 365076 305396 365128 305448
rect 237748 305260 237800 305312
rect 238668 305260 238720 305312
rect 259552 305260 259604 305312
rect 260196 305260 260248 305312
rect 260932 305260 260984 305312
rect 261944 305260 261996 305312
rect 350816 305260 350868 305312
rect 358728 305260 358780 305312
rect 359464 305056 359516 305108
rect 360108 305056 360160 305108
rect 335452 304648 335504 304700
rect 336464 304648 336516 304700
rect 317420 304512 317472 304564
rect 318340 304512 318392 304564
rect 308588 304376 308640 304428
rect 390560 304376 390612 304428
rect 301044 304308 301096 304360
rect 301228 304308 301280 304360
rect 314108 304308 314160 304360
rect 418160 304308 418212 304360
rect 217416 304240 217468 304292
rect 352656 304240 352708 304292
rect 317604 304172 317656 304224
rect 317880 304172 317932 304224
rect 322940 304172 322992 304224
rect 323308 304172 323360 304224
rect 324596 304172 324648 304224
rect 325608 304172 325660 304224
rect 255320 304104 255372 304156
rect 255688 304104 255740 304156
rect 258080 303696 258132 303748
rect 258356 303696 258408 303748
rect 320272 303696 320324 303748
rect 320640 303696 320692 303748
rect 212448 303560 212500 303612
rect 280160 303560 280212 303612
rect 353576 303560 353628 303612
rect 372804 303560 372856 303612
rect 213552 303492 213604 303544
rect 282092 303492 282144 303544
rect 352380 303492 352432 303544
rect 372896 303492 372948 303544
rect 213092 303424 213144 303476
rect 282552 303424 282604 303476
rect 351736 303424 351788 303476
rect 371608 303424 371660 303476
rect 217968 303356 218020 303408
rect 288256 303356 288308 303408
rect 347596 303356 347648 303408
rect 371976 303356 372028 303408
rect 213644 303288 213696 303340
rect 283104 303288 283156 303340
rect 306656 303288 306708 303340
rect 379520 303288 379572 303340
rect 211068 303220 211120 303272
rect 282276 303220 282328 303272
rect 307208 303220 307260 303272
rect 382280 303220 382332 303272
rect 212356 303152 212408 303204
rect 283012 303152 283064 303204
rect 301044 303152 301096 303204
rect 301872 303152 301924 303204
rect 308036 303152 308088 303204
rect 386420 303152 386472 303204
rect 213368 303084 213420 303136
rect 346860 303084 346912 303136
rect 348516 303084 348568 303136
rect 370688 303084 370740 303136
rect 306564 303016 306616 303068
rect 307392 303016 307444 303068
rect 353116 303016 353168 303068
rect 374276 303016 374328 303068
rect 211896 302948 211948 303000
rect 347780 302948 347832 303000
rect 349620 302948 349672 303000
rect 372712 302948 372764 303000
rect 210608 302880 210660 302932
rect 348056 302880 348108 302932
rect 348700 302880 348752 302932
rect 374184 302880 374236 302932
rect 217876 302812 217928 302864
rect 283932 302812 283984 302864
rect 349436 302812 349488 302864
rect 367652 302812 367704 302864
rect 215944 302744 215996 302796
rect 280896 302744 280948 302796
rect 350356 302744 350408 302796
rect 366548 302744 366600 302796
rect 218796 302676 218848 302728
rect 281540 302676 281592 302728
rect 356336 302676 356388 302728
rect 370596 302676 370648 302728
rect 217508 302608 217560 302660
rect 351920 302608 351972 302660
rect 305276 302336 305328 302388
rect 305552 302336 305604 302388
rect 305644 301792 305696 301844
rect 375380 301792 375432 301844
rect 217600 301724 217652 301776
rect 345020 301724 345072 301776
rect 217048 301656 217100 301708
rect 350632 301656 350684 301708
rect 341616 301588 341668 301640
rect 560300 301588 560352 301640
rect 342812 301520 342864 301572
rect 564440 301520 564492 301572
rect 344376 301452 344428 301504
rect 574100 301452 574152 301504
rect 243176 300840 243228 300892
rect 243360 300840 243412 300892
rect 216036 300772 216088 300824
rect 285864 300772 285916 300824
rect 214380 300704 214432 300756
rect 285772 300704 285824 300756
rect 212172 300636 212224 300688
rect 284300 300636 284352 300688
rect 213184 300568 213236 300620
rect 280988 300568 281040 300620
rect 210976 300500 211028 300552
rect 284392 300500 284444 300552
rect 210884 300432 210936 300484
rect 284760 300432 284812 300484
rect 305368 300432 305420 300484
rect 372620 300432 372672 300484
rect 212264 300364 212316 300416
rect 285680 300364 285732 300416
rect 321928 300364 321980 300416
rect 456800 300364 456852 300416
rect 210516 300296 210568 300348
rect 350540 300296 350592 300348
rect 210700 300228 210752 300280
rect 284668 300228 284720 300280
rect 338580 300228 338632 300280
rect 542360 300228 542412 300280
rect 210792 300160 210844 300212
rect 284484 300160 284536 300212
rect 339776 300160 339828 300212
rect 549260 300160 549312 300212
rect 213460 300092 213512 300144
rect 288440 300092 288492 300144
rect 340236 300092 340288 300144
rect 553400 300092 553452 300144
rect 215852 300024 215904 300076
rect 286416 300024 286468 300076
rect 217784 299956 217836 300008
rect 283288 299956 283340 300008
rect 219348 299888 219400 299940
rect 284576 299888 284628 299940
rect 321008 298936 321060 298988
rect 454040 298936 454092 298988
rect 336096 298868 336148 298920
rect 531320 298868 531372 298920
rect 337200 298800 337252 298852
rect 535460 298800 535512 298852
rect 337108 298732 337160 298784
rect 539600 298732 539652 298784
rect 330668 297576 330720 297628
rect 503720 297576 503772 297628
rect 331680 297508 331732 297560
rect 506480 297508 506532 297560
rect 331588 297440 331640 297492
rect 510620 297440 510672 297492
rect 342628 297372 342680 297424
rect 567200 297372 567252 297424
rect 218612 296216 218664 296268
rect 349160 296216 349212 296268
rect 327540 296148 327592 296200
rect 489920 296148 489972 296200
rect 328920 296080 328972 296132
rect 492680 296080 492732 296132
rect 330116 296012 330168 296064
rect 499580 296012 499632 296064
rect 341248 295944 341300 295996
rect 556160 295944 556212 295996
rect 218520 294856 218572 294908
rect 348240 294856 348292 294908
rect 321836 294788 321888 294840
rect 463700 294788 463752 294840
rect 324688 294720 324740 294772
rect 473360 294720 473412 294772
rect 326068 294652 326120 294704
rect 481640 294652 481692 294704
rect 124220 294584 124272 294636
rect 256700 294584 256752 294636
rect 335728 294584 335780 294636
rect 528560 294584 528612 294636
rect 314936 293428 314988 293480
rect 427820 293428 427872 293480
rect 117320 293360 117372 293412
rect 255688 293360 255740 293412
rect 317880 293360 317932 293412
rect 441620 293360 441672 293412
rect 110420 293292 110472 293344
rect 254308 293292 254360 293344
rect 321744 293292 321796 293344
rect 459560 293292 459612 293344
rect 102140 293224 102192 293276
rect 252928 293224 252980 293276
rect 324596 293224 324648 293276
rect 477500 293224 477552 293276
rect 112444 292000 112496 292052
rect 251180 292000 251232 292052
rect 312084 292000 312136 292052
rect 409880 292000 409932 292052
rect 92480 291932 92532 291984
rect 250168 291932 250220 291984
rect 312176 291932 312228 291984
rect 414020 291932 414072 291984
rect 88340 291864 88392 291916
rect 249800 291864 249852 291916
rect 314844 291864 314896 291916
rect 423680 291864 423732 291916
rect 85580 291796 85632 291848
rect 248788 291796 248840 291848
rect 316316 291796 316368 291848
rect 434720 291796 434772 291848
rect 104164 290640 104216 290692
rect 247500 290640 247552 290692
rect 309416 290640 309468 290692
rect 398840 290640 398892 290692
rect 77300 290572 77352 290624
rect 247408 290572 247460 290624
rect 310704 290572 310756 290624
rect 402980 290572 403032 290624
rect 74540 290504 74592 290556
rect 246028 290504 246080 290556
rect 310796 290504 310848 290556
rect 407212 290504 407264 290556
rect 70400 290436 70452 290488
rect 246120 290436 246172 290488
rect 313648 290436 313700 290488
rect 420920 290436 420972 290488
rect 122840 289280 122892 289332
rect 255504 289280 255556 289332
rect 306656 289280 306708 289332
rect 382372 289280 382424 289332
rect 118700 289212 118752 289264
rect 255596 289212 255648 289264
rect 308036 289212 308088 289264
rect 391940 289212 391992 289264
rect 115940 289144 115992 289196
rect 254216 289144 254268 289196
rect 309324 289144 309376 289196
rect 396080 289144 396132 289196
rect 63500 289076 63552 289128
rect 244648 289076 244700 289128
rect 323308 289076 323360 289128
rect 470600 289076 470652 289128
rect 111800 287852 111852 287904
rect 254124 287852 254176 287904
rect 303988 287852 304040 287904
rect 371240 287852 371292 287904
rect 109040 287784 109092 287836
rect 252836 287784 252888 287836
rect 305276 287784 305328 287836
rect 374000 287784 374052 287836
rect 104900 287716 104952 287768
rect 252744 287716 252796 287768
rect 305184 287716 305236 287768
rect 378140 287716 378192 287768
rect 52460 287648 52512 287700
rect 241980 287648 242032 287700
rect 319260 287648 319312 287700
rect 445760 287648 445812 287700
rect 102232 286492 102284 286544
rect 251548 286492 251600 286544
rect 319168 286492 319220 286544
rect 447140 286492 447192 286544
rect 98000 286424 98052 286476
rect 251456 286424 251508 286476
rect 344008 286424 344060 286476
rect 543004 286424 543056 286476
rect 91100 286356 91152 286408
rect 250076 286356 250128 286408
rect 345204 286356 345256 286408
rect 552664 286356 552716 286408
rect 49700 286288 49752 286340
rect 241888 286288 241940 286340
rect 343916 286288 343968 286340
rect 569960 286288 570012 286340
rect 114560 285200 114612 285252
rect 254032 285200 254084 285252
rect 93860 285132 93912 285184
rect 249984 285132 250036 285184
rect 327448 285132 327500 285184
rect 485780 285132 485832 285184
rect 86960 285064 87012 285116
rect 248696 285064 248748 285116
rect 341156 285064 341208 285116
rect 538864 285064 538916 285116
rect 77392 284996 77444 285048
rect 247316 284996 247368 285048
rect 342444 284996 342496 285048
rect 563060 284996 563112 285048
rect 38660 284928 38712 284980
rect 239128 284928 239180 284980
rect 342536 284928 342588 284980
rect 565820 284928 565872 284980
rect 110512 283840 110564 283892
rect 254400 283840 254452 283892
rect 107660 283772 107712 283824
rect 252652 283772 252704 283824
rect 316224 283772 316276 283824
rect 431960 283772 432012 283824
rect 100760 283704 100812 283756
rect 251364 283704 251416 283756
rect 335636 283704 335688 283756
rect 531412 283704 531464 283756
rect 73160 283636 73212 283688
rect 245936 283636 245988 283688
rect 339684 283636 339736 283688
rect 547880 283636 547932 283688
rect 43536 283568 43588 283620
rect 240508 283568 240560 283620
rect 339776 283568 339828 283620
rect 552020 283568 552072 283620
rect 160100 282412 160152 282464
rect 264060 282412 264112 282464
rect 103520 282344 103572 282396
rect 253020 282344 253072 282396
rect 313556 282344 313608 282396
rect 416780 282344 416832 282396
rect 96620 282276 96672 282328
rect 251272 282276 251324 282328
rect 333060 282276 333112 282328
rect 516140 282276 516192 282328
rect 93952 282208 94004 282260
rect 249892 282208 249944 282260
rect 334440 282208 334492 282260
rect 520280 282208 520332 282260
rect 69020 282140 69072 282192
rect 245844 282140 245896 282192
rect 335544 282140 335596 282192
rect 527180 282140 527232 282192
rect 201500 281052 201552 281104
rect 272248 281052 272300 281104
rect 155960 280984 156012 281036
rect 262496 280984 262548 281036
rect 328828 280984 328880 281036
rect 498200 280984 498252 281036
rect 151820 280916 151872 280968
rect 262588 280916 262640 280968
rect 331404 280916 331456 280968
rect 506572 280916 506624 280968
rect 66260 280848 66312 280900
rect 244556 280848 244608 280900
rect 331496 280848 331548 280900
rect 509240 280848 509292 280900
rect 31760 280780 31812 280832
rect 237748 280780 237800 280832
rect 341064 280780 341116 280832
rect 556252 280780 556304 280832
rect 198740 279760 198792 279812
rect 270868 279760 270920 279812
rect 196624 279692 196676 279744
rect 270960 279692 271012 279744
rect 191840 279624 191892 279676
rect 269488 279624 269540 279676
rect 325976 279624 326028 279676
rect 484400 279624 484452 279676
rect 149060 279556 149112 279608
rect 261300 279556 261352 279608
rect 327356 279556 327408 279608
rect 491300 279556 491352 279608
rect 89720 279488 89772 279540
rect 250260 279488 250312 279540
rect 328736 279488 328788 279540
rect 495440 279488 495492 279540
rect 26884 279420 26936 279472
rect 236276 279420 236328 279472
rect 338488 279420 338540 279472
rect 545120 279420 545172 279472
rect 187700 278264 187752 278316
rect 269396 278264 269448 278316
rect 184940 278196 184992 278248
rect 268200 278196 268252 278248
rect 320548 278196 320600 278248
rect 455420 278196 455472 278248
rect 180800 278128 180852 278180
rect 268108 278128 268160 278180
rect 321652 278128 321704 278180
rect 462320 278128 462372 278180
rect 144920 278060 144972 278112
rect 261208 278060 261260 278112
rect 325884 278060 325936 278112
rect 481732 278060 481784 278112
rect 62120 277992 62172 278044
rect 244464 277992 244516 278044
rect 327264 277992 327316 278044
rect 488540 277992 488592 278044
rect 176660 276904 176712 276956
rect 266636 276904 266688 276956
rect 173900 276836 173952 276888
rect 266728 276836 266780 276888
rect 316132 276836 316184 276888
rect 433340 276836 433392 276888
rect 169760 276768 169812 276820
rect 265440 276768 265492 276820
rect 317788 276768 317840 276820
rect 437480 276768 437532 276820
rect 142160 276700 142212 276752
rect 259920 276700 259972 276752
rect 320456 276700 320508 276752
rect 451280 276700 451332 276752
rect 61384 276632 61436 276684
rect 243360 276632 243412 276684
rect 332968 276632 333020 276684
rect 513380 276632 513432 276684
rect 167000 275408 167052 275460
rect 265348 275408 265400 275460
rect 313372 275408 313424 275460
rect 415492 275408 415544 275460
rect 162860 275340 162912 275392
rect 263968 275340 264020 275392
rect 313464 275340 313516 275392
rect 419540 275340 419592 275392
rect 57244 275272 57296 275324
rect 243268 275272 243320 275324
rect 319076 275272 319128 275324
rect 448520 275272 448572 275324
rect 211804 274252 211856 274304
rect 272064 274252 272116 274304
rect 211160 274184 211212 274236
rect 273628 274184 273680 274236
rect 206284 274116 206336 274168
rect 272156 274116 272208 274168
rect 309232 274116 309284 274168
rect 398932 274116 398984 274168
rect 158720 274048 158772 274100
rect 262404 274048 262456 274100
rect 310612 274048 310664 274100
rect 401600 274048 401652 274100
rect 138020 273980 138072 274032
rect 259828 273980 259880 274032
rect 311992 273980 312044 274032
rect 412640 273980 412692 274032
rect 36544 273912 36596 273964
rect 239036 273912 239088 273964
rect 314752 273912 314804 273964
rect 426440 273912 426492 273964
rect 367744 273164 367796 273216
rect 580172 273164 580224 273216
rect 201592 272824 201644 272876
rect 270684 272824 270736 272876
rect 197360 272756 197412 272808
rect 270776 272756 270828 272808
rect 193220 272688 193272 272740
rect 269304 272688 269356 272740
rect 154580 272620 154632 272672
rect 262312 272620 262364 272672
rect 307944 272620 307996 272672
rect 387800 272620 387852 272672
rect 131120 272552 131172 272604
rect 258356 272552 258408 272604
rect 307852 272552 307904 272604
rect 390652 272552 390704 272604
rect 30380 272484 30432 272536
rect 237656 272484 237708 272536
rect 309140 272484 309192 272536
rect 394700 272484 394752 272536
rect 188344 271464 188396 271516
rect 268016 271464 268068 271516
rect 183560 271396 183612 271448
rect 267924 271396 267976 271448
rect 179420 271328 179472 271380
rect 266544 271328 266596 271380
rect 305092 271328 305144 271380
rect 376760 271328 376812 271380
rect 143540 271260 143592 271312
rect 259736 271260 259788 271312
rect 306472 271260 306524 271312
rect 380900 271260 380952 271312
rect 85672 271192 85724 271244
rect 248604 271192 248656 271244
rect 306564 271192 306616 271244
rect 383660 271192 383712 271244
rect 27620 271124 27672 271176
rect 237564 271124 237616 271176
rect 318984 271124 319036 271176
rect 444380 271124 444432 271176
rect 178776 270104 178828 270156
rect 266452 270104 266504 270156
rect 172520 270036 172572 270088
rect 265256 270036 265308 270088
rect 168380 269968 168432 270020
rect 265164 269968 265216 270020
rect 305000 269968 305052 270020
rect 374092 269968 374144 270020
rect 140780 269900 140832 269952
rect 259644 269900 259696 269952
rect 320364 269900 320416 269952
rect 449900 269900 449952 269952
rect 82820 269832 82872 269884
rect 248512 269832 248564 269884
rect 342352 269832 342404 269884
rect 520924 269832 520976 269884
rect 13820 269764 13872 269816
rect 235080 269764 235132 269816
rect 343824 269764 343876 269816
rect 525064 269764 525116 269816
rect 165620 268608 165672 268660
rect 263784 268608 263836 268660
rect 303712 268608 303764 268660
rect 365720 268608 365772 268660
rect 161480 268540 161532 268592
rect 263876 268540 263928 268592
rect 339500 268540 339552 268592
rect 508504 268540 508556 268592
rect 157340 268472 157392 268524
rect 262680 268472 262732 268524
rect 339592 268472 339644 268524
rect 516784 268472 516836 268524
rect 136640 268404 136692 268456
rect 258264 268404 258316 268456
rect 332876 268404 332928 268456
rect 514852 268404 514904 268456
rect 52552 268336 52604 268388
rect 241796 268336 241848 268388
rect 338396 268336 338448 268388
rect 547972 268336 548024 268388
rect 3240 267656 3292 267708
rect 228364 267656 228416 267708
rect 153200 267180 153252 267232
rect 260104 267180 260156 267232
rect 335452 267180 335504 267232
rect 496084 267180 496136 267232
rect 150440 267112 150492 267164
rect 261116 267112 261168 267164
rect 336924 267112 336976 267164
rect 502984 267112 503036 267164
rect 64880 267044 64932 267096
rect 244372 267044 244424 267096
rect 334348 267044 334400 267096
rect 523132 267044 523184 267096
rect 22100 266976 22152 267028
rect 236184 266976 236236 267028
rect 337016 266976 337068 267028
rect 539692 266976 539744 267028
rect 209780 265820 209832 265872
rect 273444 265820 273496 265872
rect 311900 265820 311952 265872
rect 408500 265820 408552 265872
rect 146300 265752 146352 265804
rect 261024 265752 261076 265804
rect 332784 265752 332836 265804
rect 440884 265752 440936 265804
rect 133880 265684 133932 265736
rect 258172 265684 258224 265736
rect 334256 265684 334308 265736
rect 446404 265684 446456 265736
rect 48320 265616 48372 265668
rect 241704 265616 241756 265668
rect 334164 265616 334216 265668
rect 525800 265616 525852 265668
rect 207020 264528 207072 264580
rect 271972 264528 272024 264580
rect 195980 264460 196032 264512
rect 270592 264460 270644 264512
rect 193312 264392 193364 264444
rect 269212 264392 269264 264444
rect 332692 264392 332744 264444
rect 432604 264392 432656 264444
rect 143632 264324 143684 264376
rect 259552 264324 259604 264376
rect 317696 264324 317748 264376
rect 440240 264324 440292 264376
rect 126980 264256 127032 264308
rect 257068 264256 257120 264308
rect 331220 264256 331272 264308
rect 507860 264256 507912 264308
rect 44180 264188 44232 264240
rect 240416 264188 240468 264240
rect 331312 264188 331364 264240
rect 512000 264188 512052 264240
rect 175280 263100 175332 263152
rect 253296 263100 253348 263152
rect 185032 263032 185084 263084
rect 267740 263032 267792 263084
rect 330024 263032 330076 263084
rect 417424 263032 417476 263084
rect 182180 262964 182232 263016
rect 267832 262964 267884 263016
rect 316040 262964 316092 263016
rect 432052 262964 432104 263016
rect 139400 262896 139452 262948
rect 259460 262896 259512 262948
rect 328644 262896 328696 262948
rect 498292 262896 498344 262948
rect 40040 262828 40092 262880
rect 240324 262828 240376 262880
rect 343732 262828 343784 262880
rect 575480 262828 575532 262880
rect 207664 261808 207716 261860
rect 266820 261808 266872 261860
rect 171140 261740 171192 261792
rect 264980 261740 265032 261792
rect 168472 261672 168524 261724
rect 265072 261672 265124 261724
rect 327080 261672 327132 261724
rect 487160 261672 487212 261724
rect 164240 261604 164292 261656
rect 263692 261604 263744 261656
rect 327172 261604 327224 261656
rect 490012 261604 490064 261656
rect 128360 261536 128412 261588
rect 256976 261536 257028 261588
rect 328552 261536 328604 261588
rect 494060 261536 494112 261588
rect 35256 261468 35308 261520
rect 238944 261468 238996 261520
rect 338304 261468 338356 261520
rect 543740 261468 543792 261520
rect 160192 260312 160244 260364
rect 263600 260312 263652 260364
rect 125600 260244 125652 260296
rect 256884 260244 256936 260296
rect 60740 260176 60792 260228
rect 244740 260176 244792 260228
rect 325792 260176 325844 260228
rect 483020 260176 483072 260228
rect 8300 260108 8352 260160
rect 233516 260108 233568 260160
rect 335360 260108 335412 260160
rect 529940 260108 529992 260160
rect 51080 258884 51132 258936
rect 241612 258884 241664 258936
rect 35900 258816 35952 258868
rect 238852 258816 238904 258868
rect 3700 258748 3752 258800
rect 231124 258748 231176 258800
rect 4804 258680 4856 258732
rect 231860 258680 231912 258732
rect 217140 257320 217192 257372
rect 345480 257320 345532 257372
rect 321560 256164 321612 256216
rect 460940 256164 460992 256216
rect 24860 256096 24912 256148
rect 236092 256096 236144 256148
rect 323216 256096 323268 256148
rect 465080 256096 465132 256148
rect 17224 256028 17276 256080
rect 234988 256028 235040 256080
rect 324412 256028 324464 256080
rect 474740 256028 474792 256080
rect 7564 255960 7616 256012
rect 233424 255960 233476 256012
rect 325700 255960 325752 256012
rect 478880 255960 478932 256012
rect 116584 254804 116636 254856
rect 240600 254804 240652 254856
rect 79324 254736 79376 254788
rect 243084 254736 243136 254788
rect 302424 254736 302476 254788
rect 361580 254736 361632 254788
rect 56600 254668 56652 254720
rect 243176 254668 243228 254720
rect 313280 254668 313332 254720
rect 385684 254668 385736 254720
rect 44272 254600 44324 254652
rect 240232 254600 240284 254652
rect 318892 254600 318944 254652
rect 443000 254600 443052 254652
rect 39304 254532 39356 254584
rect 239220 254532 239272 254584
rect 345388 254532 345440 254584
rect 578240 254532 578292 254584
rect 2780 254328 2832 254380
rect 4896 254328 4948 254380
rect 301228 253512 301280 253564
rect 361672 253512 361724 253564
rect 84200 253444 84252 253496
rect 248420 253444 248472 253496
rect 301320 253444 301372 253496
rect 365812 253444 365864 253496
rect 80060 253376 80112 253428
rect 247224 253376 247276 253428
rect 332600 253376 332652 253428
rect 517520 253376 517572 253428
rect 17960 253308 18012 253360
rect 234804 253308 234856 253360
rect 334072 253308 334124 253360
rect 521660 253308 521712 253360
rect 12440 253240 12492 253292
rect 234896 253240 234948 253292
rect 333980 253240 334032 253292
rect 524420 253240 524472 253292
rect 9680 253172 9732 253224
rect 233332 253172 233384 253224
rect 343640 253172 343692 253224
rect 571340 253172 571392 253224
rect 121460 252084 121512 252136
rect 255412 252084 255464 252136
rect 118792 252016 118844 252068
rect 255780 252016 255832 252068
rect 318800 252016 318852 252068
rect 448612 252016 448664 252068
rect 31024 251948 31076 252000
rect 237472 251948 237524 252000
rect 320272 251948 320324 252000
rect 452660 251948 452712 252000
rect 26240 251880 26292 251932
rect 237840 251880 237892 251932
rect 320180 251880 320232 251932
rect 456892 251880 456944 251932
rect 20720 251812 20772 251864
rect 236368 251812 236420 251864
rect 323032 251812 323084 251864
rect 466460 251812 466512 251864
rect 299756 251132 299808 251184
rect 364708 251132 364760 251184
rect 299940 251064 299992 251116
rect 366180 251064 366232 251116
rect 292948 250996 293000 251048
rect 360200 250996 360252 251048
rect 298284 250928 298336 250980
rect 365904 250928 365956 250980
rect 298376 250860 298428 250912
rect 366088 250860 366140 250912
rect 297180 250792 297232 250844
rect 366272 250792 366324 250844
rect 174544 250724 174596 250776
rect 251640 250724 251692 250776
rect 294144 250724 294196 250776
rect 363512 250724 363564 250776
rect 78680 250656 78732 250708
rect 247132 250656 247184 250708
rect 294052 250656 294104 250708
rect 365996 250656 366048 250708
rect 75920 250588 75972 250640
rect 247040 250588 247092 250640
rect 291568 250588 291620 250640
rect 368480 250588 368532 250640
rect 71780 250520 71832 250572
rect 245752 250520 245804 250572
rect 306380 250520 306432 250572
rect 385040 250520 385092 250572
rect 16580 250452 16632 250504
rect 234712 250452 234764 250504
rect 307760 250452 307812 250504
rect 389180 250452 389232 250504
rect 299848 250384 299900 250436
rect 362960 250384 363012 250436
rect 295800 250316 295852 250368
rect 358820 250316 358872 250368
rect 295708 250248 295760 250300
rect 357440 250248 357492 250300
rect 209872 249228 209924 249280
rect 273260 249228 273312 249280
rect 317512 249228 317564 249280
rect 436100 249228 436152 249280
rect 205640 249160 205692 249212
rect 272340 249160 272392 249212
rect 338120 249160 338172 249212
rect 534724 249160 534776 249212
rect 135260 249092 135312 249144
rect 258448 249092 258500 249144
rect 336832 249092 336884 249144
rect 534080 249092 534132 249144
rect 13084 249024 13136 249076
rect 234620 249024 234672 249076
rect 336740 249024 336792 249076
rect 538220 249024 538272 249076
rect 295616 248344 295668 248396
rect 361764 248344 361816 248396
rect 297088 248276 297140 248328
rect 363420 248276 363472 248328
rect 298100 248208 298152 248260
rect 364616 248208 364668 248260
rect 292672 248140 292724 248192
rect 359188 248140 359240 248192
rect 296996 248072 297048 248124
rect 364432 248072 364484 248124
rect 296812 248004 296864 248056
rect 364524 248004 364576 248056
rect 151912 247936 151964 247988
rect 260932 247936 260984 247988
rect 292764 247936 292816 247988
rect 360752 247936 360804 247988
rect 147680 247868 147732 247920
rect 260840 247868 260892 247920
rect 292856 247868 292908 247920
rect 362224 247868 362276 247920
rect 127072 247800 127124 247852
rect 256792 247800 256844 247852
rect 293960 247800 294012 247852
rect 368664 247800 368716 247852
rect 69112 247732 69164 247784
rect 245660 247732 245712 247784
rect 288808 247732 288860 247784
rect 367100 247732 367152 247784
rect 2780 247664 2832 247716
rect 232136 247664 232188 247716
rect 288716 247664 288768 247716
rect 368572 247664 368624 247716
rect 298192 247596 298244 247648
rect 364340 247596 364392 247648
rect 291476 247528 291528 247580
rect 356704 247528 356756 247580
rect 299664 247460 299716 247512
rect 364800 247460 364852 247512
rect 291384 246644 291436 246696
rect 366364 246644 366416 246696
rect 192484 246576 192536 246628
rect 269580 246576 269632 246628
rect 310520 246576 310572 246628
rect 405740 246576 405792 246628
rect 129740 246508 129792 246560
rect 257160 246508 257212 246560
rect 331864 246508 331916 246560
rect 430580 246508 430632 246560
rect 57980 246440 58032 246492
rect 242992 246440 243044 246492
rect 314660 246440 314712 246492
rect 423772 246440 423824 246492
rect 53840 246372 53892 246424
rect 242900 246372 242952 246424
rect 317420 246372 317472 246424
rect 440332 246372 440384 246424
rect 48964 246304 49016 246356
rect 241520 246304 241572 246356
rect 328460 246304 328512 246356
rect 496820 246304 496872 246356
rect 300952 245556 301004 245608
rect 357440 245556 357492 245608
rect 357256 245488 357308 245540
rect 369860 245488 369912 245540
rect 301044 245420 301096 245472
rect 362132 245420 362184 245472
rect 299572 245352 299624 245404
rect 363328 245352 363380 245404
rect 214840 245284 214892 245336
rect 288624 245284 288676 245336
rect 295340 245284 295392 245336
rect 360660 245284 360712 245336
rect 213000 245216 213052 245268
rect 288532 245216 288584 245268
rect 292580 245216 292632 245268
rect 357992 245216 358044 245268
rect 358084 245216 358136 245268
rect 369952 245216 370004 245268
rect 135352 245148 135404 245200
rect 253204 245148 253256 245200
rect 291292 245148 291344 245200
rect 367192 245148 367244 245200
rect 132500 245080 132552 245132
rect 257344 245080 257396 245132
rect 329840 245080 329892 245132
rect 502340 245080 502392 245132
rect 6920 245012 6972 245064
rect 233240 245012 233292 245064
rect 340972 245012 341024 245064
rect 557540 245012 557592 245064
rect 4896 244944 4948 244996
rect 232044 244944 232096 244996
rect 340880 244944 340932 244996
rect 561680 244944 561732 244996
rect 2872 244876 2924 244928
rect 231952 244876 232004 244928
rect 342260 244876 342312 244928
rect 564532 244876 564584 244928
rect 357072 244808 357124 244860
rect 364892 244808 364944 244860
rect 356980 244604 357032 244656
rect 363696 244604 363748 244656
rect 357164 244468 357216 244520
rect 362316 244468 362368 244520
rect 355324 244060 355376 244112
rect 362408 244060 362460 244112
rect 355416 243992 355468 244044
rect 359280 243992 359332 244044
rect 219164 243720 219216 243772
rect 287336 243720 287388 243772
rect 290004 243720 290056 243772
rect 358084 243720 358136 243772
rect 217232 243652 217284 243704
rect 286048 243652 286100 243704
rect 289820 243652 289872 243704
rect 360844 243652 360896 243704
rect 219256 243584 219308 243636
rect 288900 243584 288952 243636
rect 289912 243584 289964 243636
rect 363604 243584 363656 243636
rect 215760 243516 215812 243568
rect 287428 243516 287480 243568
rect 291200 243516 291252 243568
rect 364984 243516 365036 243568
rect 3332 215228 3384 215280
rect 210424 215228 210476 215280
rect 214380 195236 214432 195288
rect 217324 195236 217376 195288
rect 215760 193128 215812 193180
rect 217416 193128 217468 193180
rect 210516 193060 210568 193112
rect 216680 193060 216732 193112
rect 215852 189252 215904 189304
rect 218612 189252 218664 189304
rect 210608 188980 210660 189032
rect 216680 188980 216732 189032
rect 213000 169532 213052 169584
rect 217508 169532 217560 169584
rect 351920 159672 351972 159724
rect 357900 159672 357952 159724
rect 213092 159604 213144 159656
rect 256700 159604 256752 159656
rect 325884 159604 325936 159656
rect 357808 159604 357860 159656
rect 217876 159536 217928 159588
rect 263600 159536 263652 159588
rect 313280 159536 313332 159588
rect 356796 159536 356848 159588
rect 214472 159468 214524 159520
rect 260840 159468 260892 159520
rect 310980 159468 311032 159520
rect 359004 159468 359056 159520
rect 217784 159400 217836 159452
rect 264980 159400 265032 159452
rect 291108 159400 291160 159452
rect 359096 159400 359148 159452
rect 216128 159332 216180 159384
rect 284392 159332 284444 159384
rect 285680 159332 285732 159384
rect 360568 159332 360620 159384
rect 279240 159128 279292 159180
rect 363236 159196 363288 159248
rect 278136 159060 278188 159112
rect 363144 159128 363196 159180
rect 355232 159060 355284 159112
rect 361948 159060 362000 159112
rect 277032 158992 277084 159044
rect 362040 158992 362092 159044
rect 273352 158924 273404 158976
rect 360476 158924 360528 158976
rect 275836 158856 275888 158908
rect 355232 158856 355284 158908
rect 274456 158788 274508 158840
rect 361028 158856 361080 158908
rect 211896 158720 211948 158772
rect 239588 158720 239640 158772
rect 261116 158720 261168 158772
rect 359372 158788 359424 158840
rect 213368 158652 213420 158704
rect 238116 158652 238168 158704
rect 269948 158652 270000 158704
rect 291108 158652 291160 158704
rect 295984 158652 296036 158704
rect 357624 158720 357676 158772
rect 214564 158584 214616 158636
rect 233240 158584 233292 158636
rect 315856 158584 315908 158636
rect 361856 158584 361908 158636
rect 218980 158516 219032 158568
rect 238760 158516 238812 158568
rect 272248 158516 272300 158568
rect 285680 158516 285732 158568
rect 293592 158516 293644 158568
rect 351920 158516 351972 158568
rect 211988 158448 212040 158500
rect 237380 158448 237432 158500
rect 298560 158448 298612 158500
rect 358360 158448 358412 158500
rect 216404 158380 216456 158432
rect 242992 158380 243044 158432
rect 300952 158380 301004 158432
rect 358912 158380 358964 158432
rect 213276 158312 213328 158364
rect 241520 158312 241572 158364
rect 303528 158312 303580 158364
rect 358176 158312 358228 158364
rect 216496 158244 216548 158296
rect 245660 158244 245712 158296
rect 306104 158244 306156 158296
rect 358268 158244 358320 158296
rect 214656 158176 214708 158228
rect 247040 158176 247092 158228
rect 308680 158176 308732 158228
rect 360384 158176 360436 158228
rect 215944 158108 215996 158160
rect 248420 158108 248472 158160
rect 268752 158108 268804 158160
rect 310980 158108 311032 158160
rect 311072 158108 311124 158160
rect 360292 158108 360344 158160
rect 216312 158040 216364 158092
rect 249800 158040 249852 158092
rect 288256 158040 288308 158092
rect 313280 158040 313332 158092
rect 313464 158040 313516 158092
rect 359648 158040 359700 158092
rect 218704 157972 218756 158024
rect 252560 157972 252612 158024
rect 318616 157972 318668 158024
rect 359556 157972 359608 158024
rect 212080 157904 212132 157956
rect 230480 157904 230532 157956
rect 323400 157904 323452 157956
rect 363052 157904 363104 157956
rect 216220 157836 216272 157888
rect 229100 157836 229152 157888
rect 321008 157836 321060 157888
rect 359464 157836 359516 157888
rect 219072 157768 219124 157820
rect 231860 157768 231912 157820
rect 265440 157768 265492 157820
rect 325884 157768 325936 157820
rect 325976 157768 326028 157820
rect 360936 157768 360988 157820
rect 242440 157292 242492 157344
rect 372712 157292 372764 157344
rect 244648 157224 244700 157276
rect 370044 157224 370096 157276
rect 248328 157156 248380 157208
rect 369308 157156 369360 157208
rect 245568 157088 245620 157140
rect 363788 157088 363840 157140
rect 252376 157020 252428 157072
rect 369216 157020 369268 157072
rect 255872 156952 255924 157004
rect 367284 156952 367336 157004
rect 257252 156884 257304 156936
rect 367376 156884 367428 156936
rect 261760 156816 261812 156868
rect 370136 156816 370188 156868
rect 265992 156748 266044 156800
rect 372896 156748 372948 156800
rect 266544 156680 266596 156732
rect 368848 156680 368900 156732
rect 270960 156612 271012 156664
rect 372804 156612 372856 156664
rect 276112 156544 276164 156596
rect 371792 156544 371844 156596
rect 281080 156476 281132 156528
rect 371884 156476 371936 156528
rect 217968 156408 218020 156460
rect 285680 156408 285732 156460
rect 291016 156408 291068 156460
rect 371700 156408 371752 156460
rect 241428 155864 241480 155916
rect 374184 155864 374236 155916
rect 246672 155796 246724 155848
rect 370228 155796 370280 155848
rect 251088 155728 251140 155780
rect 371976 155728 372028 155780
rect 247960 155660 248012 155712
rect 368940 155660 368992 155712
rect 248696 155592 248748 155644
rect 370320 155592 370372 155644
rect 250444 155524 250496 155576
rect 369032 155524 369084 155576
rect 252468 155456 252520 155508
rect 370412 155456 370464 155508
rect 218796 155388 218848 155440
rect 251180 155388 251232 155440
rect 253480 155388 253532 155440
rect 365076 155388 365128 155440
rect 210792 155320 210844 155372
rect 267740 155320 267792 155372
rect 268384 155320 268436 155372
rect 374276 155320 374328 155372
rect 212172 155252 212224 155304
rect 271880 155252 271932 155304
rect 273720 155252 273772 155304
rect 371516 155252 371568 155304
rect 210700 155184 210752 155236
rect 270500 155184 270552 155236
rect 271328 155184 271380 155236
rect 368756 155184 368808 155236
rect 216036 155116 216088 155168
rect 277400 155116 277452 155168
rect 278504 155116 278556 155168
rect 371424 155116 371476 155168
rect 214748 155048 214800 155100
rect 282920 155048 282972 155100
rect 283656 155048 283708 155100
rect 371332 155048 371384 155100
rect 217232 154980 217284 155032
rect 278780 154980 278832 155032
rect 256240 154504 256292 154556
rect 367652 154504 367704 154556
rect 263692 154436 263744 154488
rect 371608 154436 371660 154488
rect 286048 154368 286100 154420
rect 370596 154368 370648 154420
rect 218612 152600 218664 152652
rect 276112 152600 276164 152652
rect 212264 152532 212316 152584
rect 273260 152532 273312 152584
rect 213460 152464 213512 152516
rect 288440 152464 288492 152516
rect 3516 150356 3568 150408
rect 43444 150356 43496 150408
rect 3516 137912 3568 137964
rect 180064 137912 180116 137964
rect 143540 11704 143592 11756
rect 144736 11704 144788 11756
rect 168380 11704 168432 11756
rect 169576 11704 169628 11756
rect 201500 11704 201552 11756
rect 202696 11704 202748 11756
rect 234620 11704 234672 11756
rect 235816 11704 235868 11756
rect 151728 9596 151780 9648
rect 153016 9596 153068 9648
rect 209688 9596 209740 9648
rect 210976 9596 211028 9648
rect 300768 9596 300820 9648
rect 360844 9596 360896 9648
rect 301964 9528 302016 9580
rect 362408 9528 362460 9580
rect 309048 9460 309100 9512
rect 369860 9460 369912 9512
rect 306748 9392 306800 9444
rect 368480 9392 368532 9444
rect 305552 9324 305604 9376
rect 367192 9324 367244 9376
rect 304356 9256 304408 9308
rect 366364 9256 366416 9308
rect 303160 9188 303212 9240
rect 364984 9188 365036 9240
rect 296076 9120 296128 9172
rect 358084 9120 358136 9172
rect 299664 9052 299716 9104
rect 362316 9052 362368 9104
rect 294880 8984 294932 9036
rect 369952 8984 370004 9036
rect 293684 8916 293736 8968
rect 368572 8916 368624 8968
rect 298468 8848 298520 8900
rect 359280 8848 359332 8900
rect 312636 8780 312688 8832
rect 360752 8780 360804 8832
rect 316224 8712 316276 8764
rect 363512 8712 363564 8764
rect 330392 6808 330444 6860
rect 363420 6808 363472 6860
rect 333888 6740 333940 6792
rect 366272 6740 366324 6792
rect 323308 6672 323360 6724
rect 357532 6672 357584 6724
rect 313832 6604 313884 6656
rect 360200 6604 360252 6656
rect 319720 6536 319772 6588
rect 365996 6536 366048 6588
rect 318524 6468 318576 6520
rect 364892 6468 364944 6520
rect 317328 6400 317380 6452
rect 363696 6400 363748 6452
rect 315028 6332 315080 6384
rect 362224 6332 362276 6384
rect 311440 6264 311492 6316
rect 359188 6264 359240 6316
rect 310244 6196 310296 6248
rect 357992 6196 358044 6248
rect 292580 6128 292632 6180
rect 367100 6128 367152 6180
rect 326804 6060 326856 6112
rect 358820 6060 358872 6112
rect 337476 5992 337528 6044
rect 366088 5992 366140 6044
rect 340972 5924 341024 5976
rect 365904 5924 365956 5976
rect 6460 4088 6512 4140
rect 7564 4088 7616 4140
rect 15936 4088 15988 4140
rect 17224 4088 17276 4140
rect 24216 4088 24268 4140
rect 26884 4088 26936 4140
rect 213644 4088 213696 4140
rect 220452 4088 220504 4140
rect 34796 4020 34848 4072
rect 36544 4020 36596 4072
rect 213736 4020 213788 4072
rect 258264 4088 258316 4140
rect 355232 4088 355284 4140
rect 365812 4088 365864 4140
rect 220820 4020 220872 4072
rect 260656 4020 260708 4072
rect 350448 4020 350500 4072
rect 362960 4020 363012 4072
rect 219348 3952 219400 4004
rect 266544 3952 266596 4004
rect 349252 3952 349304 4004
rect 363328 3952 363380 4004
rect 214932 3884 214984 3936
rect 262956 3884 263008 3936
rect 343364 3884 343416 3936
rect 364340 3884 364392 3936
rect 503076 3884 503128 3936
rect 537208 3884 537260 3936
rect 217324 3816 217376 3868
rect 276020 3816 276072 3868
rect 339868 3816 339920 3868
rect 364616 3816 364668 3868
rect 496084 3816 496136 3868
rect 533712 3816 533764 3868
rect 538864 3816 538916 3868
rect 559748 3816 559800 3868
rect 219164 3748 219216 3800
rect 280712 3748 280764 3800
rect 336280 3748 336332 3800
rect 364524 3748 364576 3800
rect 516784 3748 516836 3800
rect 43076 3680 43128 3732
rect 50344 3680 50396 3732
rect 217416 3680 217468 3732
rect 284300 3680 284352 3732
rect 332692 3680 332744 3732
rect 364432 3680 364484 3732
rect 508504 3680 508556 3732
rect 551468 3680 551520 3732
rect 11152 3612 11204 3664
rect 12348 3544 12400 3596
rect 13084 3544 13136 3596
rect 35164 3612 35216 3664
rect 35992 3612 36044 3664
rect 46204 3612 46256 3664
rect 46664 3612 46716 3664
rect 30104 3544 30156 3596
rect 31024 3544 31076 3596
rect 33600 3544 33652 3596
rect 35256 3544 35308 3596
rect 52460 3544 52512 3596
rect 53380 3544 53432 3596
rect 60832 3612 60884 3664
rect 79324 3612 79376 3664
rect 96252 3612 96304 3664
rect 112444 3612 112496 3664
rect 114008 3612 114060 3664
rect 182824 3612 182876 3664
rect 116584 3544 116636 3596
rect 118700 3544 118752 3596
rect 119896 3544 119948 3596
rect 121092 3544 121144 3596
rect 189724 3612 189776 3664
rect 213828 3612 213880 3664
rect 281908 3612 281960 3664
rect 329196 3612 329248 3664
rect 361764 3612 361816 3664
rect 446404 3612 446456 3664
rect 523040 3612 523092 3664
rect 543004 3612 543056 3664
rect 552572 3612 552624 3664
rect 187332 3544 187384 3596
rect 188344 3544 188396 3596
rect 193220 3544 193272 3596
rect 194416 3544 194468 3596
rect 195612 3544 195664 3596
rect 196624 3544 196676 3596
rect 208584 3544 208636 3596
rect 211804 3544 211856 3596
rect 219256 3544 219308 3596
rect 287796 3544 287848 3596
rect 328000 3544 328052 3596
rect 360660 3544 360712 3596
rect 385684 3544 385736 3596
rect 398840 3544 398892 3596
rect 400128 3544 400180 3596
rect 572 3476 624 3528
rect 4804 3476 4856 3528
rect 5264 3476 5316 3528
rect 75184 3476 75236 3528
rect 77300 3476 77352 3528
rect 78220 3476 78272 3528
rect 82084 3476 82136 3528
rect 104164 3476 104216 3528
rect 106924 3476 106976 3528
rect 2780 3408 2832 3460
rect 3700 3408 3752 3460
rect 20628 3408 20680 3460
rect 68284 3408 68336 3460
rect 69020 3408 69072 3460
rect 69940 3408 69992 3460
rect 93860 3408 93912 3460
rect 94780 3408 94832 3460
rect 102140 3408 102192 3460
rect 103336 3408 103388 3460
rect 28908 3340 28960 3392
rect 32404 3340 32456 3392
rect 56048 3340 56100 3392
rect 57244 3340 57296 3392
rect 59636 3340 59688 3392
rect 61384 3340 61436 3392
rect 99840 3340 99892 3392
rect 174544 3408 174596 3460
rect 176660 3476 176712 3528
rect 177856 3476 177908 3528
rect 190828 3476 190880 3528
rect 192484 3476 192536 3528
rect 205088 3476 205140 3528
rect 206284 3476 206336 3528
rect 217508 3476 217560 3528
rect 291384 3476 291436 3528
rect 307944 3476 307996 3528
rect 356704 3476 356756 3528
rect 365720 3476 365772 3528
rect 367008 3476 367060 3528
rect 374000 3476 374052 3528
rect 375288 3476 375340 3528
rect 382280 3476 382332 3528
rect 383568 3476 383620 3528
rect 178684 3408 178736 3460
rect 179052 3408 179104 3460
rect 207664 3408 207716 3460
rect 214840 3408 214892 3460
rect 290188 3408 290240 3460
rect 297272 3408 297324 3460
rect 363604 3408 363656 3460
rect 390652 3476 390704 3528
rect 391848 3476 391900 3528
rect 392676 3476 392728 3528
rect 426164 3544 426216 3596
rect 432604 3544 432656 3596
rect 415492 3476 415544 3528
rect 416688 3476 416740 3528
rect 423680 3476 423732 3528
rect 424968 3476 425020 3528
rect 432052 3476 432104 3528
rect 433248 3476 433300 3528
rect 440884 3544 440936 3596
rect 519544 3544 519596 3596
rect 525064 3544 525116 3596
rect 531320 3544 531372 3596
rect 532148 3544 532200 3596
rect 534724 3544 534776 3596
rect 541992 3544 542044 3596
rect 547880 3544 547932 3596
rect 548708 3544 548760 3596
rect 552756 3748 552808 3800
rect 554044 3680 554096 3732
rect 558184 3748 558236 3800
rect 583392 3748 583444 3800
rect 554964 3544 555016 3596
rect 556160 3544 556212 3596
rect 556988 3544 557040 3596
rect 577412 3680 577464 3732
rect 557172 3612 557224 3664
rect 573916 3612 573968 3664
rect 582196 3544 582248 3596
rect 515956 3476 516008 3528
rect 572720 3476 572772 3528
rect 417516 3408 417568 3460
rect 505376 3408 505428 3460
rect 506480 3408 506532 3460
rect 507308 3408 507360 3460
rect 520924 3408 520976 3460
rect 569132 3408 569184 3460
rect 212448 3340 212500 3392
rect 245200 3340 245252 3392
rect 251180 3340 251232 3392
rect 252376 3340 252428 3392
rect 352840 3340 352892 3392
rect 363880 3340 363932 3392
rect 415492 3340 415544 3392
rect 440332 3340 440384 3392
rect 441528 3340 441580 3392
rect 448612 3340 448664 3392
rect 449808 3340 449860 3392
rect 456800 3340 456852 3392
rect 458088 3340 458140 3392
rect 473360 3340 473412 3392
rect 474188 3340 474240 3392
rect 481640 3340 481692 3392
rect 482468 3340 482520 3392
rect 498200 3340 498252 3392
rect 499028 3340 499080 3392
rect 552572 3340 552624 3392
rect 557172 3340 557224 3392
rect 215208 3272 215260 3324
rect 242900 3272 242952 3324
rect 354036 3272 354088 3324
rect 361028 3272 361080 3324
rect 47860 3204 47912 3256
rect 48964 3204 49016 3256
rect 215024 3204 215076 3256
rect 240508 3204 240560 3256
rect 1676 3136 1728 3188
rect 4896 3136 4948 3188
rect 38384 3136 38436 3188
rect 39304 3136 39356 3188
rect 176660 3000 176712 3052
rect 178776 3000 178828 3052
rect 356336 3000 356388 3052
rect 362132 3000 362184 3052
rect 19432 2932 19484 2984
rect 25504 2932 25556 2984
rect 41880 2864 41932 2916
rect 43536 2864 43588 2916
rect 407120 2184 407172 2236
rect 408408 2184 408460 2236
<< metal2 >>
rect 6932 703582 7972 703610
rect 2778 684312 2834 684321
rect 2778 684247 2834 684256
rect 2792 683738 2820 684247
rect 2780 683732 2832 683738
rect 2780 683674 2832 683680
rect 4804 683732 4856 683738
rect 4804 683674 4856 683680
rect 3422 671256 3478 671265
rect 3422 671191 3478 671200
rect 2780 632120 2832 632126
rect 2778 632088 2780 632097
rect 2832 632088 2834 632097
rect 2778 632023 2834 632032
rect 3330 606112 3386 606121
rect 3330 606047 3386 606056
rect 3344 605878 3372 606047
rect 3332 605872 3384 605878
rect 3332 605814 3384 605820
rect 2778 580000 2834 580009
rect 2778 579935 2780 579944
rect 2832 579935 2834 579944
rect 2780 579906 2832 579912
rect 3054 566944 3110 566953
rect 3054 566879 3110 566888
rect 3068 565894 3096 566879
rect 3056 565888 3108 565894
rect 3056 565830 3108 565836
rect 2778 553888 2834 553897
rect 2778 553823 2834 553832
rect 2792 553722 2820 553823
rect 2780 553716 2832 553722
rect 2780 553658 2832 553664
rect 3330 527912 3386 527921
rect 3330 527847 3386 527856
rect 3344 527814 3372 527847
rect 3332 527808 3384 527814
rect 3332 527750 3384 527756
rect 3330 475688 3386 475697
rect 3330 475623 3386 475632
rect 3344 474774 3372 475623
rect 3332 474768 3384 474774
rect 3332 474710 3384 474716
rect 3436 470594 3464 671191
rect 3514 658200 3570 658209
rect 3514 658135 3570 658144
rect 3528 656946 3556 658135
rect 3516 656940 3568 656946
rect 3516 656882 3568 656888
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3344 470566 3464 470594
rect 3344 454850 3372 470566
rect 3422 462632 3478 462641
rect 3422 462567 3478 462576
rect 3436 462398 3464 462567
rect 3424 462392 3476 462398
rect 3424 462334 3476 462340
rect 3332 454844 3384 454850
rect 3332 454786 3384 454792
rect 3528 454782 3556 619103
rect 3606 514856 3662 514865
rect 3606 514791 3662 514800
rect 3620 456074 3648 514791
rect 3698 501800 3754 501809
rect 3698 501735 3754 501744
rect 3712 478174 3740 501735
rect 3700 478168 3752 478174
rect 3700 478110 3752 478116
rect 3608 456068 3660 456074
rect 3608 456010 3660 456016
rect 3516 454776 3568 454782
rect 3516 454718 3568 454724
rect 4816 450634 4844 683674
rect 4896 632120 4948 632126
rect 4896 632062 4948 632068
rect 4804 450628 4856 450634
rect 4804 450570 4856 450576
rect 4908 450566 4936 632062
rect 4988 579964 5040 579970
rect 4988 579906 5040 579912
rect 5000 451926 5028 579906
rect 5080 553716 5132 553722
rect 5080 553658 5132 553664
rect 5092 454714 5120 553658
rect 5080 454708 5132 454714
rect 5080 454650 5132 454656
rect 6932 453354 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 23492 703582 24164 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 8944 527808 8996 527814
rect 8944 527750 8996 527756
rect 6920 453348 6972 453354
rect 6920 453290 6972 453296
rect 8956 451994 8984 527750
rect 8944 451988 8996 451994
rect 8944 451930 8996 451936
rect 4988 451920 5040 451926
rect 4988 451862 5040 451868
rect 4896 450560 4948 450566
rect 4896 450502 4948 450508
rect 2870 449576 2926 449585
rect 2870 449511 2926 449520
rect 2884 447846 2912 449511
rect 23492 449206 23520 703582
rect 24136 703474 24164 703582
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 24320 703474 24348 703520
rect 24136 703446 24348 703474
rect 31024 565888 31076 565894
rect 31024 565830 31076 565836
rect 31036 454918 31064 565830
rect 31024 454912 31076 454918
rect 31024 454854 31076 454860
rect 23480 449200 23532 449206
rect 23480 449142 23532 449148
rect 40052 447914 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 71792 452062 71820 702986
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 71780 452056 71832 452062
rect 71780 451998 71832 452004
rect 88352 449342 88380 702406
rect 88340 449336 88392 449342
rect 88340 449278 88392 449284
rect 104912 447982 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 136652 448050 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 702434 154160 703520
rect 170324 702434 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 153212 702406 154160 702434
rect 169772 702406 170352 702434
rect 153212 449478 153240 702406
rect 153200 449472 153252 449478
rect 153200 449414 153252 449420
rect 169772 448118 169800 702406
rect 178684 656940 178736 656946
rect 178684 656882 178736 656888
rect 178696 453422 178724 656882
rect 178684 453416 178736 453422
rect 178684 453358 178736 453364
rect 201512 448186 201540 702986
rect 203524 605872 203576 605878
rect 203524 605814 203576 605820
rect 203536 453490 203564 605814
rect 217968 565140 218020 565146
rect 217968 565082 218020 565088
rect 217874 516896 217930 516905
rect 217874 516831 217930 516840
rect 217598 515944 217654 515953
rect 217598 515879 217654 515888
rect 217506 513768 217562 513777
rect 217506 513703 217562 513712
rect 217414 488336 217470 488345
rect 217414 488271 217470 488280
rect 217428 478922 217456 488271
rect 217416 478916 217468 478922
rect 217416 478858 217468 478864
rect 217520 474026 217548 513703
rect 217612 475386 217640 515879
rect 217690 489968 217746 489977
rect 217690 489903 217746 489912
rect 217600 475380 217652 475386
rect 217600 475322 217652 475328
rect 217508 474020 217560 474026
rect 217508 473962 217560 473968
rect 203524 453484 203576 453490
rect 203524 453426 203576 453432
rect 217704 450702 217732 489903
rect 217782 488064 217838 488073
rect 217782 487999 217838 488008
rect 217692 450696 217744 450702
rect 217692 450638 217744 450644
rect 201500 448180 201552 448186
rect 201500 448122 201552 448128
rect 169760 448112 169812 448118
rect 169760 448054 169812 448060
rect 136640 448044 136692 448050
rect 136640 447986 136692 447992
rect 104900 447976 104952 447982
rect 104900 447918 104952 447924
rect 40040 447908 40092 447914
rect 40040 447850 40092 447856
rect 2872 447840 2924 447846
rect 2872 447782 2924 447788
rect 210424 446820 210476 446826
rect 210424 446762 210476 446768
rect 4896 445188 4948 445194
rect 4896 445130 4948 445136
rect 3884 445052 3936 445058
rect 3884 444994 3936 445000
rect 3792 443964 3844 443970
rect 3792 443906 3844 443912
rect 3516 443896 3568 443902
rect 3516 443838 3568 443844
rect 3424 434036 3476 434042
rect 3424 433978 3476 433984
rect 3332 423632 3384 423638
rect 3330 423600 3332 423609
rect 3384 423600 3386 423609
rect 3330 423535 3386 423544
rect 3332 411256 3384 411262
rect 3332 411198 3384 411204
rect 3344 410553 3372 411198
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 3332 372564 3384 372570
rect 3332 372506 3384 372512
rect 3344 371385 3372 372506
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 3332 358760 3384 358766
rect 3332 358702 3384 358708
rect 3344 358465 3372 358702
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3332 320136 3384 320142
rect 3332 320078 3384 320084
rect 3344 319297 3372 320078
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3240 267708 3292 267714
rect 3240 267650 3292 267656
rect 3252 267209 3280 267650
rect 3238 267200 3294 267209
rect 3238 267135 3294 267144
rect 2780 254380 2832 254386
rect 2780 254322 2832 254328
rect 2792 254153 2820 254322
rect 2778 254144 2834 254153
rect 2778 254079 2834 254088
rect 2780 247716 2832 247722
rect 2780 247658 2832 247664
rect 572 3528 624 3534
rect 572 3470 624 3476
rect 584 480 612 3470
rect 2792 3466 2820 247658
rect 2872 244928 2924 244934
rect 2872 244870 2924 244876
rect 2780 3460 2832 3466
rect 2780 3402 2832 3408
rect 1676 3188 1728 3194
rect 1676 3130 1728 3136
rect 1688 480 1716 3130
rect 2884 480 2912 244870
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3436 97617 3464 433978
rect 3528 188873 3556 443838
rect 3608 443828 3660 443834
rect 3608 443770 3660 443776
rect 3620 241097 3648 443770
rect 3700 443692 3752 443698
rect 3700 443634 3752 443640
rect 3712 293185 3740 443634
rect 3804 306241 3832 443906
rect 3896 345409 3924 444994
rect 3976 443760 4028 443766
rect 3976 443702 4028 443708
rect 3988 397497 4016 443702
rect 3974 397488 4030 397497
rect 3974 397423 4030 397432
rect 3882 345400 3938 345409
rect 3882 345335 3938 345344
rect 3790 306232 3846 306241
rect 3790 306167 3846 306176
rect 3698 293176 3754 293185
rect 3698 293111 3754 293120
rect 3700 258800 3752 258806
rect 3700 258742 3752 258748
rect 3606 241088 3662 241097
rect 3606 241023 3662 241032
rect 3712 201929 3740 258742
rect 4804 258732 4856 258738
rect 4804 258674 4856 258680
rect 3698 201920 3754 201929
rect 3698 201855 3754 201864
rect 3514 188864 3570 188873
rect 3514 188799 3570 188808
rect 3516 150408 3568 150414
rect 3516 150350 3568 150356
rect 3528 149841 3556 150350
rect 3514 149832 3570 149841
rect 3514 149767 3570 149776
rect 3516 137964 3568 137970
rect 3516 137906 3568 137912
rect 3528 136785 3556 137906
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 4816 3534 4844 258674
rect 4908 254386 4936 445130
rect 40684 445120 40736 445126
rect 40684 445062 40736 445068
rect 40696 423638 40724 445062
rect 174544 444712 174596 444718
rect 174544 444654 174596 444660
rect 106924 444644 106976 444650
rect 106924 444586 106976 444592
rect 43444 444508 43496 444514
rect 43444 444450 43496 444456
rect 40684 423632 40736 423638
rect 40684 423574 40736 423580
rect 32404 308508 32456 308514
rect 32404 308450 32456 308456
rect 25504 308440 25556 308446
rect 25504 308382 25556 308388
rect 13820 269816 13872 269822
rect 13820 269758 13872 269764
rect 8300 260160 8352 260166
rect 8300 260102 8352 260108
rect 7564 256012 7616 256018
rect 7564 255954 7616 255960
rect 4896 254380 4948 254386
rect 4896 254322 4948 254328
rect 6920 245064 6972 245070
rect 6920 245006 6972 245012
rect 4896 244996 4948 245002
rect 4896 244938 4948 244944
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 3700 3460 3752 3466
rect 3700 3402 3752 3408
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3712 354 3740 3402
rect 4908 3194 4936 244938
rect 6932 16574 6960 245006
rect 6932 16546 7512 16574
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 4896 3188 4948 3194
rect 4896 3130 4948 3136
rect 5276 480 5304 3470
rect 6472 480 6500 4082
rect 7484 3482 7512 16546
rect 7576 4146 7604 255954
rect 8312 16574 8340 260102
rect 12440 253292 12492 253298
rect 12440 253234 12492 253240
rect 9680 253224 9732 253230
rect 9680 253166 9732 253172
rect 8312 16546 8800 16574
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7484 3454 7696 3482
rect 7668 480 7696 3454
rect 8772 480 8800 16546
rect 4038 354 4150 480
rect 3712 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 253166
rect 12452 16574 12480 253234
rect 13084 249076 13136 249082
rect 13084 249018 13136 249024
rect 12452 16546 13032 16574
rect 11152 3664 11204 3670
rect 11152 3606 11204 3612
rect 11164 480 11192 3606
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 12360 480 12388 3538
rect 13004 3482 13032 16546
rect 13096 3602 13124 249018
rect 13832 16574 13860 269758
rect 22100 267028 22152 267034
rect 22100 266970 22152 266976
rect 17224 256080 17276 256086
rect 17224 256022 17276 256028
rect 16580 250504 16632 250510
rect 16580 250446 16632 250452
rect 16592 16574 16620 250446
rect 13832 16546 14320 16574
rect 16592 16546 17080 16574
rect 13084 3596 13136 3602
rect 13084 3538 13136 3544
rect 13004 3454 13584 3482
rect 13556 480 13584 3454
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 15936 4140 15988 4146
rect 15936 4082 15988 4088
rect 15948 480 15976 4082
rect 17052 480 17080 16546
rect 17236 4146 17264 256022
rect 17960 253360 18012 253366
rect 17960 253302 18012 253308
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 253302
rect 20720 251864 20772 251870
rect 20720 251806 20772 251812
rect 20732 16574 20760 251806
rect 22112 16574 22140 266970
rect 24860 256148 24912 256154
rect 24860 256090 24912 256096
rect 24872 16574 24900 256090
rect 20732 16546 21864 16574
rect 22112 16546 22600 16574
rect 24872 16546 25360 16574
rect 20628 3460 20680 3466
rect 20628 3402 20680 3408
rect 19432 2984 19484 2990
rect 19432 2926 19484 2932
rect 19444 480 19472 2926
rect 20640 480 20668 3402
rect 21836 480 21864 16546
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 24216 4140 24268 4146
rect 24216 4082 24268 4088
rect 24228 480 24256 4082
rect 25332 480 25360 16546
rect 25516 2990 25544 308382
rect 31760 280832 31812 280838
rect 31760 280774 31812 280780
rect 26884 279472 26936 279478
rect 26884 279414 26936 279420
rect 26240 251932 26292 251938
rect 26240 251874 26292 251880
rect 25504 2984 25556 2990
rect 25504 2926 25556 2932
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 251874
rect 26896 4146 26924 279414
rect 30380 272536 30432 272542
rect 30380 272478 30432 272484
rect 27620 271176 27672 271182
rect 27620 271118 27672 271124
rect 27632 16574 27660 271118
rect 30392 16574 30420 272478
rect 31024 252000 31076 252006
rect 31024 251942 31076 251948
rect 27632 16546 27752 16574
rect 30392 16546 30880 16574
rect 26884 4140 26936 4146
rect 26884 4082 26936 4088
rect 27724 480 27752 16546
rect 30104 3596 30156 3602
rect 30104 3538 30156 3544
rect 28908 3392 28960 3398
rect 28908 3334 28960 3340
rect 28920 480 28948 3334
rect 30116 480 30144 3538
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31036 3602 31064 251942
rect 31772 16574 31800 280774
rect 31772 16546 31984 16574
rect 31024 3596 31076 3602
rect 31024 3538 31076 3544
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 32416 3398 32444 308450
rect 35162 308408 35218 308417
rect 35162 308343 35218 308352
rect 34796 4072 34848 4078
rect 34796 4014 34848 4020
rect 33600 3596 33652 3602
rect 33600 3538 33652 3544
rect 32404 3392 32456 3398
rect 32404 3334 32456 3340
rect 33612 480 33640 3538
rect 34808 480 34836 4014
rect 35176 3670 35204 308343
rect 38660 284980 38712 284986
rect 38660 284922 38712 284928
rect 36544 273964 36596 273970
rect 36544 273906 36596 273912
rect 35256 261520 35308 261526
rect 35256 261462 35308 261468
rect 35164 3664 35216 3670
rect 35164 3606 35216 3612
rect 35268 3602 35296 261462
rect 35900 258868 35952 258874
rect 35900 258810 35952 258816
rect 35912 16574 35940 258810
rect 35912 16546 36492 16574
rect 35992 3664 36044 3670
rect 35992 3606 36044 3612
rect 35256 3596 35308 3602
rect 35256 3538 35308 3544
rect 36004 480 36032 3606
rect 36464 490 36492 16546
rect 36556 4078 36584 273906
rect 38672 16574 38700 284922
rect 40040 262880 40092 262886
rect 40040 262822 40092 262828
rect 39304 254584 39356 254590
rect 39304 254526 39356 254532
rect 38672 16546 39160 16574
rect 36544 4072 36596 4078
rect 36544 4014 36596 4020
rect 38384 3188 38436 3194
rect 38384 3130 38436 3136
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 36464 462 36860 490
rect 38396 480 38424 3130
rect 36832 354 36860 462
rect 37158 354 37270 480
rect 36832 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 39316 3194 39344 254526
rect 40052 16574 40080 262822
rect 43456 150414 43484 444450
rect 106936 372570 106964 444586
rect 106924 372564 106976 372570
rect 106924 372506 106976 372512
rect 174556 320142 174584 444654
rect 180064 443148 180116 443154
rect 180064 443090 180116 443096
rect 174544 320136 174596 320142
rect 174544 320078 174596 320084
rect 178684 308780 178736 308786
rect 178684 308722 178736 308728
rect 68284 308712 68336 308718
rect 68284 308654 68336 308660
rect 50344 308644 50396 308650
rect 50344 308586 50396 308592
rect 46204 308576 46256 308582
rect 46204 308518 46256 308524
rect 43536 283620 43588 283626
rect 43536 283562 43588 283568
rect 43444 150408 43496 150414
rect 43444 150350 43496 150356
rect 40052 16546 40264 16574
rect 39304 3188 39356 3194
rect 39304 3130 39356 3136
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 43076 3732 43128 3738
rect 43076 3674 43128 3680
rect 41880 2916 41932 2922
rect 41880 2858 41932 2864
rect 41892 480 41920 2858
rect 43088 480 43116 3674
rect 43548 2922 43576 283562
rect 44180 264240 44232 264246
rect 44180 264182 44232 264188
rect 44192 6914 44220 264182
rect 44272 254652 44324 254658
rect 44272 254594 44324 254600
rect 44284 16574 44312 254594
rect 44284 16546 45048 16574
rect 44192 6886 44312 6914
rect 43536 2916 43588 2922
rect 43536 2858 43588 2864
rect 44284 480 44312 6886
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45020 354 45048 16546
rect 46216 3670 46244 308518
rect 49700 286340 49752 286346
rect 49700 286282 49752 286288
rect 48320 265668 48372 265674
rect 48320 265610 48372 265616
rect 48332 16574 48360 265610
rect 48964 246356 49016 246362
rect 48964 246298 49016 246304
rect 48332 16546 48544 16574
rect 46204 3664 46256 3670
rect 46204 3606 46256 3612
rect 46664 3664 46716 3670
rect 46664 3606 46716 3612
rect 46676 480 46704 3606
rect 47860 3256 47912 3262
rect 47860 3198 47912 3204
rect 47872 480 47900 3198
rect 45438 354 45550 480
rect 45020 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48516 354 48544 16546
rect 48976 3262 49004 246298
rect 49712 16574 49740 286282
rect 49712 16546 50200 16574
rect 48964 3256 49016 3262
rect 48964 3198 49016 3204
rect 50172 480 50200 16546
rect 50356 3738 50384 308586
rect 67640 307080 67692 307086
rect 67640 307022 67692 307028
rect 63500 289128 63552 289134
rect 63500 289070 63552 289076
rect 52460 287700 52512 287706
rect 52460 287642 52512 287648
rect 51080 258936 51132 258942
rect 51080 258878 51132 258884
rect 50344 3732 50396 3738
rect 50344 3674 50396 3680
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51092 354 51120 258878
rect 52472 3602 52500 287642
rect 62120 278044 62172 278050
rect 62120 277986 62172 277992
rect 61384 276684 61436 276690
rect 61384 276626 61436 276632
rect 57244 275324 57296 275330
rect 57244 275266 57296 275272
rect 52552 268388 52604 268394
rect 52552 268330 52604 268336
rect 52460 3596 52512 3602
rect 52460 3538 52512 3544
rect 52564 480 52592 268330
rect 56600 254720 56652 254726
rect 56600 254662 56652 254668
rect 53840 246424 53892 246430
rect 53840 246366 53892 246372
rect 53852 16574 53880 246366
rect 56612 16574 56640 254662
rect 53852 16546 54984 16574
rect 56612 16546 56824 16574
rect 53380 3596 53432 3602
rect 53380 3538 53432 3544
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53392 354 53420 3538
rect 54956 480 54984 16546
rect 56048 3392 56100 3398
rect 56048 3334 56100 3340
rect 56060 480 56088 3334
rect 53718 354 53830 480
rect 53392 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 57256 3398 57284 275266
rect 60740 260228 60792 260234
rect 60740 260170 60792 260176
rect 57980 246492 58032 246498
rect 57980 246434 58032 246440
rect 57992 16574 58020 246434
rect 60752 16574 60780 260170
rect 57992 16546 58480 16574
rect 60752 16546 61332 16574
rect 57244 3392 57296 3398
rect 57244 3334 57296 3340
rect 58452 480 58480 16546
rect 60832 3664 60884 3670
rect 60832 3606 60884 3612
rect 59636 3392 59688 3398
rect 59636 3334 59688 3340
rect 59648 480 59676 3334
rect 60844 480 60872 3606
rect 61304 490 61332 16546
rect 61396 3398 61424 276626
rect 62132 16574 62160 277986
rect 63512 16574 63540 289070
rect 66260 280900 66312 280906
rect 66260 280842 66312 280848
rect 64880 267096 64932 267102
rect 64880 267038 64932 267044
rect 64892 16574 64920 267038
rect 66272 16574 66300 280842
rect 62132 16546 63264 16574
rect 63512 16546 64368 16574
rect 64892 16546 65104 16574
rect 66272 16546 66760 16574
rect 61384 3392 61436 3398
rect 61384 3334 61436 3340
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61304 462 61700 490
rect 63236 480 63264 16546
rect 64340 480 64368 16546
rect 61672 354 61700 462
rect 61998 354 62110 480
rect 61672 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66732 480 66760 16546
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 307022
rect 68296 3466 68324 308654
rect 75182 308544 75238 308553
rect 75182 308479 75238 308488
rect 74540 290556 74592 290562
rect 74540 290498 74592 290504
rect 70400 290488 70452 290494
rect 70400 290430 70452 290436
rect 69020 282192 69072 282198
rect 69020 282134 69072 282140
rect 69032 3466 69060 282134
rect 69112 247784 69164 247790
rect 69112 247726 69164 247732
rect 68284 3460 68336 3466
rect 68284 3402 68336 3408
rect 69020 3460 69072 3466
rect 69020 3402 69072 3408
rect 69124 480 69152 247726
rect 70412 16574 70440 290430
rect 73160 283688 73212 283694
rect 73160 283630 73212 283636
rect 71780 250572 71832 250578
rect 71780 250514 71832 250520
rect 71792 16574 71820 250514
rect 73172 16574 73200 283630
rect 74552 16574 74580 290498
rect 70412 16546 71544 16574
rect 71792 16546 72648 16574
rect 73172 16546 73384 16574
rect 74552 16546 75040 16574
rect 69940 3460 69992 3466
rect 69940 3402 69992 3408
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69952 354 69980 3402
rect 71516 480 71544 16546
rect 72620 480 72648 16546
rect 70278 354 70390 480
rect 69952 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 16546
rect 75012 480 75040 16546
rect 75196 3534 75224 308479
rect 124220 294636 124272 294642
rect 124220 294578 124272 294584
rect 117320 293412 117372 293418
rect 117320 293354 117372 293360
rect 110420 293344 110472 293350
rect 110420 293286 110472 293292
rect 102140 293276 102192 293282
rect 102140 293218 102192 293224
rect 92480 291984 92532 291990
rect 92480 291926 92532 291932
rect 88340 291916 88392 291922
rect 88340 291858 88392 291864
rect 85580 291848 85632 291854
rect 85580 291790 85632 291796
rect 77300 290624 77352 290630
rect 77300 290566 77352 290572
rect 75920 250640 75972 250646
rect 75920 250582 75972 250588
rect 75184 3528 75236 3534
rect 75184 3470 75236 3476
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 250582
rect 77312 3534 77340 290566
rect 77392 285048 77444 285054
rect 77392 284990 77444 284996
rect 77300 3528 77352 3534
rect 77300 3470 77352 3476
rect 77404 480 77432 284990
rect 82820 269884 82872 269890
rect 82820 269826 82872 269832
rect 79324 254788 79376 254794
rect 79324 254730 79376 254736
rect 78680 250708 78732 250714
rect 78680 250650 78732 250656
rect 78692 16574 78720 250650
rect 78692 16546 79272 16574
rect 78220 3528 78272 3534
rect 78220 3470 78272 3476
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78232 354 78260 3470
rect 78558 354 78670 480
rect 78232 326 78670 354
rect 79244 354 79272 16546
rect 79336 3670 79364 254730
rect 80060 253428 80112 253434
rect 80060 253370 80112 253376
rect 80072 16574 80100 253370
rect 82832 16574 82860 269826
rect 84200 253496 84252 253502
rect 84200 253438 84252 253444
rect 80072 16546 80928 16574
rect 82832 16546 83320 16574
rect 79324 3664 79376 3670
rect 79324 3606 79376 3612
rect 80900 480 80928 16546
rect 82084 3528 82136 3534
rect 82084 3470 82136 3476
rect 82096 480 82124 3470
rect 83292 480 83320 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84212 354 84240 253438
rect 85592 6914 85620 291790
rect 86960 285116 87012 285122
rect 86960 285058 87012 285064
rect 85672 271244 85724 271250
rect 85672 271186 85724 271192
rect 85684 16574 85712 271186
rect 86972 16574 87000 285058
rect 88352 16574 88380 291858
rect 91100 286408 91152 286414
rect 91100 286350 91152 286356
rect 89720 279540 89772 279546
rect 89720 279482 89772 279488
rect 89732 16574 89760 279482
rect 91112 16574 91140 286350
rect 85684 16546 86448 16574
rect 86972 16546 87552 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 85592 6886 85712 6914
rect 85684 480 85712 6886
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86420 354 86448 16546
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 87524 354 87552 16546
rect 89180 480 89208 16546
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 291926
rect 98000 286476 98052 286482
rect 98000 286418 98052 286424
rect 93860 285184 93912 285190
rect 93860 285126 93912 285132
rect 93872 3466 93900 285126
rect 96620 282328 96672 282334
rect 96620 282270 96672 282276
rect 93952 282260 94004 282266
rect 93952 282202 94004 282208
rect 93860 3460 93912 3466
rect 93860 3402 93912 3408
rect 93964 480 93992 282202
rect 96632 16574 96660 282270
rect 98012 16574 98040 286418
rect 100760 283756 100812 283762
rect 100760 283698 100812 283704
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 96252 3664 96304 3670
rect 96252 3606 96304 3612
rect 94780 3460 94832 3466
rect 94780 3402 94832 3408
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94792 354 94820 3402
rect 96264 480 96292 3606
rect 97460 480 97488 16546
rect 95118 354 95230 480
rect 94792 326 95230 354
rect 95118 -960 95230 326
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99840 3392 99892 3398
rect 99840 3334 99892 3340
rect 99852 480 99880 3334
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 283698
rect 102152 3466 102180 293218
rect 104164 290692 104216 290698
rect 104164 290634 104216 290640
rect 102232 286544 102284 286550
rect 102232 286486 102284 286492
rect 102140 3460 102192 3466
rect 102140 3402 102192 3408
rect 102244 480 102272 286486
rect 103520 282396 103572 282402
rect 103520 282338 103572 282344
rect 103532 16574 103560 282338
rect 103532 16546 104112 16574
rect 103336 3460 103388 3466
rect 103336 3402 103388 3408
rect 103348 480 103376 3402
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 104176 3534 104204 290634
rect 109040 287836 109092 287842
rect 109040 287778 109092 287784
rect 104900 287768 104952 287774
rect 104900 287710 104952 287716
rect 104912 16574 104940 287710
rect 107660 283824 107712 283830
rect 107660 283766 107712 283772
rect 107672 16574 107700 283766
rect 104912 16546 105768 16574
rect 107672 16546 108160 16574
rect 104164 3528 104216 3534
rect 104164 3470 104216 3476
rect 105740 480 105768 16546
rect 106924 3528 106976 3534
rect 106924 3470 106976 3476
rect 106936 480 106964 3470
rect 108132 480 108160 16546
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109052 354 109080 287778
rect 110432 6914 110460 293286
rect 112444 292052 112496 292058
rect 112444 291994 112496 292000
rect 111800 287904 111852 287910
rect 111800 287846 111852 287852
rect 110512 283892 110564 283898
rect 110512 283834 110564 283840
rect 110524 16574 110552 283834
rect 111812 16574 111840 287846
rect 110524 16546 111656 16574
rect 111812 16546 112392 16574
rect 110432 6886 110552 6914
rect 110524 480 110552 6886
rect 111628 480 111656 16546
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 112456 3670 112484 291994
rect 115940 289196 115992 289202
rect 115940 289138 115992 289144
rect 114560 285252 114612 285258
rect 114560 285194 114612 285200
rect 114572 16574 114600 285194
rect 115952 16574 115980 289138
rect 116584 254856 116636 254862
rect 116584 254798 116636 254804
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 112444 3664 112496 3670
rect 112444 3606 112496 3612
rect 114008 3664 114060 3670
rect 114008 3606 114060 3612
rect 114020 480 114048 3606
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 116596 3602 116624 254798
rect 116584 3596 116636 3602
rect 116584 3538 116636 3544
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 293354
rect 122840 289332 122892 289338
rect 122840 289274 122892 289280
rect 118700 289264 118752 289270
rect 118700 289206 118752 289212
rect 118712 3602 118740 289206
rect 121460 252136 121512 252142
rect 121460 252078 121512 252084
rect 118792 252068 118844 252074
rect 118792 252010 118844 252016
rect 118700 3596 118752 3602
rect 118700 3538 118752 3544
rect 118804 480 118832 252010
rect 121472 16574 121500 252078
rect 122852 16574 122880 289274
rect 124232 16574 124260 294578
rect 160100 282464 160152 282470
rect 160100 282406 160152 282412
rect 155960 281036 156012 281042
rect 155960 280978 156012 280984
rect 151820 280968 151872 280974
rect 151820 280910 151872 280916
rect 149060 279608 149112 279614
rect 149060 279550 149112 279556
rect 144920 278112 144972 278118
rect 144920 278054 144972 278060
rect 142160 276752 142212 276758
rect 142160 276694 142212 276700
rect 138020 274032 138072 274038
rect 138020 273974 138072 273980
rect 131120 272604 131172 272610
rect 131120 272546 131172 272552
rect 126980 264308 127032 264314
rect 126980 264250 127032 264256
rect 125600 260296 125652 260302
rect 125600 260238 125652 260244
rect 121472 16546 122328 16574
rect 122852 16546 123064 16574
rect 124232 16546 124720 16574
rect 119896 3596 119948 3602
rect 119896 3538 119948 3544
rect 121092 3596 121144 3602
rect 121092 3538 121144 3544
rect 119908 480 119936 3538
rect 121104 480 121132 3538
rect 122300 480 122328 16546
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124692 480 124720 16546
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125612 354 125640 260238
rect 126992 480 127020 264250
rect 128360 261588 128412 261594
rect 128360 261530 128412 261536
rect 127072 247852 127124 247858
rect 127072 247794 127124 247800
rect 127084 16574 127112 247794
rect 128372 16574 128400 261530
rect 129740 246560 129792 246566
rect 129740 246502 129792 246508
rect 129752 16574 129780 246502
rect 131132 16574 131160 272546
rect 136640 268456 136692 268462
rect 136640 268398 136692 268404
rect 133880 265736 133932 265742
rect 133880 265678 133932 265684
rect 132500 245132 132552 245138
rect 132500 245074 132552 245080
rect 132512 16574 132540 245074
rect 127084 16546 128216 16574
rect 128372 16546 128952 16574
rect 129752 16546 130608 16574
rect 131132 16546 131344 16574
rect 132512 16546 133000 16574
rect 128188 480 128216 16546
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 16546
rect 130580 480 130608 16546
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 132972 480 133000 16546
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 133892 354 133920 265678
rect 135260 249144 135312 249150
rect 135260 249086 135312 249092
rect 135272 480 135300 249086
rect 135352 245200 135404 245206
rect 135352 245142 135404 245148
rect 135364 16574 135392 245142
rect 136652 16574 136680 268398
rect 138032 16574 138060 273974
rect 140780 269952 140832 269958
rect 140780 269894 140832 269900
rect 139400 262948 139452 262954
rect 139400 262890 139452 262896
rect 139412 16574 139440 262890
rect 140792 16574 140820 269894
rect 135364 16546 136496 16574
rect 136652 16546 137232 16574
rect 138032 16546 138888 16574
rect 139412 16546 139624 16574
rect 140792 16546 141280 16574
rect 136468 480 136496 16546
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 16546
rect 138860 480 138888 16546
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 139596 354 139624 16546
rect 141252 480 141280 16546
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142172 354 142200 276694
rect 143540 271312 143592 271318
rect 143540 271254 143592 271260
rect 143552 11762 143580 271254
rect 143632 264376 143684 264382
rect 143632 264318 143684 264324
rect 143540 11756 143592 11762
rect 143540 11698 143592 11704
rect 143644 6914 143672 264318
rect 144932 16574 144960 278054
rect 146300 265804 146352 265810
rect 146300 265746 146352 265752
rect 146312 16574 146340 265746
rect 147680 247920 147732 247926
rect 147680 247862 147732 247868
rect 147692 16574 147720 247862
rect 149072 16574 149100 279550
rect 150440 267164 150492 267170
rect 150440 267106 150492 267112
rect 150452 16574 150480 267106
rect 144932 16546 145512 16574
rect 146312 16546 147168 16574
rect 147692 16546 147904 16574
rect 149072 16546 149560 16574
rect 150452 16546 150664 16574
rect 144736 11756 144788 11762
rect 144736 11698 144788 11704
rect 143552 6886 143672 6914
rect 143552 480 143580 6886
rect 144748 480 144776 11698
rect 142406 354 142518 480
rect 142172 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 147140 480 147168 16546
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 149532 480 149560 16546
rect 150636 480 150664 16546
rect 151832 9674 151860 280910
rect 154580 272672 154632 272678
rect 154580 272614 154632 272620
rect 153200 267232 153252 267238
rect 153200 267174 153252 267180
rect 151912 247988 151964 247994
rect 151912 247930 151964 247936
rect 151740 9654 151860 9674
rect 151728 9648 151860 9654
rect 151780 9646 151860 9648
rect 151728 9590 151780 9596
rect 151924 6914 151952 247930
rect 153212 16574 153240 267174
rect 154592 16574 154620 272614
rect 155972 16574 156000 280978
rect 158720 274100 158772 274106
rect 158720 274042 158772 274048
rect 157340 268524 157392 268530
rect 157340 268466 157392 268472
rect 157352 16574 157380 268466
rect 158732 16574 158760 274042
rect 153212 16546 153792 16574
rect 154592 16546 155448 16574
rect 155972 16546 156184 16574
rect 157352 16546 157840 16574
rect 158732 16546 158944 16574
rect 153016 9648 153068 9654
rect 153016 9590 153068 9596
rect 151832 6886 151952 6914
rect 151832 480 151860 6886
rect 153028 480 153056 9590
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 16546
rect 155420 480 155448 16546
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156156 354 156184 16546
rect 157812 480 157840 16546
rect 158916 480 158944 16546
rect 160112 480 160140 282406
rect 176660 276956 176712 276962
rect 176660 276898 176712 276904
rect 173900 276888 173952 276894
rect 173900 276830 173952 276836
rect 169760 276820 169812 276826
rect 169760 276762 169812 276768
rect 167000 275460 167052 275466
rect 167000 275402 167052 275408
rect 162860 275392 162912 275398
rect 162860 275334 162912 275340
rect 161480 268592 161532 268598
rect 161480 268534 161532 268540
rect 160192 260364 160244 260370
rect 160192 260306 160244 260312
rect 160204 16574 160232 260306
rect 161492 16574 161520 268534
rect 162872 16574 162900 275334
rect 165620 268660 165672 268666
rect 165620 268602 165672 268608
rect 164240 261656 164292 261662
rect 164240 261598 164292 261604
rect 164252 16574 164280 261598
rect 165632 16574 165660 268602
rect 167012 16574 167040 275402
rect 168380 270020 168432 270026
rect 168380 269962 168432 269968
rect 160204 16546 161336 16574
rect 161492 16546 162072 16574
rect 162872 16546 163728 16574
rect 164252 16546 164464 16574
rect 165632 16546 166120 16574
rect 167012 16546 167224 16574
rect 161308 480 161336 16546
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 354 162072 16546
rect 163700 480 163728 16546
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164436 354 164464 16546
rect 166092 480 166120 16546
rect 167196 480 167224 16546
rect 168392 11762 168420 269962
rect 168472 261724 168524 261730
rect 168472 261666 168524 261672
rect 168380 11756 168432 11762
rect 168380 11698 168432 11704
rect 168484 6914 168512 261666
rect 169772 16574 169800 276762
rect 172520 270088 172572 270094
rect 172520 270030 172572 270036
rect 171140 261792 171192 261798
rect 171140 261734 171192 261740
rect 171152 16574 171180 261734
rect 172532 16574 172560 270030
rect 169772 16546 170352 16574
rect 171152 16546 172008 16574
rect 172532 16546 172744 16574
rect 169576 11756 169628 11762
rect 169576 11698 169628 11704
rect 168392 6886 168512 6914
rect 168392 480 168420 6886
rect 169588 480 169616 11698
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170324 354 170352 16546
rect 171980 480 172008 16546
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173912 354 173940 276830
rect 175280 263152 175332 263158
rect 175280 263094 175332 263100
rect 174544 250776 174596 250782
rect 174544 250718 174596 250724
rect 174556 3466 174584 250718
rect 175292 16574 175320 263094
rect 175292 16546 175504 16574
rect 174544 3460 174596 3466
rect 174544 3402 174596 3408
rect 175476 480 175504 16546
rect 176672 3534 176700 276898
rect 176660 3528 176712 3534
rect 176660 3470 176712 3476
rect 177856 3528 177908 3534
rect 177856 3470 177908 3476
rect 176660 3052 176712 3058
rect 176660 2994 176712 3000
rect 176672 480 176700 2994
rect 177868 480 177896 3470
rect 178696 3466 178724 308722
rect 179420 271380 179472 271386
rect 179420 271322 179472 271328
rect 178776 270156 178828 270162
rect 178776 270098 178828 270104
rect 178684 3460 178736 3466
rect 178684 3402 178736 3408
rect 178788 3058 178816 270098
rect 179432 16574 179460 271322
rect 180076 137970 180104 443090
rect 189724 308984 189776 308990
rect 189724 308926 189776 308932
rect 182824 308916 182876 308922
rect 182824 308858 182876 308864
rect 180800 278180 180852 278186
rect 180800 278122 180852 278128
rect 180064 137964 180116 137970
rect 180064 137906 180116 137912
rect 180812 16574 180840 278122
rect 182180 263016 182232 263022
rect 182180 262958 182232 262964
rect 179432 16546 180288 16574
rect 180812 16546 181024 16574
rect 179052 3460 179104 3466
rect 179052 3402 179104 3408
rect 178776 3052 178828 3058
rect 178776 2994 178828 3000
rect 179064 480 179092 3402
rect 180260 480 180288 16546
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 173134 -960 173246 326
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 182192 354 182220 262958
rect 182836 3670 182864 308858
rect 189080 307148 189132 307154
rect 189080 307090 189132 307096
rect 187700 278316 187752 278322
rect 187700 278258 187752 278264
rect 184940 278248 184992 278254
rect 184940 278190 184992 278196
rect 183560 271448 183612 271454
rect 183560 271390 183612 271396
rect 183572 16574 183600 271390
rect 183572 16546 183784 16574
rect 182824 3664 182876 3670
rect 182824 3606 182876 3612
rect 183756 480 183784 16546
rect 184952 480 184980 278190
rect 185032 263084 185084 263090
rect 185032 263026 185084 263032
rect 185044 16574 185072 263026
rect 187712 16574 187740 278258
rect 188344 271516 188396 271522
rect 188344 271458 188396 271464
rect 185044 16546 186176 16574
rect 187712 16546 188292 16574
rect 186148 480 186176 16546
rect 187332 3596 187384 3602
rect 187332 3538 187384 3544
rect 187344 480 187372 3538
rect 188264 3482 188292 16546
rect 188356 3602 188384 271458
rect 189092 16574 189120 307090
rect 189092 16546 189304 16574
rect 188344 3596 188396 3602
rect 188344 3538 188396 3544
rect 188264 3454 188568 3482
rect 188540 480 188568 3454
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189276 354 189304 16546
rect 189736 3670 189764 308926
rect 202880 307216 202932 307222
rect 202880 307158 202932 307164
rect 201500 281104 201552 281110
rect 201500 281046 201552 281052
rect 198740 279812 198792 279818
rect 198740 279754 198792 279760
rect 196624 279744 196676 279750
rect 196624 279686 196676 279692
rect 191840 279676 191892 279682
rect 191840 279618 191892 279624
rect 191852 16574 191880 279618
rect 193220 272740 193272 272746
rect 193220 272682 193272 272688
rect 192484 246628 192536 246634
rect 192484 246570 192536 246576
rect 191852 16546 192064 16574
rect 189724 3664 189776 3670
rect 189724 3606 189776 3612
rect 190828 3528 190880 3534
rect 190828 3470 190880 3476
rect 190840 480 190868 3470
rect 192036 480 192064 16546
rect 192496 3534 192524 246570
rect 193232 3602 193260 272682
rect 195980 264512 196032 264518
rect 195980 264454 196032 264460
rect 193312 264444 193364 264450
rect 193312 264386 193364 264392
rect 193220 3596 193272 3602
rect 193220 3538 193272 3544
rect 192484 3528 192536 3534
rect 193324 3482 193352 264386
rect 195992 16574 196020 264454
rect 195992 16546 196572 16574
rect 194416 3596 194468 3602
rect 194416 3538 194468 3544
rect 195612 3596 195664 3602
rect 195612 3538 195664 3544
rect 192484 3470 192536 3476
rect 193232 3454 193352 3482
rect 193232 480 193260 3454
rect 194428 480 194456 3538
rect 195624 480 195652 3538
rect 196544 3482 196572 16546
rect 196636 3602 196664 279686
rect 197360 272808 197412 272814
rect 197360 272750 197412 272756
rect 197372 16574 197400 272750
rect 197372 16546 197952 16574
rect 196624 3596 196676 3602
rect 196624 3538 196676 3544
rect 196544 3454 196848 3482
rect 196820 480 196848 3454
rect 197924 480 197952 16546
rect 189694 354 189806 480
rect 189276 326 189806 354
rect 189694 -960 189806 326
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 279754
rect 201512 11762 201540 281046
rect 201592 272876 201644 272882
rect 201592 272818 201644 272824
rect 201500 11756 201552 11762
rect 201500 11698 201552 11704
rect 201604 6914 201632 272818
rect 202892 16574 202920 307158
rect 206284 274168 206336 274174
rect 206284 274110 206336 274116
rect 205640 249212 205692 249218
rect 205640 249154 205692 249160
rect 205652 16574 205680 249154
rect 202892 16546 203472 16574
rect 205652 16546 206232 16574
rect 202696 11756 202748 11762
rect 202696 11698 202748 11704
rect 201512 6886 201632 6914
rect 200302 3360 200358 3369
rect 200302 3295 200358 3304
rect 200316 480 200344 3295
rect 201512 480 201540 6886
rect 202708 480 202736 11698
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203444 354 203472 16546
rect 205088 3528 205140 3534
rect 205088 3470 205140 3476
rect 205100 480 205128 3470
rect 206204 480 206232 16546
rect 206296 3534 206324 274110
rect 209780 265872 209832 265878
rect 209780 265814 209832 265820
rect 207020 264580 207072 264586
rect 207020 264522 207072 264528
rect 206284 3528 206336 3534
rect 206284 3470 206336 3476
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 264522
rect 207664 261860 207716 261866
rect 207664 261802 207716 261808
rect 207676 3466 207704 261802
rect 209792 9674 209820 265814
rect 209872 249280 209924 249286
rect 209872 249222 209924 249228
rect 209700 9654 209820 9674
rect 209688 9648 209820 9654
rect 209740 9646 209820 9648
rect 209688 9590 209740 9596
rect 209884 6914 209912 249222
rect 210436 215286 210464 446762
rect 217796 446486 217824 487999
rect 217888 457502 217916 516831
rect 217876 457496 217928 457502
rect 217876 457438 217928 457444
rect 217980 446894 218008 565082
rect 218072 454986 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 234632 565146 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 700330 267688 703520
rect 283852 700398 283880 703520
rect 300136 700466 300164 703520
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 300124 700460 300176 700466
rect 300124 700402 300176 700408
rect 283840 700392 283892 700398
rect 283840 700334 283892 700340
rect 267648 700324 267700 700330
rect 267648 700266 267700 700272
rect 331232 565146 331260 702986
rect 348804 700534 348832 703520
rect 348792 700528 348844 700534
rect 348792 700470 348844 700476
rect 358912 700528 358964 700534
rect 358912 700470 358964 700476
rect 357532 700460 357584 700466
rect 357532 700402 357584 700408
rect 357440 700324 357492 700330
rect 357440 700266 357492 700272
rect 234620 565140 234672 565146
rect 234620 565082 234672 565088
rect 331220 565140 331272 565146
rect 331220 565082 331272 565088
rect 219070 512816 219126 512825
rect 219070 512751 219126 512760
rect 219084 475454 219112 512751
rect 219162 511048 219218 511057
rect 219162 510983 219218 510992
rect 219072 475448 219124 475454
rect 219072 475390 219124 475396
rect 219176 472666 219204 510983
rect 219346 509960 219402 509969
rect 219346 509895 219402 509904
rect 219254 508192 219310 508201
rect 219254 508127 219310 508136
rect 219164 472660 219216 472666
rect 219164 472602 219216 472608
rect 219268 456210 219296 508127
rect 219256 456204 219308 456210
rect 219256 456146 219308 456152
rect 219360 456142 219388 509895
rect 220084 478916 220136 478922
rect 220084 478858 220136 478864
rect 219348 456136 219400 456142
rect 219348 456078 219400 456084
rect 218060 454980 218112 454986
rect 218060 454922 218112 454928
rect 217968 446888 218020 446894
rect 217968 446830 218020 446836
rect 220096 446554 220124 478858
rect 311900 478236 311952 478242
rect 311900 478178 311952 478184
rect 264978 477320 265034 477329
rect 264978 477255 265034 477264
rect 268014 477320 268070 477329
rect 268014 477255 268070 477264
rect 255318 477184 255374 477193
rect 255318 477119 255374 477128
rect 252558 476776 252614 476785
rect 252558 476711 252614 476720
rect 252572 476678 252600 476711
rect 241612 476672 241664 476678
rect 252560 476672 252612 476678
rect 241612 476614 241664 476620
rect 244278 476640 244334 476649
rect 238760 476536 238812 476542
rect 238760 476478 238812 476484
rect 236092 476468 236144 476474
rect 236092 476410 236144 476416
rect 234712 476332 234764 476338
rect 234712 476274 234764 476280
rect 234620 476128 234672 476134
rect 234620 476070 234672 476076
rect 234252 450696 234304 450702
rect 234252 450638 234304 450644
rect 220084 446548 220136 446554
rect 220084 446490 220136 446496
rect 232780 446548 232832 446554
rect 232780 446490 232832 446496
rect 217784 446480 217836 446486
rect 217784 446422 217836 446428
rect 232320 446140 232372 446146
rect 232320 446082 232372 446088
rect 231124 446004 231176 446010
rect 231124 445946 231176 445952
rect 228364 444848 228416 444854
rect 228364 444790 228416 444796
rect 218428 444780 218480 444786
rect 218428 444722 218480 444728
rect 215208 309120 215260 309126
rect 215208 309062 215260 309068
rect 213828 308848 213880 308854
rect 213828 308790 213880 308796
rect 213736 305924 213788 305930
rect 213736 305866 213788 305872
rect 212448 303612 212500 303618
rect 212448 303554 212500 303560
rect 211068 303272 211120 303278
rect 211068 303214 211120 303220
rect 210608 302932 210660 302938
rect 210608 302874 210660 302880
rect 210516 300348 210568 300354
rect 210516 300290 210568 300296
rect 210424 215280 210476 215286
rect 210424 215222 210476 215228
rect 210528 193118 210556 300290
rect 210516 193112 210568 193118
rect 210516 193054 210568 193060
rect 210620 189038 210648 302874
rect 210976 300552 211028 300558
rect 210976 300494 211028 300500
rect 210884 300484 210936 300490
rect 210884 300426 210936 300432
rect 210700 300280 210752 300286
rect 210700 300222 210752 300228
rect 210608 189032 210660 189038
rect 210608 188974 210660 188980
rect 210712 155242 210740 300222
rect 210792 300212 210844 300218
rect 210792 300154 210844 300160
rect 210804 155378 210832 300154
rect 210896 155553 210924 300426
rect 210882 155544 210938 155553
rect 210882 155479 210938 155488
rect 210988 155417 211016 300494
rect 211080 155825 211108 303214
rect 212356 303204 212408 303210
rect 212356 303146 212408 303152
rect 212078 303104 212134 303113
rect 212078 303039 212134 303048
rect 211896 303000 211948 303006
rect 211896 302942 211948 302948
rect 211804 274304 211856 274310
rect 211804 274246 211856 274252
rect 211160 274236 211212 274242
rect 211160 274178 211212 274184
rect 211066 155816 211122 155825
rect 211066 155751 211122 155760
rect 210974 155408 211030 155417
rect 210792 155372 210844 155378
rect 210974 155343 211030 155352
rect 210792 155314 210844 155320
rect 210700 155236 210752 155242
rect 210700 155178 210752 155184
rect 211172 16574 211200 274178
rect 211172 16546 211752 16574
rect 210976 9648 211028 9654
rect 210976 9590 211028 9596
rect 209792 6886 209912 6914
rect 208584 3596 208636 3602
rect 208584 3538 208636 3544
rect 207664 3460 207716 3466
rect 207664 3402 207716 3408
rect 208596 480 208624 3538
rect 209792 480 209820 6886
rect 210988 480 211016 9590
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 16546
rect 211816 3602 211844 274246
rect 211908 158778 211936 302942
rect 211986 302832 212042 302841
rect 211986 302767 212042 302776
rect 211896 158772 211948 158778
rect 211896 158714 211948 158720
rect 212000 158506 212028 302767
rect 211988 158500 212040 158506
rect 211988 158442 212040 158448
rect 212092 157962 212120 303039
rect 212172 300688 212224 300694
rect 212172 300630 212224 300636
rect 212080 157956 212132 157962
rect 212080 157898 212132 157904
rect 212184 155310 212212 300630
rect 212264 300416 212316 300422
rect 212264 300358 212316 300364
rect 212172 155304 212224 155310
rect 212172 155246 212224 155252
rect 212276 152590 212304 300358
rect 212368 155689 212396 303146
rect 212354 155680 212410 155689
rect 212354 155615 212410 155624
rect 212264 152584 212316 152590
rect 212264 152526 212316 152532
rect 211804 3596 211856 3602
rect 211804 3538 211856 3544
rect 212460 3398 212488 303554
rect 213552 303544 213604 303550
rect 213552 303486 213604 303492
rect 213092 303476 213144 303482
rect 213092 303418 213144 303424
rect 213000 245268 213052 245274
rect 213000 245210 213052 245216
rect 213012 169590 213040 245210
rect 213000 169584 213052 169590
rect 213000 169526 213052 169532
rect 213104 159662 213132 303418
rect 213368 303136 213420 303142
rect 213368 303078 213420 303084
rect 213274 302968 213330 302977
rect 213274 302903 213330 302912
rect 213184 300620 213236 300626
rect 213184 300562 213236 300568
rect 213092 159656 213144 159662
rect 213092 159598 213144 159604
rect 213196 155281 213224 300562
rect 213288 158370 213316 302903
rect 213380 158710 213408 303078
rect 213460 300144 213512 300150
rect 213460 300086 213512 300092
rect 213368 158704 213420 158710
rect 213368 158646 213420 158652
rect 213276 158364 213328 158370
rect 213276 158306 213328 158312
rect 213182 155272 213238 155281
rect 213182 155207 213238 155216
rect 213472 152522 213500 300086
rect 213564 155961 213592 303486
rect 213644 303340 213696 303346
rect 213644 303282 213696 303288
rect 213550 155952 213606 155961
rect 213550 155887 213606 155896
rect 213460 152516 213512 152522
rect 213460 152458 213512 152464
rect 213656 4146 213684 303282
rect 213644 4140 213696 4146
rect 213644 4082 213696 4088
rect 213748 4078 213776 305866
rect 213736 4072 213788 4078
rect 213736 4014 213788 4020
rect 213840 3670 213868 308790
rect 214564 306196 214616 306202
rect 214564 306138 214616 306144
rect 214472 305856 214524 305862
rect 214472 305798 214524 305804
rect 214380 300756 214432 300762
rect 214380 300698 214432 300704
rect 214392 195294 214420 300698
rect 214380 195288 214432 195294
rect 214380 195230 214432 195236
rect 214484 159526 214512 305798
rect 214472 159520 214524 159526
rect 214472 159462 214524 159468
rect 214576 158642 214604 306138
rect 215024 306060 215076 306066
rect 215024 306002 215076 306008
rect 214656 305992 214708 305998
rect 214656 305934 214708 305940
rect 214564 158636 214616 158642
rect 214564 158578 214616 158584
rect 214668 158234 214696 305934
rect 214748 305720 214800 305726
rect 214748 305662 214800 305668
rect 214656 158228 214708 158234
rect 214656 158170 214708 158176
rect 214760 155106 214788 305662
rect 214930 300112 214986 300121
rect 214930 300047 214986 300056
rect 214840 245336 214892 245342
rect 214840 245278 214892 245284
rect 214748 155100 214800 155106
rect 214748 155042 214800 155048
rect 213828 3664 213880 3670
rect 213828 3606 213880 3612
rect 213366 3496 213422 3505
rect 213366 3431 213422 3440
rect 214470 3496 214526 3505
rect 214852 3466 214880 245278
rect 214944 3942 214972 300047
rect 214932 3936 214984 3942
rect 214932 3878 214984 3884
rect 214470 3431 214526 3440
rect 214840 3460 214892 3466
rect 212448 3392 212500 3398
rect 212448 3334 212500 3340
rect 213380 480 213408 3431
rect 214484 480 214512 3431
rect 214840 3402 214892 3408
rect 215036 3262 215064 306002
rect 215116 305584 215168 305590
rect 215116 305526 215168 305532
rect 215024 3256 215076 3262
rect 215128 3233 215156 305526
rect 215220 3330 215248 309062
rect 216496 309052 216548 309058
rect 216496 308994 216548 309000
rect 216404 306332 216456 306338
rect 216404 306274 216456 306280
rect 216312 306128 216364 306134
rect 216312 306070 216364 306076
rect 216128 305788 216180 305794
rect 216128 305730 216180 305736
rect 215944 302796 215996 302802
rect 215944 302738 215996 302744
rect 215852 300076 215904 300082
rect 215852 300018 215904 300024
rect 215760 243568 215812 243574
rect 215760 243510 215812 243516
rect 215772 193186 215800 243510
rect 215760 193180 215812 193186
rect 215760 193122 215812 193128
rect 215864 189310 215892 300018
rect 215852 189304 215904 189310
rect 215852 189246 215904 189252
rect 215956 158166 215984 302738
rect 216036 300824 216088 300830
rect 216036 300766 216088 300772
rect 215944 158160 215996 158166
rect 215944 158102 215996 158108
rect 216048 155174 216076 300766
rect 216140 159390 216168 305730
rect 216220 305448 216272 305454
rect 216220 305390 216272 305396
rect 216128 159384 216180 159390
rect 216128 159326 216180 159332
rect 216232 157894 216260 305390
rect 216324 158098 216352 306070
rect 216416 158438 216444 306274
rect 216404 158432 216456 158438
rect 216404 158374 216456 158380
rect 216508 158302 216536 308994
rect 217692 305652 217744 305658
rect 217692 305594 217744 305600
rect 216588 305516 216640 305522
rect 216588 305458 216640 305464
rect 216496 158296 216548 158302
rect 216496 158238 216548 158244
rect 216312 158092 216364 158098
rect 216312 158034 216364 158040
rect 216220 157888 216272 157894
rect 216220 157830 216272 157836
rect 216036 155168 216088 155174
rect 216036 155110 216088 155116
rect 215666 3496 215722 3505
rect 215666 3431 215722 3440
rect 215208 3324 215260 3330
rect 215208 3266 215260 3272
rect 215024 3198 215076 3204
rect 215114 3224 215170 3233
rect 215114 3159 215170 3168
rect 215680 480 215708 3431
rect 216600 3097 216628 305458
rect 217416 304292 217468 304298
rect 217416 304234 217468 304240
rect 217048 301708 217100 301714
rect 217048 301650 217100 301656
rect 217060 193769 217088 301650
rect 217140 257372 217192 257378
rect 217140 257314 217192 257320
rect 217046 193760 217102 193769
rect 217046 193695 217102 193704
rect 216680 193112 216732 193118
rect 216680 193054 216732 193060
rect 216692 192817 216720 193054
rect 216678 192808 216734 192817
rect 216678 192743 216734 192752
rect 216680 189032 216732 189038
rect 216680 188974 216732 188980
rect 216692 188193 216720 188974
rect 216678 188184 216734 188193
rect 216678 188119 216734 188128
rect 217152 169969 217180 257314
rect 217232 243704 217284 243710
rect 217232 243646 217284 243652
rect 217138 169960 217194 169969
rect 217138 169895 217194 169904
rect 217244 155038 217272 243646
rect 217428 196897 217456 304234
rect 217508 302660 217560 302666
rect 217508 302602 217560 302608
rect 217414 196888 217470 196897
rect 217414 196823 217470 196832
rect 217520 195945 217548 302602
rect 217600 301776 217652 301782
rect 217600 301718 217652 301724
rect 217506 195936 217562 195945
rect 217506 195871 217562 195880
rect 217324 195288 217376 195294
rect 217324 195230 217376 195236
rect 217232 155032 217284 155038
rect 217232 154974 217284 154980
rect 217336 3874 217364 195230
rect 217416 193180 217468 193186
rect 217416 193122 217468 193128
rect 217324 3868 217376 3874
rect 217324 3810 217376 3816
rect 217428 3738 217456 193122
rect 217508 169584 217560 169590
rect 217508 169526 217560 169532
rect 217416 3732 217468 3738
rect 217416 3674 217468 3680
rect 217520 3534 217548 169526
rect 217612 168337 217640 301718
rect 217598 168328 217654 168337
rect 217598 168263 217654 168272
rect 217704 168065 217732 305594
rect 217968 303408 218020 303414
rect 217968 303350 218020 303356
rect 217876 302864 217928 302870
rect 217876 302806 217928 302812
rect 217784 300008 217836 300014
rect 217784 299950 217836 299956
rect 217690 168056 217746 168065
rect 217690 167991 217746 168000
rect 217796 159458 217824 299950
rect 217888 159594 217916 302806
rect 217876 159588 217928 159594
rect 217876 159530 217928 159536
rect 217784 159452 217836 159458
rect 217784 159394 217836 159400
rect 217980 156466 218008 303350
rect 218440 243409 218468 444722
rect 218980 308372 219032 308378
rect 218980 308314 219032 308320
rect 218888 308236 218940 308242
rect 218888 308178 218940 308184
rect 218704 306264 218756 306270
rect 218704 306206 218756 306212
rect 218612 296268 218664 296274
rect 218612 296210 218664 296216
rect 218520 294908 218572 294914
rect 218520 294850 218572 294856
rect 218426 243400 218482 243409
rect 218426 243335 218482 243344
rect 218532 189961 218560 294850
rect 218624 191049 218652 296210
rect 218610 191040 218666 191049
rect 218610 190975 218666 190984
rect 218518 189952 218574 189961
rect 218518 189887 218574 189896
rect 218612 189304 218664 189310
rect 218612 189246 218664 189252
rect 217968 156460 218020 156466
rect 217968 156402 218020 156408
rect 218624 152658 218652 189246
rect 218716 158030 218744 306206
rect 218796 302728 218848 302734
rect 218796 302670 218848 302676
rect 218704 158024 218756 158030
rect 218704 157966 218756 157972
rect 218808 155446 218836 302670
rect 218900 158545 218928 308178
rect 218992 158574 219020 308314
rect 219072 308304 219124 308310
rect 219072 308246 219124 308252
rect 218980 158568 219032 158574
rect 218886 158536 218942 158545
rect 218980 158510 219032 158516
rect 218886 158471 218942 158480
rect 219084 157826 219112 308246
rect 219348 299940 219400 299946
rect 219348 299882 219400 299888
rect 219164 243772 219216 243778
rect 219164 243714 219216 243720
rect 219072 157820 219124 157826
rect 219072 157762 219124 157768
rect 218796 155440 218848 155446
rect 218796 155382 218848 155388
rect 218612 152652 218664 152658
rect 218612 152594 218664 152600
rect 219176 3806 219204 243714
rect 219256 243636 219308 243642
rect 219256 243578 219308 243584
rect 219164 3800 219216 3806
rect 219164 3742 219216 3748
rect 218058 3632 218114 3641
rect 219268 3602 219296 243578
rect 219360 4010 219388 299882
rect 228376 267714 228404 444790
rect 228364 267708 228416 267714
rect 228364 267650 228416 267656
rect 231136 258806 231164 445946
rect 232228 445936 232280 445942
rect 232228 445878 232280 445884
rect 231216 444916 231268 444922
rect 231216 444858 231268 444864
rect 231228 358766 231256 444858
rect 232240 434042 232268 445878
rect 232228 434036 232280 434042
rect 232228 433978 232280 433984
rect 232332 412634 232360 446082
rect 232792 443972 232820 446490
rect 233516 446480 233568 446486
rect 233516 446422 233568 446428
rect 233528 443972 233556 446422
rect 233792 446072 233844 446078
rect 233792 446014 233844 446020
rect 233804 443970 233832 446014
rect 233884 445868 233936 445874
rect 233884 445810 233936 445816
rect 233792 443964 233844 443970
rect 233792 443906 233844 443912
rect 233896 443902 233924 445810
rect 234264 443972 234292 450638
rect 234632 443986 234660 476070
rect 234724 460934 234752 476274
rect 235906 476232 235962 476241
rect 235906 476167 235962 476176
rect 235920 476134 235948 476167
rect 235908 476128 235960 476134
rect 235908 476070 235960 476076
rect 236104 460934 236132 476410
rect 237378 476368 237434 476377
rect 237378 476303 237434 476312
rect 234724 460906 235488 460934
rect 236104 460906 236224 460934
rect 235460 443986 235488 460906
rect 236196 443986 236224 460906
rect 234632 443958 235106 443986
rect 235460 443958 235842 443986
rect 236196 443958 236670 443986
rect 237392 443972 237420 476303
rect 237470 476232 237526 476241
rect 237470 476167 237526 476176
rect 237484 460934 237512 476167
rect 237484 460906 237880 460934
rect 237852 443986 237880 460906
rect 238772 443986 238800 476478
rect 238852 476400 238904 476406
rect 238852 476342 238904 476348
rect 238864 460934 238892 476342
rect 241520 476264 241572 476270
rect 240138 476232 240194 476241
rect 240138 476167 240194 476176
rect 241426 476232 241482 476241
rect 241520 476206 241572 476212
rect 241426 476167 241482 476176
rect 238864 460906 239352 460934
rect 239324 443986 239352 460906
rect 240152 443986 240180 476167
rect 241440 476134 241468 476167
rect 241428 476128 241480 476134
rect 241428 476070 241480 476076
rect 240968 456204 241020 456210
rect 240968 456146 241020 456152
rect 240980 443986 241008 456146
rect 241532 443986 241560 476206
rect 241624 460934 241652 476614
rect 244278 476575 244334 476584
rect 247038 476640 247094 476649
rect 247038 476575 247094 476584
rect 249798 476640 249854 476649
rect 252560 476614 252612 476620
rect 249798 476575 249854 476584
rect 244292 476542 244320 476575
rect 244280 476536 244332 476542
rect 244280 476478 244332 476484
rect 247052 476474 247080 476575
rect 249812 476542 249840 476575
rect 249800 476536 249852 476542
rect 249800 476478 249852 476484
rect 252652 476536 252704 476542
rect 252652 476478 252704 476484
rect 247040 476468 247092 476474
rect 247040 476410 247092 476416
rect 251180 476468 251232 476474
rect 251180 476410 251232 476416
rect 242898 476368 242954 476377
rect 242898 476303 242900 476312
rect 242952 476303 242954 476312
rect 244278 476368 244334 476377
rect 244278 476303 244334 476312
rect 245752 476332 245804 476338
rect 242900 476274 242952 476280
rect 244292 476270 244320 476303
rect 245752 476274 245804 476280
rect 244280 476264 244332 476270
rect 242806 476232 242862 476241
rect 244280 476206 244332 476212
rect 245658 476232 245714 476241
rect 242806 476167 242808 476176
rect 242860 476167 242862 476176
rect 244924 476196 244976 476202
rect 242808 476138 242860 476144
rect 245658 476167 245714 476176
rect 244924 476138 244976 476144
rect 242900 476128 242952 476134
rect 242900 476070 242952 476076
rect 244280 476128 244332 476134
rect 244280 476070 244332 476076
rect 242912 460934 242940 476070
rect 241624 460906 242480 460934
rect 242912 460906 243216 460934
rect 242452 443986 242480 460906
rect 243188 443986 243216 460906
rect 244292 447302 244320 476070
rect 244936 460934 244964 476138
rect 245672 476134 245700 476167
rect 245660 476128 245712 476134
rect 245660 476070 245712 476076
rect 244936 460906 245056 460934
rect 244372 456136 244424 456142
rect 244372 456078 244424 456084
rect 244280 447296 244332 447302
rect 244280 447238 244332 447244
rect 237852 443958 238234 443986
rect 238772 443958 238970 443986
rect 239324 443958 239798 443986
rect 240152 443958 240534 443986
rect 240980 443958 241362 443986
rect 241532 443958 242098 443986
rect 242452 443958 242834 443986
rect 243188 443958 243662 443986
rect 244384 443972 244412 456078
rect 244924 447296 244976 447302
rect 244924 447238 244976 447244
rect 244936 443986 244964 447238
rect 245028 447098 245056 460906
rect 245016 447092 245068 447098
rect 245016 447034 245068 447040
rect 245764 443986 245792 476274
rect 248420 476264 248472 476270
rect 247222 476232 247278 476241
rect 248420 476206 248472 476212
rect 249798 476232 249854 476241
rect 247222 476167 247278 476176
rect 247132 472660 247184 472666
rect 247132 472602 247184 472608
rect 246764 447092 246816 447098
rect 246764 447034 246816 447040
rect 244936 443958 245226 443986
rect 245764 443958 245962 443986
rect 246776 443972 246804 447034
rect 247144 443986 247172 472602
rect 247236 460934 247264 476167
rect 248432 460934 248460 476206
rect 249798 476167 249854 476176
rect 251086 476232 251142 476241
rect 251086 476167 251142 476176
rect 247236 460906 248000 460934
rect 248432 460906 248736 460934
rect 247972 443986 248000 460906
rect 248708 443986 248736 460906
rect 249812 447302 249840 476167
rect 251100 476134 251128 476167
rect 251088 476128 251140 476134
rect 251088 476070 251140 476076
rect 249892 475448 249944 475454
rect 249892 475390 249944 475396
rect 249800 447296 249852 447302
rect 249800 447238 249852 447244
rect 247144 443958 247526 443986
rect 247972 443958 248354 443986
rect 248708 443958 249090 443986
rect 249904 443972 249932 475390
rect 250260 447296 250312 447302
rect 250260 447238 250312 447244
rect 250272 443986 250300 447238
rect 251192 443986 251220 476410
rect 252374 476368 252430 476377
rect 252374 476303 252430 476312
rect 252388 476202 252416 476303
rect 252466 476232 252522 476241
rect 252376 476196 252428 476202
rect 252466 476167 252522 476176
rect 252376 476138 252428 476144
rect 251272 474020 251324 474026
rect 251272 473962 251324 473968
rect 251284 460934 251312 473962
rect 251284 460906 251864 460934
rect 251836 443986 251864 460906
rect 252480 447098 252508 476167
rect 252560 476128 252612 476134
rect 252560 476070 252612 476076
rect 252468 447092 252520 447098
rect 252468 447034 252520 447040
rect 252572 443986 252600 476070
rect 252664 460934 252692 476478
rect 255332 476338 255360 477119
rect 259366 476912 259422 476921
rect 259366 476847 259422 476856
rect 255412 476672 255464 476678
rect 255412 476614 255464 476620
rect 258262 476640 258318 476649
rect 255320 476332 255372 476338
rect 255320 476274 255372 476280
rect 253846 476232 253902 476241
rect 253846 476167 253902 476176
rect 255226 476232 255282 476241
rect 255226 476167 255282 476176
rect 252664 460906 253336 460934
rect 253308 443986 253336 460906
rect 253860 447030 253888 476167
rect 253940 475380 253992 475386
rect 253940 475322 253992 475328
rect 253952 460934 253980 475322
rect 253952 460906 254072 460934
rect 253848 447024 253900 447030
rect 253848 446966 253900 446972
rect 254044 443986 254072 460906
rect 255240 446962 255268 476167
rect 255424 460934 255452 476614
rect 258262 476575 258318 476584
rect 258172 476400 258224 476406
rect 258172 476342 258224 476348
rect 256606 476232 256662 476241
rect 257986 476232 258042 476241
rect 256606 476167 256662 476176
rect 256700 476196 256752 476202
rect 255424 460906 255728 460934
rect 255320 447092 255372 447098
rect 255320 447034 255372 447040
rect 255228 446956 255280 446962
rect 255228 446898 255280 446904
rect 250272 443958 250654 443986
rect 251192 443958 251390 443986
rect 251836 443958 252218 443986
rect 252572 443958 252954 443986
rect 253308 443958 253782 443986
rect 254044 443958 254518 443986
rect 255332 443972 255360 447034
rect 255700 443986 255728 460906
rect 256620 446622 256648 476167
rect 257986 476167 258042 476176
rect 256700 476138 256752 476144
rect 256608 446616 256660 446622
rect 256608 446558 256660 446564
rect 256712 446418 256740 476138
rect 256792 457496 256844 457502
rect 256792 457438 256844 457444
rect 256700 446412 256752 446418
rect 256700 446354 256752 446360
rect 256804 443986 256832 457438
rect 258000 446486 258028 476167
rect 257988 446480 258040 446486
rect 257988 446422 258040 446428
rect 257252 446412 257304 446418
rect 257252 446354 257304 446360
rect 257264 443986 257292 446354
rect 258184 443986 258212 476342
rect 258276 476202 258304 476575
rect 258264 476196 258316 476202
rect 258264 476138 258316 476144
rect 259380 447030 259408 476847
rect 264992 476678 265020 477255
rect 264980 476672 265032 476678
rect 263598 476640 263654 476649
rect 259552 476604 259604 476610
rect 264980 476614 265032 476620
rect 263598 476575 263654 476584
rect 259552 476546 259604 476552
rect 259184 447024 259236 447030
rect 259184 446966 259236 446972
rect 259368 447024 259420 447030
rect 259368 446966 259420 446972
rect 255700 443958 256082 443986
rect 256804 443958 256910 443986
rect 257264 443958 257646 443986
rect 258184 443958 258474 443986
rect 259196 443972 259224 446966
rect 259564 443986 259592 476546
rect 263612 476542 263640 476575
rect 263600 476536 263652 476542
rect 260838 476504 260894 476513
rect 263600 476478 263652 476484
rect 265072 476536 265124 476542
rect 265072 476478 265124 476484
rect 260838 476439 260840 476448
rect 260892 476439 260894 476448
rect 260840 476410 260892 476416
rect 261482 476368 261538 476377
rect 260932 476332 260984 476338
rect 261482 476303 261538 476312
rect 263506 476368 263562 476377
rect 263506 476303 263562 476312
rect 263692 476332 263744 476338
rect 260932 476274 260984 476280
rect 260746 476232 260802 476241
rect 260746 476167 260802 476176
rect 260380 446956 260432 446962
rect 260380 446898 260432 446904
rect 260392 443986 260420 446898
rect 260760 446554 260788 476167
rect 260944 460934 260972 476274
rect 260944 460906 261064 460934
rect 260748 446548 260800 446554
rect 260748 446490 260800 446496
rect 261036 443986 261064 460906
rect 261496 446962 261524 476303
rect 262404 476264 262456 476270
rect 262404 476206 262456 476212
rect 262862 476232 262918 476241
rect 262416 460934 262444 476206
rect 262862 476167 262918 476176
rect 262416 460906 262720 460934
rect 261484 446956 261536 446962
rect 261484 446898 261536 446904
rect 262312 446616 262364 446622
rect 262312 446558 262364 446564
rect 259564 443958 259946 443986
rect 260392 443958 260774 443986
rect 261036 443958 261510 443986
rect 262324 443972 262352 446558
rect 262692 443986 262720 460906
rect 262876 447098 262904 476167
rect 263520 476134 263548 476303
rect 263692 476274 263744 476280
rect 263508 476128 263560 476134
rect 263508 476070 263560 476076
rect 263704 460934 263732 476274
rect 264886 476232 264942 476241
rect 264886 476167 264942 476176
rect 263704 460906 264192 460934
rect 262864 447092 262916 447098
rect 262864 447034 262916 447040
rect 263876 446480 263928 446486
rect 263876 446422 263928 446428
rect 262692 443958 263074 443986
rect 263888 443972 263916 446422
rect 264164 443986 264192 460906
rect 264900 446486 264928 476167
rect 265084 460934 265112 476478
rect 268028 476474 268056 477255
rect 280158 477048 280214 477057
rect 280158 476983 280214 476992
rect 304998 477048 305054 477057
rect 304998 476983 305054 476992
rect 307758 477048 307814 477057
rect 307758 476983 307814 476992
rect 277858 476912 277914 476921
rect 277858 476847 277914 476856
rect 270498 476776 270554 476785
rect 270498 476711 270554 476720
rect 270512 476610 270540 476711
rect 270500 476604 270552 476610
rect 270500 476546 270552 476552
rect 273258 476504 273314 476513
rect 268016 476468 268068 476474
rect 273258 476439 273314 476448
rect 268016 476410 268068 476416
rect 273272 476406 273300 476439
rect 273260 476400 273312 476406
rect 267554 476368 267610 476377
rect 273260 476342 273312 476348
rect 274546 476368 274602 476377
rect 267554 476303 267610 476312
rect 274546 476303 274602 476312
rect 276018 476368 276074 476377
rect 277872 476338 277900 476847
rect 278042 476776 278098 476785
rect 278042 476711 278098 476720
rect 276018 476303 276074 476312
rect 277860 476332 277912 476338
rect 266266 476232 266322 476241
rect 266266 476167 266322 476176
rect 265084 460906 265848 460934
rect 265440 447024 265492 447030
rect 265440 446966 265492 446972
rect 264888 446480 264940 446486
rect 264888 446422 264940 446428
rect 264164 443958 264638 443986
rect 265452 443972 265480 446966
rect 265820 443986 265848 460906
rect 266280 458998 266308 476167
rect 267004 476128 267056 476134
rect 267004 476070 267056 476076
rect 266268 458992 266320 458998
rect 266268 458934 266320 458940
rect 267016 446690 267044 476070
rect 267568 458930 267596 476303
rect 267646 476232 267702 476241
rect 269026 476232 269082 476241
rect 267646 476167 267702 476176
rect 267740 476196 267792 476202
rect 267556 458924 267608 458930
rect 267556 458866 267608 458872
rect 267660 457502 267688 476167
rect 269026 476167 269082 476176
rect 270406 476232 270462 476241
rect 270406 476167 270462 476176
rect 271786 476232 271842 476241
rect 271786 476167 271842 476176
rect 273166 476232 273222 476241
rect 273166 476167 273222 476176
rect 267740 476138 267792 476144
rect 267648 457496 267700 457502
rect 267648 457438 267700 457444
rect 267004 446684 267056 446690
rect 267004 446626 267056 446632
rect 267004 446548 267056 446554
rect 267004 446490 267056 446496
rect 265820 443958 266202 443986
rect 267016 443972 267044 446490
rect 267752 443972 267780 476138
rect 269040 457774 269068 476167
rect 269028 457768 269080 457774
rect 269028 457710 269080 457716
rect 270420 457706 270448 476167
rect 270592 460216 270644 460222
rect 270592 460158 270644 460164
rect 270408 457700 270460 457706
rect 270408 457642 270460 457648
rect 269212 456136 269264 456142
rect 269212 456078 269264 456084
rect 268476 447024 268528 447030
rect 268476 446966 268528 446972
rect 268488 443972 268516 446966
rect 269224 443986 269252 456078
rect 270040 447092 270092 447098
rect 270040 447034 270092 447040
rect 269224 443958 269330 443986
rect 270052 443972 270080 447034
rect 270604 443986 270632 460158
rect 271800 458862 271828 476167
rect 271972 461712 272024 461718
rect 271972 461654 272024 461660
rect 271984 460934 272012 461654
rect 271984 460906 272104 460934
rect 271788 458856 271840 458862
rect 271788 458798 271840 458804
rect 271604 446684 271656 446690
rect 271604 446626 271656 446632
rect 270604 443958 270894 443986
rect 271616 443972 271644 446626
rect 272076 443986 272104 460906
rect 273180 460290 273208 476167
rect 273260 461644 273312 461650
rect 273260 461586 273312 461592
rect 273272 460934 273300 461586
rect 273272 460906 273576 460934
rect 273168 460284 273220 460290
rect 273168 460226 273220 460232
rect 273168 446480 273220 446486
rect 273168 446422 273220 446428
rect 272076 443958 272458 443986
rect 273180 443972 273208 446422
rect 273548 443986 273576 460906
rect 274560 460358 274588 476303
rect 276032 476270 276060 476303
rect 277860 476274 277912 476280
rect 276020 476264 276072 476270
rect 275282 476232 275338 476241
rect 276020 476206 276072 476212
rect 276662 476232 276718 476241
rect 275282 476167 275338 476176
rect 276662 476167 276718 476176
rect 274548 460352 274600 460358
rect 274548 460294 274600 460300
rect 274640 458992 274692 458998
rect 274640 458934 274692 458940
rect 274652 443986 274680 458934
rect 275192 457632 275244 457638
rect 275192 457574 275244 457580
rect 275204 443986 275232 457574
rect 275296 446554 275324 476167
rect 276020 458924 276072 458930
rect 276020 458866 276072 458872
rect 275284 446548 275336 446554
rect 275284 446490 275336 446496
rect 276032 443986 276060 458866
rect 276572 457564 276624 457570
rect 276572 457506 276624 457512
rect 276584 444122 276612 457506
rect 276676 446622 276704 476167
rect 277400 457496 277452 457502
rect 277400 457438 277452 457444
rect 277952 457496 278004 457502
rect 277952 457438 278004 457444
rect 276664 446616 276716 446622
rect 276664 446558 276716 446564
rect 276584 444094 276704 444122
rect 276676 443986 276704 444094
rect 277412 443986 277440 457438
rect 277964 444122 277992 457438
rect 278056 446486 278084 476711
rect 280172 476542 280200 476983
rect 302238 476776 302294 476785
rect 280252 476740 280304 476746
rect 302238 476711 302240 476720
rect 280252 476682 280304 476688
rect 302292 476711 302294 476720
rect 302240 476682 302292 476688
rect 280160 476536 280212 476542
rect 280160 476478 280212 476484
rect 278686 476232 278742 476241
rect 278686 476167 278742 476176
rect 280066 476232 280122 476241
rect 280066 476167 280122 476176
rect 278700 456210 278728 476167
rect 280080 476134 280108 476167
rect 280068 476128 280120 476134
rect 280068 476070 280120 476076
rect 280264 470594 280292 476682
rect 305012 476678 305040 476983
rect 281540 476672 281592 476678
rect 281540 476614 281592 476620
rect 305000 476672 305052 476678
rect 305000 476614 305052 476620
rect 280172 470566 280292 470594
rect 279056 457768 279108 457774
rect 279056 457710 279108 457716
rect 278688 456204 278740 456210
rect 278688 456146 278740 456152
rect 278044 446480 278096 446486
rect 278044 446422 278096 446428
rect 277964 444094 278176 444122
rect 278148 443986 278176 444094
rect 279068 443986 279096 457710
rect 273548 443958 274022 443986
rect 274652 443958 274758 443986
rect 275204 443958 275586 443986
rect 276032 443958 276322 443986
rect 276676 443958 277058 443986
rect 277412 443958 277886 443986
rect 278148 443958 278622 443986
rect 279068 443958 279450 443986
rect 280172 443972 280200 470566
rect 280528 457700 280580 457706
rect 280528 457642 280580 457648
rect 280540 443986 280568 457642
rect 281552 443986 281580 476614
rect 307772 476610 307800 476983
rect 310518 476912 310574 476921
rect 310518 476847 310574 476856
rect 283104 476604 283156 476610
rect 283104 476546 283156 476552
rect 307760 476604 307812 476610
rect 307760 476546 307812 476552
rect 282918 476232 282974 476241
rect 282918 476167 282920 476176
rect 282972 476167 282974 476176
rect 282920 476138 282972 476144
rect 282184 476128 282236 476134
rect 282184 476070 282236 476076
rect 282092 458856 282144 458862
rect 282092 458798 282144 458804
rect 282104 444122 282132 458798
rect 282196 446690 282224 476070
rect 283012 460284 283064 460290
rect 283012 460226 283064 460232
rect 283024 447302 283052 460226
rect 283012 447296 283064 447302
rect 283012 447238 283064 447244
rect 282184 446684 282236 446690
rect 282184 446626 282236 446632
rect 282104 444094 282224 444122
rect 282196 443986 282224 444094
rect 283116 443986 283144 476546
rect 310532 476542 310560 476847
rect 284300 476536 284352 476542
rect 284300 476478 284352 476484
rect 310520 476536 310572 476542
rect 310520 476478 310572 476484
rect 283748 447296 283800 447302
rect 283748 447238 283800 447244
rect 283760 443986 283788 447238
rect 284312 443986 284340 476478
rect 285680 476468 285732 476474
rect 285680 476410 285732 476416
rect 285128 460352 285180 460358
rect 285128 460294 285180 460300
rect 285140 443986 285168 460294
rect 285692 451274 285720 476410
rect 287244 476400 287296 476406
rect 287244 476342 287296 476348
rect 285770 476232 285826 476241
rect 285770 476167 285826 476176
rect 287150 476232 287206 476241
rect 287150 476167 287206 476176
rect 285784 456142 285812 476167
rect 287164 460222 287192 476167
rect 287256 460934 287284 476342
rect 288532 476332 288584 476338
rect 288532 476274 288584 476280
rect 288544 460934 288572 476274
rect 292764 476264 292816 476270
rect 289910 476232 289966 476241
rect 292670 476232 292726 476241
rect 289910 476167 289966 476176
rect 290004 476196 290056 476202
rect 289924 461718 289952 476167
rect 292764 476206 292816 476212
rect 295338 476232 295394 476241
rect 292670 476167 292726 476176
rect 290004 476138 290056 476144
rect 289912 461712 289964 461718
rect 289912 461654 289964 461660
rect 290016 460934 290044 476138
rect 292684 461650 292712 476167
rect 292672 461644 292724 461650
rect 292672 461586 292724 461592
rect 287256 460906 287560 460934
rect 288544 460906 289216 460934
rect 290016 460906 290688 460934
rect 287152 460216 287204 460222
rect 287152 460158 287204 460164
rect 285772 456136 285824 456142
rect 285772 456078 285824 456084
rect 285692 451246 286088 451274
rect 286060 443986 286088 451246
rect 287152 446548 287204 446554
rect 287152 446490 287204 446496
rect 280540 443958 281014 443986
rect 281552 443958 281750 443986
rect 282196 443958 282578 443986
rect 283116 443958 283314 443986
rect 283760 443958 284142 443986
rect 284312 443958 284878 443986
rect 285140 443958 285614 443986
rect 286060 443958 286442 443986
rect 287164 443972 287192 446490
rect 287532 443986 287560 460906
rect 288716 446616 288768 446622
rect 288716 446558 288768 446564
rect 288348 446208 288400 446214
rect 288348 446150 288400 446156
rect 288360 444106 288388 446150
rect 288348 444100 288400 444106
rect 288348 444042 288400 444048
rect 287532 443958 288006 443986
rect 288728 443972 288756 446558
rect 289188 443986 289216 460906
rect 290280 446480 290332 446486
rect 290280 446422 290332 446428
rect 289188 443958 289570 443986
rect 290292 443972 290320 446422
rect 290660 443986 290688 460906
rect 291384 456204 291436 456210
rect 291384 456146 291436 456152
rect 291396 443986 291424 456146
rect 292776 443986 292804 476206
rect 295338 476167 295394 476176
rect 298098 476232 298154 476241
rect 298098 476167 298154 476176
rect 300858 476232 300914 476241
rect 300858 476167 300914 476176
rect 293960 476128 294012 476134
rect 293960 476070 294012 476076
rect 293408 446684 293460 446690
rect 293408 446626 293460 446632
rect 290660 443958 291134 443986
rect 291396 443958 291870 443986
rect 292698 443958 292804 443986
rect 293420 443972 293448 446626
rect 293972 443986 294000 476070
rect 295352 457638 295380 476167
rect 295340 457632 295392 457638
rect 295340 457574 295392 457580
rect 298112 457570 298140 476167
rect 298100 457564 298152 457570
rect 298100 457506 298152 457512
rect 300872 457502 300900 476167
rect 311912 460934 311940 478178
rect 354680 478168 354732 478174
rect 354680 478110 354732 478116
rect 322938 476776 322994 476785
rect 322938 476711 322994 476720
rect 313278 476504 313334 476513
rect 313278 476439 313280 476448
rect 313332 476439 313334 476448
rect 314658 476504 314714 476513
rect 314658 476439 314714 476448
rect 313280 476410 313332 476416
rect 314672 476406 314700 476439
rect 314660 476400 314712 476406
rect 314660 476342 314712 476348
rect 317418 476368 317474 476377
rect 317418 476303 317420 476312
rect 317472 476303 317474 476312
rect 320178 476368 320234 476377
rect 320178 476303 320234 476312
rect 317420 476274 317472 476280
rect 320192 476202 320220 476303
rect 322952 476270 322980 476711
rect 322940 476264 322992 476270
rect 322940 476206 322992 476212
rect 325790 476232 325846 476241
rect 320180 476196 320232 476202
rect 325790 476167 325846 476176
rect 320180 476138 320232 476144
rect 325804 476134 325832 476167
rect 325792 476128 325844 476134
rect 325792 476070 325844 476076
rect 333980 474768 334032 474774
rect 333980 474710 334032 474716
rect 333992 460934 334020 474710
rect 335360 462392 335412 462398
rect 335360 462334 335412 462340
rect 335372 460934 335400 462334
rect 311912 460906 312400 460934
rect 333992 460906 334296 460934
rect 335372 460906 335768 460934
rect 300860 457496 300912 457502
rect 300860 457438 300912 457444
rect 300860 456272 300912 456278
rect 300860 456214 300912 456220
rect 298376 456136 298428 456142
rect 298376 456078 298428 456084
rect 297272 450696 297324 450702
rect 297272 450638 297324 450644
rect 296534 446176 296590 446185
rect 296534 446111 296590 446120
rect 294970 446040 295026 446049
rect 294970 445975 295026 445984
rect 293972 443958 294170 443986
rect 294984 443972 295012 445975
rect 295706 445904 295762 445913
rect 295706 445839 295762 445848
rect 295720 443972 295748 445839
rect 296548 443972 296576 446111
rect 297284 443972 297312 450638
rect 298388 443986 298416 456078
rect 299664 450764 299716 450770
rect 299664 450706 299716 450712
rect 298388 443958 298862 443986
rect 299676 443972 299704 450706
rect 300398 444544 300454 444553
rect 300398 444479 300454 444488
rect 300412 443972 300440 444479
rect 300872 443986 300900 456214
rect 303160 456204 303212 456210
rect 303160 456146 303212 456152
rect 301964 450832 302016 450838
rect 301964 450774 302016 450780
rect 300872 443958 301254 443986
rect 301976 443972 302004 450774
rect 303172 443986 303200 456146
rect 310888 453552 310940 453558
rect 310888 453494 310940 453500
rect 303896 452260 303948 452266
rect 303896 452202 303948 452208
rect 303908 443986 303936 452202
rect 308496 452192 308548 452198
rect 308496 452134 308548 452140
rect 306380 452124 306432 452130
rect 306380 452066 306432 452072
rect 305828 449268 305880 449274
rect 305828 449210 305880 449216
rect 305092 445800 305144 445806
rect 305092 445742 305144 445748
rect 303172 443958 303554 443986
rect 303908 443958 304290 443986
rect 305104 443972 305132 445742
rect 305840 443972 305868 449210
rect 306392 443986 306420 452066
rect 308220 449404 308272 449410
rect 308220 449346 308272 449352
rect 307392 446616 307444 446622
rect 307392 446558 307444 446564
rect 306392 443958 306682 443986
rect 307404 443972 307432 446558
rect 308232 443972 308260 449346
rect 308508 443986 308536 452134
rect 310520 449540 310572 449546
rect 310520 449482 310572 449488
rect 309784 446412 309836 446418
rect 309784 446354 309836 446360
rect 308508 443958 308982 443986
rect 309796 443972 309824 446354
rect 310532 443972 310560 449482
rect 310900 443986 310928 453494
rect 312084 444984 312136 444990
rect 312084 444926 312136 444932
rect 310900 443958 311374 443986
rect 312096 443972 312124 444926
rect 312372 443986 312400 460906
rect 333520 456068 333572 456074
rect 333520 456010 333572 456016
rect 317420 454980 317472 454986
rect 317420 454922 317472 454928
rect 315948 446888 316000 446894
rect 315948 446830 316000 446836
rect 315212 446548 315264 446554
rect 315212 446490 315264 446496
rect 313648 446480 313700 446486
rect 313648 446422 313700 446428
rect 312372 443958 312846 443986
rect 313660 443972 313688 446422
rect 314384 446276 314436 446282
rect 314384 446218 314436 446224
rect 314396 443972 314424 446218
rect 315224 443972 315252 446490
rect 315960 443972 315988 446830
rect 316776 444576 316828 444582
rect 316776 444518 316828 444524
rect 316788 443972 316816 444518
rect 317432 443986 317460 454922
rect 331220 454912 331272 454918
rect 331220 454854 331272 454860
rect 325700 454844 325752 454850
rect 325700 454786 325752 454792
rect 325792 454844 325844 454850
rect 325792 454786 325844 454792
rect 323400 453688 323452 453694
rect 323400 453630 323452 453636
rect 321008 453620 321060 453626
rect 321008 453562 321060 453568
rect 319904 449472 319956 449478
rect 319904 449414 319956 449420
rect 318340 448112 318392 448118
rect 318340 448054 318392 448060
rect 317432 443958 317538 443986
rect 318352 443972 318380 448054
rect 318708 446344 318760 446350
rect 318708 446286 318760 446292
rect 318720 445058 318748 446286
rect 318708 445052 318760 445058
rect 318708 444994 318760 445000
rect 319076 444440 319128 444446
rect 319076 444382 319128 444388
rect 319088 443972 319116 444382
rect 319916 443972 319944 449414
rect 320640 447976 320692 447982
rect 320640 447918 320692 447924
rect 320652 443972 320680 447918
rect 321020 443986 321048 453562
rect 322204 449336 322256 449342
rect 322204 449278 322256 449284
rect 321020 443958 321402 443986
rect 322216 443972 322244 449278
rect 322940 447908 322992 447914
rect 322940 447850 322992 447856
rect 322952 443972 322980 447850
rect 323412 443986 323440 453630
rect 325332 450628 325384 450634
rect 325332 450570 325384 450576
rect 324504 449200 324556 449206
rect 324504 449142 324556 449148
rect 323412 443958 323794 443986
rect 324516 443972 324544 449142
rect 325344 443972 325372 450570
rect 325712 447302 325740 454786
rect 325700 447296 325752 447302
rect 325700 447238 325752 447244
rect 325804 443986 325832 454786
rect 328736 454776 328788 454782
rect 328736 454718 328788 454724
rect 329840 454776 329892 454782
rect 329840 454718 329892 454724
rect 327632 450560 327684 450566
rect 327632 450502 327684 450508
rect 326620 447296 326672 447302
rect 326620 447238 326672 447244
rect 326632 443986 326660 447238
rect 325804 443958 326094 443986
rect 326632 443958 326922 443986
rect 327644 443972 327672 450502
rect 328460 447908 328512 447914
rect 328460 447850 328512 447856
rect 328472 443972 328500 447850
rect 328748 443986 328776 454718
rect 329852 447302 329880 454718
rect 329932 451920 329984 451926
rect 329932 451862 329984 451868
rect 329840 447296 329892 447302
rect 329840 447238 329892 447244
rect 328748 443958 329222 443986
rect 329944 443972 329972 451862
rect 330484 447296 330536 447302
rect 330484 447238 330536 447244
rect 330496 443986 330524 447238
rect 331232 443986 331260 454854
rect 331864 451988 331916 451994
rect 331864 451930 331916 451936
rect 331876 443986 331904 451930
rect 333060 447976 333112 447982
rect 333060 447918 333112 447924
rect 330496 443958 330786 443986
rect 331232 443958 331522 443986
rect 331876 443958 332350 443986
rect 333072 443972 333100 447918
rect 333532 443986 333560 456010
rect 334268 443986 334296 460906
rect 335452 450560 335504 450566
rect 335452 450502 335504 450508
rect 333532 443958 333914 443986
rect 334268 443958 334650 443986
rect 335464 443972 335492 450502
rect 335740 443986 335768 460906
rect 337384 454912 337436 454918
rect 337384 454854 337436 454860
rect 337016 445120 337068 445126
rect 337016 445062 337068 445068
rect 335740 443958 336214 443986
rect 337028 443972 337056 445062
rect 337396 443986 337424 454854
rect 353760 453484 353812 453490
rect 353760 453426 353812 453432
rect 353392 453416 353444 453422
rect 353392 453358 353444 453364
rect 351368 453348 351420 453354
rect 351368 453290 351420 453296
rect 349252 452056 349304 452062
rect 349252 451998 349304 452004
rect 344744 448180 344796 448186
rect 344744 448122 344796 448128
rect 340052 446684 340104 446690
rect 340052 446626 340104 446632
rect 338488 446140 338540 446146
rect 338488 446082 338540 446088
rect 337396 443958 337778 443986
rect 338500 443972 338528 446082
rect 338764 445800 338816 445806
rect 338764 445742 338816 445748
rect 338776 445058 338804 445742
rect 338764 445052 338816 445058
rect 338764 444994 338816 445000
rect 339316 444644 339368 444650
rect 339316 444586 339368 444592
rect 339328 443972 339356 444586
rect 340064 443972 340092 446626
rect 340880 446616 340932 446622
rect 340880 446558 340932 446564
rect 342444 446616 342496 446622
rect 342444 446558 342496 446564
rect 340892 445126 340920 446558
rect 340880 445120 340932 445126
rect 340880 445062 340932 445068
rect 340880 444916 340932 444922
rect 340880 444858 340932 444864
rect 340892 443972 340920 444858
rect 341616 444712 341668 444718
rect 341616 444654 341668 444660
rect 341628 443972 341656 444654
rect 342456 443972 342484 446558
rect 343180 446072 343232 446078
rect 343180 446014 343232 446020
rect 343272 446072 343324 446078
rect 343272 446014 343324 446020
rect 343192 443972 343220 446014
rect 233884 443896 233936 443902
rect 233884 443838 233936 443844
rect 343284 443766 343312 446014
rect 344008 444848 344060 444854
rect 344008 444790 344060 444796
rect 344020 443972 344048 444790
rect 344756 443972 344784 448122
rect 347044 448044 347096 448050
rect 347044 447986 347096 447992
rect 345940 446820 345992 446826
rect 345940 446762 345992 446768
rect 345572 445188 345624 445194
rect 345572 445130 345624 445136
rect 345584 443972 345612 445130
rect 345952 443986 345980 446762
rect 346308 446412 346360 446418
rect 346308 446354 346360 446360
rect 346320 445194 346348 446354
rect 346308 445188 346360 445194
rect 346308 445130 346360 445136
rect 345952 443958 346334 443986
rect 347056 443972 347084 447986
rect 347872 446004 347924 446010
rect 347872 445946 347924 445952
rect 347884 443972 347912 445946
rect 348608 444780 348660 444786
rect 348608 444722 348660 444728
rect 348620 443972 348648 444722
rect 349264 443986 349292 451998
rect 350172 444508 350224 444514
rect 350172 444450 350224 444456
rect 349264 443958 349462 443986
rect 350184 443972 350212 444450
rect 350998 444408 351054 444417
rect 350998 444343 351054 444352
rect 351012 443972 351040 444343
rect 351380 443986 351408 453290
rect 352564 445936 352616 445942
rect 352564 445878 352616 445884
rect 351920 445800 351972 445806
rect 351920 445742 351972 445748
rect 351380 443958 351762 443986
rect 343272 443760 343324 443766
rect 343272 443702 343324 443708
rect 351932 443698 351960 445742
rect 352576 443972 352604 445878
rect 353404 443986 353432 453358
rect 353326 443958 353432 443986
rect 353772 443986 353800 453426
rect 354692 447302 354720 478110
rect 354772 454708 354824 454714
rect 354772 454650 354824 454656
rect 354680 447296 354732 447302
rect 354680 447238 354732 447244
rect 354784 443986 354812 454650
rect 356428 447840 356480 447846
rect 356428 447782 356480 447788
rect 355324 447296 355376 447302
rect 355324 447238 355376 447244
rect 355336 443986 355364 447238
rect 353772 443958 354154 443986
rect 354784 443958 354890 443986
rect 355336 443958 355626 443986
rect 356440 443972 356468 447782
rect 357452 446622 357480 700266
rect 357440 446616 357492 446622
rect 357440 446558 357492 446564
rect 357544 446486 357572 700402
rect 358820 700392 358872 700398
rect 358820 700334 358872 700340
rect 358084 700324 358136 700330
rect 358084 700266 358136 700272
rect 358096 452266 358124 700266
rect 358176 670744 358228 670750
rect 358176 670686 358228 670692
rect 358084 452260 358136 452266
rect 358084 452202 358136 452208
rect 358188 450838 358216 670686
rect 358268 536852 358320 536858
rect 358268 536794 358320 536800
rect 358280 453694 358308 536794
rect 358360 484424 358412 484430
rect 358360 484366 358412 484372
rect 358268 453688 358320 453694
rect 358268 453630 358320 453636
rect 358372 453626 358400 484366
rect 358360 453620 358412 453626
rect 358360 453562 358412 453568
rect 358176 450832 358228 450838
rect 358176 450774 358228 450780
rect 358832 446554 358860 700334
rect 358924 478242 358952 700470
rect 359464 700392 359516 700398
rect 359464 700334 359516 700340
rect 359004 565140 359056 565146
rect 359004 565082 359056 565088
rect 358912 478236 358964 478242
rect 358912 478178 358964 478184
rect 359016 446690 359044 565082
rect 359476 454918 359504 700334
rect 364996 699718 365024 703520
rect 397472 700398 397500 703520
rect 397460 700392 397512 700398
rect 397460 700334 397512 700340
rect 360844 699712 360896 699718
rect 360844 699654 360896 699660
rect 364984 699712 365036 699718
rect 364984 699654 365036 699660
rect 359556 696992 359608 696998
rect 359556 696934 359608 696940
rect 359464 454912 359516 454918
rect 359464 454854 359516 454860
rect 359568 454782 359596 696934
rect 359648 616888 359700 616894
rect 359648 616830 359700 616836
rect 359556 454776 359608 454782
rect 359556 454718 359608 454724
rect 359660 450770 359688 616830
rect 360856 453558 360884 699654
rect 362224 630692 362276 630698
rect 362224 630634 362276 630640
rect 362236 456278 362264 630634
rect 362316 590708 362368 590714
rect 362316 590650 362368 590656
rect 362224 456272 362276 456278
rect 362224 456214 362276 456220
rect 362328 454850 362356 590650
rect 371884 563100 371936 563106
rect 371884 563042 371936 563048
rect 362316 454844 362368 454850
rect 362316 454786 362368 454792
rect 360844 453552 360896 453558
rect 360844 453494 360896 453500
rect 359648 450764 359700 450770
rect 359648 450706 359700 450712
rect 371896 450702 371924 563042
rect 371884 450696 371936 450702
rect 371884 450638 371936 450644
rect 412652 449546 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 429212 452198 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 429200 452192 429252 452198
rect 429200 452134 429252 452140
rect 462332 450566 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 462320 450560 462372 450566
rect 462320 450502 462372 450508
rect 412640 449540 412692 449546
rect 412640 449482 412692 449488
rect 477512 449410 477540 702406
rect 494072 452130 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 494060 452124 494112 452130
rect 494060 452066 494112 452072
rect 477500 449404 477552 449410
rect 477500 449346 477552 449352
rect 527192 447982 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 542372 449274 542400 702406
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580262 683904 580318 683913
rect 580262 683839 580318 683848
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579618 591016 579674 591025
rect 579618 590951 579674 590960
rect 579632 590714 579660 590951
rect 579620 590708 579672 590714
rect 579620 590650 579672 590656
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563106 580212 564295
rect 580172 563100 580224 563106
rect 580172 563042 580224 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 580276 456210 580304 683839
rect 580354 644056 580410 644065
rect 580354 643991 580410 644000
rect 580264 456204 580316 456210
rect 580264 456146 580316 456152
rect 542360 449268 542412 449274
rect 542360 449210 542412 449216
rect 527180 447976 527232 447982
rect 527180 447918 527232 447924
rect 580368 447914 580396 643991
rect 580446 577688 580502 577697
rect 580446 577623 580502 577632
rect 580460 456142 580488 577623
rect 580448 456136 580500 456142
rect 580448 456078 580500 456084
rect 580356 447908 580408 447914
rect 580356 447850 580408 447856
rect 359004 446684 359056 446690
rect 359004 446626 359056 446632
rect 358820 446548 358872 446554
rect 358820 446490 358872 446496
rect 357532 446480 357584 446486
rect 357532 446422 357584 446428
rect 357992 446344 358044 446350
rect 357992 446286 358044 446292
rect 357164 446072 357216 446078
rect 357164 446014 357216 446020
rect 357176 443972 357204 446014
rect 358004 443972 358032 446286
rect 364984 446276 365036 446282
rect 364984 446218 365036 446224
rect 359556 446208 359608 446214
rect 359556 446150 359608 446156
rect 358728 445800 358780 445806
rect 358728 445742 358780 445748
rect 358740 443972 358768 445742
rect 359568 443972 359596 446150
rect 360292 445868 360344 445874
rect 360292 445810 360344 445816
rect 360304 443972 360332 445810
rect 351920 443692 351972 443698
rect 351920 443634 351972 443640
rect 320824 443624 320876 443630
rect 320824 443566 320876 443572
rect 320836 443494 320864 443566
rect 298192 443488 298244 443494
rect 298126 443436 298192 443442
rect 303160 443488 303212 443494
rect 298126 443430 298244 443436
rect 302818 443436 303160 443442
rect 302818 443430 303212 443436
rect 320824 443488 320876 443494
rect 320824 443430 320876 443436
rect 360844 443488 360896 443494
rect 362222 443456 362278 443465
rect 360896 443436 361146 443442
rect 360844 443430 361146 443436
rect 298126 443414 298232 443430
rect 302818 443414 303200 443430
rect 360856 443414 361146 443430
rect 361882 443414 362222 443442
rect 362774 443456 362830 443465
rect 362710 443414 362774 443442
rect 362222 443391 362278 443400
rect 362774 443391 362830 443400
rect 363050 443456 363106 443465
rect 363106 443414 363446 443442
rect 363050 443391 363106 443400
rect 232240 412606 232360 412634
rect 232240 411262 232268 412606
rect 232228 411256 232280 411262
rect 232228 411198 232280 411204
rect 231216 358760 231268 358766
rect 231216 358702 231268 358708
rect 364996 325650 365024 446218
rect 558182 446176 558238 446185
rect 558182 446111 558238 446120
rect 554042 445904 554098 445913
rect 554042 445839 554098 445848
rect 367744 444984 367796 444990
rect 367744 444926 367796 444932
rect 365076 444576 365128 444582
rect 365076 444518 365128 444524
rect 365088 379506 365116 444518
rect 365168 444440 365220 444446
rect 365168 444382 365220 444388
rect 365180 431934 365208 444382
rect 365168 431928 365220 431934
rect 365168 431870 365220 431876
rect 365076 379500 365128 379506
rect 365076 379442 365128 379448
rect 364984 325644 365036 325650
rect 364984 325586 365036 325592
rect 305196 310554 305394 310570
rect 305000 310548 305052 310554
rect 305000 310490 305052 310496
rect 305184 310548 305394 310554
rect 305236 310542 305394 310548
rect 306498 310542 306696 310570
rect 309258 310554 309456 310570
rect 310638 310554 310836 310570
rect 312018 310554 312216 310570
rect 309258 310548 309468 310554
rect 309258 310542 309416 310548
rect 305184 310490 305236 310496
rect 231872 310406 232530 310434
rect 231768 308440 231820 308446
rect 231768 308382 231820 308388
rect 231780 308106 231808 308382
rect 231768 308100 231820 308106
rect 231768 308042 231820 308048
rect 231124 258800 231176 258806
rect 231124 258742 231176 258748
rect 231872 258738 231900 310406
rect 231952 308440 232004 308446
rect 232700 308394 232728 310420
rect 232792 310406 232990 310434
rect 232792 308446 232820 310406
rect 233056 308508 233108 308514
rect 233056 308450 233108 308456
rect 231952 308382 232004 308388
rect 231860 258732 231912 258738
rect 231860 258674 231912 258680
rect 231964 244934 231992 308382
rect 232056 308366 232728 308394
rect 232780 308440 232832 308446
rect 232780 308382 232832 308388
rect 232056 245002 232084 308366
rect 233068 308038 233096 308450
rect 233056 308032 233108 308038
rect 233056 307974 233108 307980
rect 233160 296714 233188 310420
rect 233436 308553 233464 310420
rect 233422 308544 233478 308553
rect 233332 308508 233384 308514
rect 233422 308479 233478 308488
rect 233332 308450 233384 308456
rect 233240 308440 233292 308446
rect 233240 308382 233292 308388
rect 232148 296686 233188 296714
rect 232148 247722 232176 296686
rect 232136 247716 232188 247722
rect 232136 247658 232188 247664
rect 233252 245070 233280 308382
rect 233344 253230 233372 308450
rect 233620 308394 233648 310420
rect 233712 310406 233910 310434
rect 233712 308446 233740 310406
rect 233436 308366 233648 308394
rect 233700 308440 233752 308446
rect 233700 308382 233752 308388
rect 233436 256018 233464 308366
rect 234080 296714 234108 310420
rect 234172 310406 234370 310434
rect 234172 308514 234200 310406
rect 234160 308508 234212 308514
rect 234160 308450 234212 308456
rect 234540 308417 234568 310420
rect 234632 310406 234830 310434
rect 234526 308408 234582 308417
rect 234526 308343 234582 308352
rect 233528 296686 234108 296714
rect 233528 260166 233556 296686
rect 233516 260160 233568 260166
rect 233516 260102 233568 260108
rect 233424 256012 233476 256018
rect 233424 255954 233476 255960
rect 233332 253224 233384 253230
rect 233332 253166 233384 253172
rect 234632 249082 234660 310406
rect 234804 306468 234856 306474
rect 234804 306410 234856 306416
rect 234712 306400 234764 306406
rect 234712 306342 234764 306348
rect 234724 250510 234752 306342
rect 234816 253366 234844 306410
rect 235000 306354 235028 310420
rect 234908 306326 235028 306354
rect 235092 310406 235290 310434
rect 234804 253360 234856 253366
rect 234804 253302 234856 253308
rect 234908 253298 234936 306326
rect 234988 305380 235040 305386
rect 234988 305322 235040 305328
rect 235000 256086 235028 305322
rect 235092 269822 235120 310406
rect 235460 305386 235488 310420
rect 235552 310406 235750 310434
rect 235552 306406 235580 310406
rect 235920 306474 235948 310420
rect 236196 308106 236224 310420
rect 236380 308718 236408 310420
rect 236472 310406 236670 310434
rect 236368 308712 236420 308718
rect 236368 308654 236420 308660
rect 236184 308100 236236 308106
rect 236184 308042 236236 308048
rect 236092 306536 236144 306542
rect 236092 306478 236144 306484
rect 235908 306468 235960 306474
rect 235908 306410 235960 306416
rect 235540 306400 235592 306406
rect 235540 306342 235592 306348
rect 235448 305380 235500 305386
rect 235448 305322 235500 305328
rect 235080 269816 235132 269822
rect 235080 269758 235132 269764
rect 236104 256154 236132 306478
rect 236184 306468 236236 306474
rect 236184 306410 236236 306416
rect 236196 267034 236224 306410
rect 236276 306400 236328 306406
rect 236276 306342 236328 306348
rect 236288 279478 236316 306342
rect 236472 296714 236500 310406
rect 236840 306474 236868 310420
rect 236932 310406 237130 310434
rect 236828 306468 236880 306474
rect 236828 306410 236880 306416
rect 236932 306406 236960 310406
rect 237300 306542 237328 310420
rect 237288 306536 237340 306542
rect 237288 306478 237340 306484
rect 237576 306474 237604 310420
rect 237564 306468 237616 306474
rect 237564 306410 237616 306416
rect 236920 306400 236972 306406
rect 236920 306342 236972 306348
rect 237472 306400 237524 306406
rect 237760 306354 237788 310420
rect 238036 308038 238064 310420
rect 238024 308032 238076 308038
rect 238024 307974 238076 307980
rect 237840 306468 237892 306474
rect 237840 306410 237892 306416
rect 237472 306342 237524 306348
rect 236380 296686 236500 296714
rect 236276 279472 236328 279478
rect 236276 279414 236328 279420
rect 236184 267028 236236 267034
rect 236184 266970 236236 266976
rect 236092 256148 236144 256154
rect 236092 256090 236144 256096
rect 234988 256080 235040 256086
rect 234988 256022 235040 256028
rect 234896 253292 234948 253298
rect 234896 253234 234948 253240
rect 236380 251870 236408 296686
rect 237484 252006 237512 306342
rect 237576 306326 237788 306354
rect 237576 271182 237604 306326
rect 237656 305380 237708 305386
rect 237656 305322 237708 305328
rect 237668 272542 237696 305322
rect 237748 305312 237800 305318
rect 237748 305254 237800 305260
rect 237760 280838 237788 305254
rect 237748 280832 237800 280838
rect 237748 280774 237800 280780
rect 237656 272536 237708 272542
rect 237656 272478 237708 272484
rect 237564 271176 237616 271182
rect 237564 271118 237616 271124
rect 237472 252000 237524 252006
rect 237472 251942 237524 251948
rect 237852 251938 237880 306410
rect 238220 306406 238248 310420
rect 238312 310406 238510 310434
rect 238208 306400 238260 306406
rect 238208 306342 238260 306348
rect 238312 305386 238340 310406
rect 238300 305380 238352 305386
rect 238300 305322 238352 305328
rect 238680 305318 238708 310420
rect 238852 306400 238904 306406
rect 238852 306342 238904 306348
rect 238668 305312 238720 305318
rect 238668 305254 238720 305260
rect 238864 258874 238892 306342
rect 238956 261526 238984 310420
rect 239140 306354 239168 310420
rect 239416 308582 239444 310420
rect 239404 308576 239456 308582
rect 239404 308518 239456 308524
rect 239600 306406 239628 310420
rect 239692 310406 239890 310434
rect 239048 306326 239168 306354
rect 239588 306400 239640 306406
rect 239588 306342 239640 306348
rect 239048 273970 239076 306326
rect 239128 305380 239180 305386
rect 239128 305322 239180 305328
rect 239140 284986 239168 305322
rect 239692 296714 239720 310406
rect 240060 305386 240088 310420
rect 240232 306468 240284 306474
rect 240232 306410 240284 306416
rect 240048 305380 240100 305386
rect 240048 305322 240100 305328
rect 239232 296686 239720 296714
rect 239128 284980 239180 284986
rect 239128 284922 239180 284928
rect 239036 273964 239088 273970
rect 239036 273906 239088 273912
rect 238944 261520 238996 261526
rect 238944 261462 238996 261468
rect 238852 258868 238904 258874
rect 238852 258810 238904 258816
rect 239232 254590 239260 296686
rect 240244 254658 240272 306410
rect 240336 262886 240364 310420
rect 240416 306400 240468 306406
rect 240416 306342 240468 306348
rect 240428 264246 240456 306342
rect 240520 283626 240548 310420
rect 240796 308650 240824 310420
rect 240784 308644 240836 308650
rect 240784 308586 240836 308592
rect 240980 306406 241008 310420
rect 241072 310406 241270 310434
rect 241072 306474 241100 310406
rect 241060 306468 241112 306474
rect 241060 306410 241112 306416
rect 240968 306400 241020 306406
rect 240968 306342 241020 306348
rect 241440 296714 241468 310420
rect 240612 296686 241468 296714
rect 241532 310406 241730 310434
rect 240508 283620 240560 283626
rect 240508 283562 240560 283568
rect 240416 264240 240468 264246
rect 240416 264182 240468 264188
rect 240324 262880 240376 262886
rect 240324 262822 240376 262828
rect 240612 254862 240640 296686
rect 240600 254856 240652 254862
rect 240600 254798 240652 254804
rect 240232 254652 240284 254658
rect 240232 254594 240284 254600
rect 239220 254584 239272 254590
rect 239220 254526 239272 254532
rect 237840 251932 237892 251938
rect 237840 251874 237892 251880
rect 236368 251864 236420 251870
rect 236368 251806 236420 251812
rect 234712 250504 234764 250510
rect 234712 250446 234764 250452
rect 234620 249076 234672 249082
rect 234620 249018 234672 249024
rect 241532 246362 241560 310406
rect 241612 306400 241664 306406
rect 241900 306354 241928 310420
rect 241612 306342 241664 306348
rect 241624 258942 241652 306342
rect 241716 306326 241928 306354
rect 241992 310406 242190 310434
rect 241716 265674 241744 306326
rect 241796 305380 241848 305386
rect 241796 305322 241848 305328
rect 241808 268394 241836 305322
rect 241992 302234 242020 310406
rect 242360 306406 242388 310420
rect 242452 310406 242650 310434
rect 242348 306400 242400 306406
rect 242348 306342 242400 306348
rect 242452 305386 242480 310406
rect 242440 305380 242492 305386
rect 242440 305322 242492 305328
rect 241900 302206 242020 302234
rect 241900 286346 241928 302206
rect 242820 296714 242848 310420
rect 241992 296686 242848 296714
rect 242912 310406 243110 310434
rect 241992 287706 242020 296686
rect 241980 287700 242032 287706
rect 241980 287642 242032 287648
rect 241888 286340 241940 286346
rect 241888 286282 241940 286288
rect 241796 268388 241848 268394
rect 241796 268330 241848 268336
rect 241704 265668 241756 265674
rect 241704 265610 241756 265616
rect 241612 258936 241664 258942
rect 241612 258878 241664 258884
rect 242912 246430 242940 310406
rect 243280 306746 243308 310420
rect 243372 310406 243570 310434
rect 243268 306740 243320 306746
rect 243268 306682 243320 306688
rect 243268 306536 243320 306542
rect 243268 306478 243320 306484
rect 243084 306468 243136 306474
rect 243084 306410 243136 306416
rect 242992 306400 243044 306406
rect 242992 306342 243044 306348
rect 243004 246498 243032 306342
rect 243096 254794 243124 306410
rect 243176 300892 243228 300898
rect 243176 300834 243228 300840
rect 243084 254788 243136 254794
rect 243084 254730 243136 254736
rect 243188 254726 243216 300834
rect 243280 275330 243308 306478
rect 243372 300898 243400 310406
rect 243740 306406 243768 310420
rect 243832 310406 244030 310434
rect 243728 306400 243780 306406
rect 243728 306342 243780 306348
rect 243360 300892 243412 300898
rect 243360 300834 243412 300840
rect 243832 296714 243860 310406
rect 244200 306474 244228 310420
rect 244384 310406 244490 310434
rect 244384 308174 244412 310406
rect 244660 308496 244688 310420
rect 244476 308468 244688 308496
rect 244752 310406 244950 310434
rect 244372 308168 244424 308174
rect 244372 308110 244424 308116
rect 244372 308032 244424 308038
rect 244372 307974 244424 307980
rect 244188 306468 244240 306474
rect 244188 306410 244240 306416
rect 243372 296686 243860 296714
rect 243372 276690 243400 296686
rect 243360 276684 243412 276690
rect 243360 276626 243412 276632
rect 243268 275324 243320 275330
rect 243268 275266 243320 275272
rect 244384 267102 244412 307974
rect 244476 278050 244504 308468
rect 244752 308394 244780 310406
rect 244660 308366 244780 308394
rect 244556 308100 244608 308106
rect 244556 308042 244608 308048
rect 244568 280906 244596 308042
rect 244660 289134 244688 308366
rect 244740 308168 244792 308174
rect 244740 308110 244792 308116
rect 244648 289128 244700 289134
rect 244648 289070 244700 289076
rect 244556 280900 244608 280906
rect 244556 280842 244608 280848
rect 244464 278044 244516 278050
rect 244464 277986 244516 277992
rect 244372 267096 244424 267102
rect 244372 267038 244424 267044
rect 244752 260234 244780 308110
rect 245120 308038 245148 310420
rect 245212 310406 245410 310434
rect 245212 308106 245240 310406
rect 245200 308100 245252 308106
rect 245200 308042 245252 308048
rect 245108 308032 245160 308038
rect 245108 307974 245160 307980
rect 245580 307086 245608 310420
rect 245672 310406 245870 310434
rect 245568 307080 245620 307086
rect 245568 307022 245620 307028
rect 244740 260228 244792 260234
rect 244740 260170 244792 260176
rect 243176 254720 243228 254726
rect 243176 254662 243228 254668
rect 245672 247790 245700 310406
rect 246040 308394 246068 310420
rect 245856 308366 246068 308394
rect 246132 310406 246330 310434
rect 245752 307012 245804 307018
rect 245752 306954 245804 306960
rect 245764 250578 245792 306954
rect 245856 282198 245884 308366
rect 245936 308168 245988 308174
rect 245936 308110 245988 308116
rect 245948 283694 245976 308110
rect 246028 308100 246080 308106
rect 246028 308042 246080 308048
rect 246040 290562 246068 308042
rect 246028 290556 246080 290562
rect 246028 290498 246080 290504
rect 246132 290494 246160 310406
rect 246500 307018 246528 310420
rect 246592 310406 246790 310434
rect 246592 308174 246620 310406
rect 246580 308168 246632 308174
rect 246580 308110 246632 308116
rect 246960 308106 246988 310420
rect 247052 310406 247250 310434
rect 246948 308100 247000 308106
rect 246948 308042 247000 308048
rect 246488 307012 246540 307018
rect 246488 306954 246540 306960
rect 246120 290488 246172 290494
rect 246120 290430 246172 290436
rect 245936 283688 245988 283694
rect 245936 283630 245988 283636
rect 245844 282192 245896 282198
rect 245844 282134 245896 282140
rect 247052 250646 247080 310406
rect 247224 308508 247276 308514
rect 247224 308450 247276 308456
rect 247132 308440 247184 308446
rect 247132 308382 247184 308388
rect 247144 250714 247172 308382
rect 247236 253434 247264 308450
rect 247420 308394 247448 310420
rect 247328 308366 247448 308394
rect 247512 310406 247710 310434
rect 247328 285054 247356 308366
rect 247512 308258 247540 310406
rect 247880 308446 247908 310420
rect 247972 310406 248170 310434
rect 247972 308514 248000 310406
rect 247960 308508 248012 308514
rect 247960 308450 248012 308456
rect 247868 308440 247920 308446
rect 247868 308382 247920 308388
rect 247420 308230 247540 308258
rect 247420 290630 247448 308230
rect 248340 296714 248368 310420
rect 248524 310406 248630 310434
rect 248420 308508 248472 308514
rect 248420 308450 248472 308456
rect 247512 296686 248368 296714
rect 247512 290698 247540 296686
rect 247500 290692 247552 290698
rect 247500 290634 247552 290640
rect 247408 290624 247460 290630
rect 247408 290566 247460 290572
rect 247316 285048 247368 285054
rect 247316 284990 247368 284996
rect 248432 253502 248460 308450
rect 248524 269890 248552 310406
rect 248604 308576 248656 308582
rect 248604 308518 248656 308524
rect 248616 271250 248644 308518
rect 248800 308514 248828 310420
rect 248892 310406 249090 310434
rect 249168 310406 249366 310434
rect 248788 308508 248840 308514
rect 248788 308450 248840 308456
rect 248696 308440 248748 308446
rect 248696 308382 248748 308388
rect 248708 285122 248736 308382
rect 248892 296714 248920 310406
rect 249168 308582 249196 310406
rect 249156 308576 249208 308582
rect 249156 308518 249208 308524
rect 249536 308446 249564 310420
rect 249524 308440 249576 308446
rect 249524 308382 249576 308388
rect 248800 296686 248920 296714
rect 248800 291854 248828 296686
rect 249812 291922 249840 310420
rect 249892 308440 249944 308446
rect 249892 308382 249944 308388
rect 249800 291916 249852 291922
rect 249800 291858 249852 291864
rect 248788 291848 248840 291854
rect 248788 291790 248840 291796
rect 248696 285116 248748 285122
rect 248696 285058 248748 285064
rect 249904 282266 249932 308382
rect 249996 308174 250024 310420
rect 250088 310406 250286 310434
rect 249984 308168 250036 308174
rect 249984 308110 250036 308116
rect 249984 308032 250036 308038
rect 249984 307974 250036 307980
rect 249996 285190 250024 307974
rect 250088 286414 250116 310406
rect 250456 308394 250484 310420
rect 250548 310406 250746 310434
rect 250548 308446 250576 310406
rect 250180 308366 250484 308394
rect 250536 308440 250588 308446
rect 250536 308382 250588 308388
rect 250180 291990 250208 308366
rect 250260 308168 250312 308174
rect 250260 308110 250312 308116
rect 250168 291984 250220 291990
rect 250168 291926 250220 291932
rect 250076 286408 250128 286414
rect 250076 286350 250128 286356
rect 249984 285184 250036 285190
rect 249984 285126 250036 285132
rect 249892 282260 249944 282266
rect 249892 282202 249944 282208
rect 250272 279546 250300 308110
rect 250916 308038 250944 310420
rect 250904 308032 250956 308038
rect 250904 307974 250956 307980
rect 251192 292058 251220 310420
rect 251376 307816 251404 310420
rect 251284 307788 251404 307816
rect 251468 310406 251666 310434
rect 251180 292052 251232 292058
rect 251180 291994 251232 292000
rect 251284 282334 251312 307788
rect 251364 307692 251416 307698
rect 251364 307634 251416 307640
rect 251376 283762 251404 307634
rect 251468 286482 251496 310406
rect 251548 308440 251600 308446
rect 251548 308382 251600 308388
rect 251560 286550 251588 308382
rect 251836 296714 251864 310420
rect 251928 310406 252126 310434
rect 251928 307698 251956 310406
rect 252296 308446 252324 310420
rect 252572 308666 252600 310420
rect 252770 310406 252968 310434
rect 252572 308638 252876 308666
rect 252744 308508 252796 308514
rect 252744 308450 252796 308456
rect 252284 308440 252336 308446
rect 252284 308382 252336 308388
rect 252652 308440 252704 308446
rect 252652 308382 252704 308388
rect 251916 307692 251968 307698
rect 251916 307634 251968 307640
rect 251652 296686 251864 296714
rect 251548 286544 251600 286550
rect 251548 286486 251600 286492
rect 251456 286476 251508 286482
rect 251456 286418 251508 286424
rect 251364 283756 251416 283762
rect 251364 283698 251416 283704
rect 251272 282328 251324 282334
rect 251272 282270 251324 282276
rect 250260 279540 250312 279546
rect 250260 279482 250312 279488
rect 248604 271244 248656 271250
rect 248604 271186 248656 271192
rect 248512 269884 248564 269890
rect 248512 269826 248564 269832
rect 248420 253496 248472 253502
rect 248420 253438 248472 253444
rect 247224 253428 247276 253434
rect 247224 253370 247276 253376
rect 251652 250782 251680 296686
rect 252664 283830 252692 308382
rect 252756 287774 252784 308450
rect 252848 308258 252876 308638
rect 252940 308394 252968 310406
rect 253032 308514 253060 310420
rect 253216 308786 253244 310420
rect 253308 310406 253506 310434
rect 253204 308780 253256 308786
rect 253204 308722 253256 308728
rect 253020 308508 253072 308514
rect 253020 308450 253072 308456
rect 253308 308446 253336 310406
rect 253388 308644 253440 308650
rect 253388 308586 253440 308592
rect 253296 308440 253348 308446
rect 252940 308366 253060 308394
rect 253296 308382 253348 308388
rect 252848 308230 252968 308258
rect 252836 308168 252888 308174
rect 252836 308110 252888 308116
rect 252848 287842 252876 308110
rect 252940 293282 252968 308230
rect 252928 293276 252980 293282
rect 252928 293218 252980 293224
rect 252836 287836 252888 287842
rect 252836 287778 252888 287784
rect 252744 287768 252796 287774
rect 252744 287710 252796 287716
rect 252652 283824 252704 283830
rect 252652 283766 252704 283772
rect 253032 282402 253060 308366
rect 253204 307896 253256 307902
rect 253204 307838 253256 307844
rect 253020 282396 253072 282402
rect 253020 282338 253072 282344
rect 251640 250776 251692 250782
rect 251640 250718 251692 250724
rect 247132 250708 247184 250714
rect 247132 250650 247184 250656
rect 247040 250640 247092 250646
rect 247040 250582 247092 250588
rect 245752 250572 245804 250578
rect 245752 250514 245804 250520
rect 245660 247784 245712 247790
rect 245660 247726 245712 247732
rect 242992 246492 243044 246498
rect 242992 246434 243044 246440
rect 242900 246424 242952 246430
rect 242900 246366 242952 246372
rect 241520 246356 241572 246362
rect 241520 246298 241572 246304
rect 253216 245206 253244 307838
rect 253400 296714 253428 308586
rect 253676 308174 253704 310420
rect 253664 308168 253716 308174
rect 253664 308110 253716 308116
rect 253952 305386 253980 310420
rect 254150 310406 254348 310434
rect 254320 307018 254348 310406
rect 254308 307012 254360 307018
rect 254308 306954 254360 306960
rect 254412 306490 254440 310420
rect 254596 308922 254624 310420
rect 254688 310406 254886 310434
rect 254584 308916 254636 308922
rect 254584 308858 254636 308864
rect 254492 307012 254544 307018
rect 254492 306954 254544 306960
rect 254032 306468 254084 306474
rect 254032 306410 254084 306416
rect 254136 306462 254440 306490
rect 253940 305380 253992 305386
rect 253940 305322 253992 305328
rect 253308 296686 253428 296714
rect 253308 263158 253336 296686
rect 254044 285258 254072 306410
rect 254136 287910 254164 306462
rect 254216 306400 254268 306406
rect 254216 306342 254268 306348
rect 254228 289202 254256 306342
rect 254308 305380 254360 305386
rect 254308 305322 254360 305328
rect 254320 293350 254348 305322
rect 254504 299474 254532 306954
rect 254688 306474 254716 310406
rect 254676 306468 254728 306474
rect 254676 306410 254728 306416
rect 255056 306406 255084 310420
rect 255044 306400 255096 306406
rect 255044 306342 255096 306348
rect 255332 304162 255360 310420
rect 255412 306468 255464 306474
rect 255412 306410 255464 306416
rect 255320 304156 255372 304162
rect 255320 304098 255372 304104
rect 254412 299446 254532 299474
rect 254308 293344 254360 293350
rect 254308 293286 254360 293292
rect 254216 289196 254268 289202
rect 254216 289138 254268 289144
rect 254124 287904 254176 287910
rect 254124 287846 254176 287852
rect 254032 285252 254084 285258
rect 254032 285194 254084 285200
rect 254412 283898 254440 299446
rect 254400 283892 254452 283898
rect 254400 283834 254452 283840
rect 253296 263152 253348 263158
rect 253296 263094 253348 263100
rect 255424 252142 255452 306410
rect 255516 306406 255544 310420
rect 255608 310406 255806 310434
rect 255504 306400 255556 306406
rect 255504 306342 255556 306348
rect 255504 305380 255556 305386
rect 255504 305322 255556 305328
rect 255516 289338 255544 305322
rect 255504 289332 255556 289338
rect 255504 289274 255556 289280
rect 255608 289270 255636 310406
rect 255976 308990 256004 310420
rect 256068 310406 256266 310434
rect 255964 308984 256016 308990
rect 255964 308926 256016 308932
rect 256068 306474 256096 310406
rect 256056 306468 256108 306474
rect 256056 306410 256108 306416
rect 255780 306400 255832 306406
rect 255780 306342 255832 306348
rect 255688 304156 255740 304162
rect 255688 304098 255740 304104
rect 255700 293418 255728 304098
rect 255688 293412 255740 293418
rect 255688 293354 255740 293360
rect 255596 289264 255648 289270
rect 255596 289206 255648 289212
rect 255412 252136 255464 252142
rect 255412 252078 255464 252084
rect 255792 252074 255820 306342
rect 256436 305386 256464 310420
rect 256424 305380 256476 305386
rect 256424 305322 256476 305328
rect 256712 294642 256740 310420
rect 256792 307964 256844 307970
rect 256792 307906 256844 307912
rect 256700 294636 256752 294642
rect 256700 294578 256752 294584
rect 255780 252068 255832 252074
rect 255780 252010 255832 252016
rect 256804 247858 256832 307906
rect 256896 260302 256924 310420
rect 257080 310406 257186 310434
rect 256976 306468 257028 306474
rect 256976 306410 257028 306416
rect 256988 261594 257016 306410
rect 257080 264314 257108 310406
rect 257356 307970 257384 310420
rect 257448 310406 257646 310434
rect 257344 307964 257396 307970
rect 257344 307906 257396 307912
rect 257344 307828 257396 307834
rect 257344 307770 257396 307776
rect 257160 306400 257212 306406
rect 257160 306342 257212 306348
rect 257068 264308 257120 264314
rect 257068 264250 257120 264256
rect 256976 261588 257028 261594
rect 256976 261530 257028 261536
rect 256884 260296 256936 260302
rect 256884 260238 256936 260244
rect 256792 247852 256844 247858
rect 256792 247794 256844 247800
rect 257172 246566 257200 306342
rect 257160 246560 257212 246566
rect 257160 246502 257212 246508
rect 253204 245200 253256 245206
rect 253204 245142 253256 245148
rect 257356 245138 257384 307770
rect 257448 306474 257476 310406
rect 257436 306468 257488 306474
rect 257436 306410 257488 306416
rect 257816 306406 257844 310420
rect 257804 306400 257856 306406
rect 257804 306342 257856 306348
rect 258092 303754 258120 310420
rect 258276 307834 258304 310420
rect 258460 310406 258566 310434
rect 258264 307828 258316 307834
rect 258264 307770 258316 307776
rect 258460 306218 258488 310406
rect 258184 306190 258488 306218
rect 258080 303748 258132 303754
rect 258080 303690 258132 303696
rect 258184 265742 258212 306190
rect 258264 305380 258316 305386
rect 258264 305322 258316 305328
rect 258276 268462 258304 305322
rect 258356 303748 258408 303754
rect 258356 303690 258408 303696
rect 258368 272610 258396 303690
rect 258736 296714 258764 310420
rect 259012 307902 259040 310420
rect 259000 307896 259052 307902
rect 259000 307838 259052 307844
rect 259196 305386 259224 310420
rect 259472 306474 259500 310420
rect 259460 306468 259512 306474
rect 259460 306410 259512 306416
rect 259656 306354 259684 310420
rect 259472 306326 259684 306354
rect 259748 310406 259946 310434
rect 259184 305380 259236 305386
rect 259184 305322 259236 305328
rect 258460 296686 258764 296714
rect 258356 272604 258408 272610
rect 258356 272546 258408 272552
rect 258264 268456 258316 268462
rect 258264 268398 258316 268404
rect 258172 265736 258224 265742
rect 258172 265678 258224 265684
rect 258460 249150 258488 296686
rect 259472 262954 259500 306326
rect 259748 306218 259776 310406
rect 259828 306468 259880 306474
rect 259828 306410 259880 306416
rect 259656 306190 259776 306218
rect 259552 305312 259604 305318
rect 259552 305254 259604 305260
rect 259564 264382 259592 305254
rect 259656 269958 259684 306190
rect 259736 305380 259788 305386
rect 259736 305322 259788 305328
rect 259748 271318 259776 305322
rect 259840 274038 259868 306410
rect 260116 302234 260144 310420
rect 260208 310406 260406 310434
rect 260208 305318 260236 310406
rect 260288 307828 260340 307834
rect 260288 307770 260340 307776
rect 260196 305312 260248 305318
rect 260196 305254 260248 305260
rect 259932 302206 260144 302234
rect 259932 276758 259960 302206
rect 260300 296714 260328 307770
rect 260576 305386 260604 310420
rect 260852 306474 260880 310420
rect 261036 307018 261064 310420
rect 261024 307012 261076 307018
rect 261024 306954 261076 306960
rect 261024 306808 261076 306814
rect 261024 306750 261076 306756
rect 260840 306468 260892 306474
rect 260840 306410 260892 306416
rect 260564 305380 260616 305386
rect 260564 305322 260616 305328
rect 260840 305380 260892 305386
rect 260840 305322 260892 305328
rect 260116 296686 260328 296714
rect 259920 276752 259972 276758
rect 259920 276694 259972 276700
rect 259828 274032 259880 274038
rect 259828 273974 259880 273980
rect 259736 271312 259788 271318
rect 259736 271254 259788 271260
rect 259644 269952 259696 269958
rect 259644 269894 259696 269900
rect 260116 267238 260144 296686
rect 260104 267232 260156 267238
rect 260104 267174 260156 267180
rect 259552 264376 259604 264382
rect 259552 264318 259604 264324
rect 259460 262948 259512 262954
rect 259460 262890 259512 262896
rect 258448 249144 258500 249150
rect 258448 249086 258500 249092
rect 260852 247926 260880 305322
rect 260932 305312 260984 305318
rect 260932 305254 260984 305260
rect 260944 247994 260972 305254
rect 261036 265810 261064 306750
rect 261208 306468 261260 306474
rect 261208 306410 261260 306416
rect 261116 306400 261168 306406
rect 261116 306342 261168 306348
rect 261128 267170 261156 306342
rect 261220 278118 261248 306410
rect 261312 305386 261340 310420
rect 261300 305380 261352 305386
rect 261300 305322 261352 305328
rect 261496 296714 261524 310420
rect 261588 310406 261786 310434
rect 261588 306406 261616 310406
rect 261576 306400 261628 306406
rect 261576 306342 261628 306348
rect 261956 305318 261984 310420
rect 262232 305386 262260 310420
rect 262416 307834 262444 310420
rect 262508 310406 262706 310434
rect 262404 307828 262456 307834
rect 262404 307770 262456 307776
rect 262508 306490 262536 310406
rect 262324 306462 262536 306490
rect 262220 305380 262272 305386
rect 262220 305322 262272 305328
rect 261944 305312 261996 305318
rect 261944 305254 261996 305260
rect 261312 296686 261524 296714
rect 261312 279614 261340 296686
rect 261300 279608 261352 279614
rect 261300 279550 261352 279556
rect 261208 278112 261260 278118
rect 261208 278054 261260 278060
rect 262324 272678 262352 306462
rect 262404 306400 262456 306406
rect 262876 306354 262904 310420
rect 262404 306342 262456 306348
rect 262416 274106 262444 306342
rect 262508 306326 262904 306354
rect 262968 310406 263166 310434
rect 262508 281042 262536 306326
rect 262588 305380 262640 305386
rect 262588 305322 262640 305328
rect 262496 281036 262548 281042
rect 262496 280978 262548 280984
rect 262600 280974 262628 305322
rect 262968 296714 262996 310406
rect 263336 306406 263364 310420
rect 263612 308530 263640 310420
rect 263520 308502 263640 308530
rect 263520 308242 263548 308502
rect 263796 308394 263824 310420
rect 263612 308366 263824 308394
rect 263888 310406 264086 310434
rect 263508 308236 263560 308242
rect 263508 308178 263560 308184
rect 263324 306400 263376 306406
rect 263324 306342 263376 306348
rect 262692 296686 262996 296714
rect 262588 280968 262640 280974
rect 262588 280910 262640 280916
rect 262404 274100 262456 274106
rect 262404 274042 262456 274048
rect 262312 272672 262364 272678
rect 262312 272614 262364 272620
rect 262692 268530 262720 296686
rect 262680 268524 262732 268530
rect 262680 268466 262732 268472
rect 261116 267164 261168 267170
rect 261116 267106 261168 267112
rect 261024 265804 261076 265810
rect 261024 265746 261076 265752
rect 263612 260370 263640 308366
rect 263692 308168 263744 308174
rect 263692 308110 263744 308116
rect 263704 261662 263732 308110
rect 263784 308032 263836 308038
rect 263784 307974 263836 307980
rect 263796 268666 263824 307974
rect 263784 268660 263836 268666
rect 263784 268602 263836 268608
rect 263888 268598 263916 310406
rect 264256 308394 264284 310420
rect 263980 308366 264284 308394
rect 264348 310406 264546 310434
rect 263980 275398 264008 308366
rect 264060 308236 264112 308242
rect 264060 308178 264112 308184
rect 264072 282470 264100 308178
rect 264348 308174 264376 310406
rect 264336 308168 264388 308174
rect 264336 308110 264388 308116
rect 264716 308038 264744 310420
rect 264992 308446 265020 310420
rect 264980 308440 265032 308446
rect 265176 308394 265204 310420
rect 264980 308382 265032 308388
rect 265084 308366 265204 308394
rect 265268 310406 265466 310434
rect 265544 310406 265742 310434
rect 264704 308032 264756 308038
rect 264704 307974 264756 307980
rect 264980 307284 265032 307290
rect 264980 307226 265032 307232
rect 264060 282464 264112 282470
rect 264060 282406 264112 282412
rect 263968 275392 264020 275398
rect 263968 275334 264020 275340
rect 263876 268592 263928 268598
rect 263876 268534 263928 268540
rect 264992 261798 265020 307226
rect 264980 261792 265032 261798
rect 264980 261734 265032 261740
rect 265084 261730 265112 308366
rect 265268 308258 265296 310406
rect 265348 308440 265400 308446
rect 265348 308382 265400 308388
rect 265176 308230 265296 308258
rect 265176 270026 265204 308230
rect 265256 308168 265308 308174
rect 265256 308110 265308 308116
rect 265268 270094 265296 308110
rect 265360 275466 265388 308382
rect 265544 296714 265572 310406
rect 265912 307290 265940 310420
rect 266004 310406 266202 310434
rect 266386 310406 266584 310434
rect 266004 308174 266032 310406
rect 266452 308440 266504 308446
rect 266452 308382 266504 308388
rect 266556 308394 266584 310406
rect 266648 308718 266676 310420
rect 266636 308712 266688 308718
rect 266636 308654 266688 308660
rect 266832 308446 266860 310420
rect 266924 310406 267122 310434
rect 266820 308440 266872 308446
rect 265992 308168 266044 308174
rect 265992 308110 266044 308116
rect 265900 307284 265952 307290
rect 265900 307226 265952 307232
rect 265452 296686 265572 296714
rect 265452 276826 265480 296686
rect 265440 276820 265492 276826
rect 265440 276762 265492 276768
rect 265348 275460 265400 275466
rect 265348 275402 265400 275408
rect 266464 270162 266492 308382
rect 266556 308366 266768 308394
rect 266820 308382 266872 308388
rect 266544 308236 266596 308242
rect 266544 308178 266596 308184
rect 266556 271386 266584 308178
rect 266636 307556 266688 307562
rect 266636 307498 266688 307504
rect 266648 276962 266676 307498
rect 266636 276956 266688 276962
rect 266636 276898 266688 276904
rect 266740 276894 266768 308366
rect 266924 307562 266952 310406
rect 266912 307556 266964 307562
rect 266912 307498 266964 307504
rect 267292 296714 267320 310420
rect 267384 310406 267582 310434
rect 267384 308242 267412 310406
rect 267372 308236 267424 308242
rect 267372 308178 267424 308184
rect 267752 308038 267780 310420
rect 267844 310406 268042 310434
rect 267740 308032 267792 308038
rect 267740 307974 267792 307980
rect 267740 307692 267792 307698
rect 267740 307634 267792 307640
rect 266832 296686 267320 296714
rect 266728 276888 266780 276894
rect 266728 276830 266780 276836
rect 266544 271380 266596 271386
rect 266544 271322 266596 271328
rect 266452 270156 266504 270162
rect 266452 270098 266504 270104
rect 265256 270088 265308 270094
rect 265256 270030 265308 270036
rect 265164 270020 265216 270026
rect 265164 269962 265216 269968
rect 266832 261866 266860 296686
rect 267752 263090 267780 307634
rect 267740 263084 267792 263090
rect 267740 263026 267792 263032
rect 267844 263022 267872 310406
rect 268212 308394 268240 310420
rect 267936 308366 268240 308394
rect 268304 310406 268502 310434
rect 267936 271454 267964 308366
rect 268016 308236 268068 308242
rect 268016 308178 268068 308184
rect 268028 271522 268056 308178
rect 268108 308032 268160 308038
rect 268108 307974 268160 307980
rect 268120 278186 268148 307974
rect 268304 296714 268332 310406
rect 268672 307698 268700 310420
rect 268764 310406 268962 310434
rect 269146 310406 269344 310434
rect 268764 308242 268792 310406
rect 269212 308440 269264 308446
rect 269212 308382 269264 308388
rect 269316 308394 269344 310406
rect 269408 308530 269436 310420
rect 269408 308502 269528 308530
rect 268752 308236 268804 308242
rect 268752 308178 268804 308184
rect 268660 307692 268712 307698
rect 268660 307634 268712 307640
rect 268212 296686 268332 296714
rect 268212 278254 268240 296686
rect 268200 278248 268252 278254
rect 268200 278190 268252 278196
rect 268108 278180 268160 278186
rect 268108 278122 268160 278128
rect 268016 271516 268068 271522
rect 268016 271458 268068 271464
rect 267924 271448 267976 271454
rect 267924 271390 267976 271396
rect 269224 264450 269252 308382
rect 269316 308366 269436 308394
rect 269304 308236 269356 308242
rect 269304 308178 269356 308184
rect 269316 272746 269344 308178
rect 269408 278322 269436 308366
rect 269500 307154 269528 308502
rect 269592 307154 269620 310420
rect 269684 310406 269882 310434
rect 269488 307148 269540 307154
rect 269488 307090 269540 307096
rect 269580 307148 269632 307154
rect 269580 307090 269632 307096
rect 269684 307034 269712 310406
rect 270052 308446 270080 310420
rect 270144 310406 270342 310434
rect 270040 308440 270092 308446
rect 270040 308382 270092 308388
rect 270144 308242 270172 310406
rect 270512 308242 270540 310420
rect 270604 310406 270802 310434
rect 270132 308236 270184 308242
rect 270132 308178 270184 308184
rect 270500 308236 270552 308242
rect 270500 308178 270552 308184
rect 270500 308100 270552 308106
rect 270500 308042 270552 308048
rect 269500 307006 269712 307034
rect 269500 279682 269528 307006
rect 269580 306944 269632 306950
rect 269580 306886 269632 306892
rect 269488 279676 269540 279682
rect 269488 279618 269540 279624
rect 269396 278316 269448 278322
rect 269396 278258 269448 278264
rect 269304 272740 269356 272746
rect 269304 272682 269356 272688
rect 269212 264444 269264 264450
rect 269212 264386 269264 264392
rect 267832 263016 267884 263022
rect 267832 262958 267884 262964
rect 266820 261860 266872 261866
rect 266820 261802 266872 261808
rect 265072 261724 265124 261730
rect 265072 261666 265124 261672
rect 263692 261656 263744 261662
rect 263692 261598 263744 261604
rect 263600 260364 263652 260370
rect 263600 260306 263652 260312
rect 260932 247988 260984 247994
rect 260932 247930 260984 247936
rect 260840 247920 260892 247926
rect 260840 247862 260892 247868
rect 269592 246634 269620 306886
rect 270512 262857 270540 308042
rect 270604 264518 270632 310406
rect 270972 308530 271000 310420
rect 270788 308502 271000 308530
rect 271064 310406 271262 310434
rect 270684 308440 270736 308446
rect 270684 308382 270736 308388
rect 270696 272882 270724 308382
rect 270684 272876 270736 272882
rect 270684 272818 270736 272824
rect 270788 272814 270816 308502
rect 271064 308394 271092 310406
rect 270880 308366 271092 308394
rect 270880 279818 270908 308366
rect 270960 308236 271012 308242
rect 270960 308178 271012 308184
rect 270868 279812 270920 279818
rect 270868 279754 270920 279760
rect 270972 279750 271000 308178
rect 271432 308106 271460 310420
rect 271524 310406 271722 310434
rect 271906 310406 272104 310434
rect 271524 308446 271552 310406
rect 271880 308508 271932 308514
rect 271880 308450 271932 308456
rect 271512 308440 271564 308446
rect 271512 308382 271564 308388
rect 271420 308100 271472 308106
rect 271420 308042 271472 308048
rect 271892 307222 271920 308450
rect 271972 308440 272024 308446
rect 271972 308382 272024 308388
rect 271880 307216 271932 307222
rect 271880 307158 271932 307164
rect 270960 279744 271012 279750
rect 270960 279686 271012 279692
rect 270776 272808 270828 272814
rect 270776 272750 270828 272756
rect 271984 264586 272012 308382
rect 272076 307154 272104 310406
rect 272168 308514 272196 310420
rect 272156 308508 272208 308514
rect 272156 308450 272208 308456
rect 272352 308394 272380 310420
rect 272168 308366 272380 308394
rect 272444 310406 272642 310434
rect 272064 307148 272116 307154
rect 272064 307090 272116 307096
rect 272064 307012 272116 307018
rect 272064 306954 272116 306960
rect 272076 274310 272104 306954
rect 272064 274304 272116 274310
rect 272064 274246 272116 274252
rect 272168 274174 272196 308366
rect 272248 307148 272300 307154
rect 272248 307090 272300 307096
rect 272260 281110 272288 307090
rect 272444 296714 272472 310406
rect 272812 308446 272840 310420
rect 272904 310406 273102 310434
rect 272800 308440 272852 308446
rect 272800 308382 272852 308388
rect 272904 307018 272932 310406
rect 272892 307012 272944 307018
rect 272892 306954 272944 306960
rect 273076 306468 273128 306474
rect 273076 306410 273128 306416
rect 273088 306270 273116 306410
rect 273076 306264 273128 306270
rect 273076 306206 273128 306212
rect 272352 296686 272472 296714
rect 272248 281104 272300 281110
rect 272248 281046 272300 281052
rect 272156 274168 272208 274174
rect 272156 274110 272208 274116
rect 271972 264580 272024 264586
rect 271972 264522 272024 264528
rect 270592 264512 270644 264518
rect 270592 264454 270644 264460
rect 270498 262848 270554 262857
rect 270498 262783 270554 262792
rect 272352 249218 272380 296686
rect 273272 249286 273300 310420
rect 273456 310406 273562 310434
rect 273352 306400 273404 306406
rect 273352 306342 273404 306348
rect 273260 249280 273312 249286
rect 273260 249222 273312 249228
rect 272340 249212 272392 249218
rect 272340 249154 272392 249160
rect 273364 249121 273392 306342
rect 273456 265878 273484 310406
rect 273536 306332 273588 306338
rect 273536 306274 273588 306280
rect 273444 265872 273496 265878
rect 273444 265814 273496 265820
rect 273548 265577 273576 306274
rect 273732 302234 273760 310420
rect 273824 310406 274022 310434
rect 273824 306406 273852 310406
rect 273812 306400 273864 306406
rect 273812 306342 273864 306348
rect 274192 306338 274220 310420
rect 274284 310406 274482 310434
rect 274180 306332 274232 306338
rect 274180 306274 274232 306280
rect 273640 302206 273760 302234
rect 273640 274242 273668 302206
rect 274284 296714 274312 310406
rect 274652 307057 274680 310420
rect 274638 307048 274694 307057
rect 274638 306983 274694 306992
rect 274928 306241 274956 310420
rect 274914 306232 274970 306241
rect 274914 306167 274970 306176
rect 275112 302234 275140 310420
rect 275388 306105 275416 310420
rect 275572 308961 275600 310420
rect 275558 308952 275614 308961
rect 275558 308887 275614 308896
rect 275374 306096 275430 306105
rect 275374 306031 275430 306040
rect 275848 305969 275876 310420
rect 275834 305960 275890 305969
rect 275834 305895 275890 305904
rect 276032 305833 276060 310420
rect 276308 308174 276336 310420
rect 276296 308168 276348 308174
rect 276296 308110 276348 308116
rect 276018 305824 276074 305833
rect 276018 305759 276074 305768
rect 276492 305590 276520 310420
rect 276480 305584 276532 305590
rect 276480 305526 276532 305532
rect 276768 303385 276796 310420
rect 276952 308825 276980 310420
rect 276938 308816 276994 308825
rect 276938 308751 276994 308760
rect 277228 305454 277256 310420
rect 277216 305448 277268 305454
rect 277216 305390 277268 305396
rect 276754 303376 276810 303385
rect 276754 303311 276810 303320
rect 277412 303113 277440 310420
rect 277688 308310 277716 310420
rect 277676 308304 277728 308310
rect 277676 308246 277728 308252
rect 277872 306202 277900 310420
rect 277860 306196 277912 306202
rect 277860 306138 277912 306144
rect 278148 303249 278176 310420
rect 278332 308689 278360 310420
rect 278318 308680 278374 308689
rect 278318 308615 278374 308624
rect 278608 305522 278636 310420
rect 278596 305516 278648 305522
rect 278596 305458 278648 305464
rect 278134 303240 278190 303249
rect 278134 303175 278190 303184
rect 277398 303104 277454 303113
rect 277398 303039 277454 303048
rect 278792 302841 278820 310420
rect 279068 308378 279096 310420
rect 279056 308372 279108 308378
rect 279056 308314 279108 308320
rect 279252 306066 279280 310420
rect 279240 306060 279292 306066
rect 279240 306002 279292 306008
rect 279528 302977 279556 310420
rect 279712 309126 279740 310420
rect 279700 309120 279752 309126
rect 279700 309062 279752 309068
rect 279988 306542 280016 310420
rect 279976 306536 280028 306542
rect 279976 306478 280028 306484
rect 280172 303618 280200 310420
rect 280448 309058 280476 310420
rect 280436 309052 280488 309058
rect 280436 308994 280488 309000
rect 280632 305998 280660 310420
rect 280620 305992 280672 305998
rect 280620 305934 280672 305940
rect 280160 303612 280212 303618
rect 280160 303554 280212 303560
rect 279514 302968 279570 302977
rect 279514 302903 279570 302912
rect 278778 302832 278834 302841
rect 280908 302802 280936 310420
rect 280988 306468 281040 306474
rect 280988 306410 281040 306416
rect 278778 302767 278834 302776
rect 280896 302796 280948 302802
rect 280896 302738 280948 302744
rect 273732 296686 274312 296714
rect 274652 302206 275140 302234
rect 273732 275233 273760 296686
rect 273718 275224 273774 275233
rect 273718 275159 273774 275168
rect 273628 274236 273680 274242
rect 273628 274178 273680 274184
rect 273534 265568 273590 265577
rect 273534 265503 273590 265512
rect 273350 249112 273406 249121
rect 273350 249047 273406 249056
rect 269580 246628 269632 246634
rect 269580 246570 269632 246576
rect 274652 246265 274680 302206
rect 281000 300626 281028 306410
rect 281092 306134 281120 310420
rect 281080 306128 281132 306134
rect 281080 306070 281132 306076
rect 281368 305697 281396 310420
rect 281354 305688 281410 305697
rect 281354 305623 281410 305632
rect 281552 302734 281580 310420
rect 281828 306338 281856 310420
rect 281816 306332 281868 306338
rect 281816 306274 281868 306280
rect 282104 303550 282132 310420
rect 282092 303544 282144 303550
rect 282092 303486 282144 303492
rect 282288 303278 282316 310420
rect 282564 303482 282592 310420
rect 282748 305930 282776 310420
rect 282736 305924 282788 305930
rect 282736 305866 282788 305872
rect 282552 303476 282604 303482
rect 282552 303418 282604 303424
rect 282276 303272 282328 303278
rect 282276 303214 282328 303220
rect 283024 303210 283052 310420
rect 283208 305402 283236 310420
rect 283484 305862 283512 310420
rect 283472 305856 283524 305862
rect 283472 305798 283524 305804
rect 283116 305374 283236 305402
rect 283116 303346 283144 305374
rect 283668 305266 283696 310420
rect 283208 305238 283696 305266
rect 283104 303340 283156 303346
rect 283104 303282 283156 303288
rect 283012 303204 283064 303210
rect 283012 303146 283064 303152
rect 281540 302728 281592 302734
rect 281540 302670 281592 302676
rect 280988 300620 281040 300626
rect 280988 300562 281040 300568
rect 283208 300121 283236 305238
rect 283944 302870 283972 310420
rect 283932 302864 283984 302870
rect 283932 302806 283984 302812
rect 284128 302234 284156 310420
rect 284300 306400 284352 306406
rect 284300 306342 284352 306348
rect 283300 302206 284156 302234
rect 283194 300112 283250 300121
rect 283194 300047 283250 300056
rect 283300 300014 283328 302206
rect 284312 300694 284340 306342
rect 284404 306270 284432 310420
rect 284588 306354 284616 310420
rect 284496 306326 284616 306354
rect 284772 310406 284878 310434
rect 284668 306332 284720 306338
rect 284392 306264 284444 306270
rect 284392 306206 284444 306212
rect 284392 306128 284444 306134
rect 284392 306070 284444 306076
rect 284300 300688 284352 300694
rect 284300 300630 284352 300636
rect 284404 300558 284432 306070
rect 284392 300552 284444 300558
rect 284392 300494 284444 300500
rect 284496 300218 284524 306326
rect 284668 306274 284720 306280
rect 284576 306264 284628 306270
rect 284576 306206 284628 306212
rect 284484 300212 284536 300218
rect 284484 300154 284536 300160
rect 283288 300008 283340 300014
rect 283288 299950 283340 299956
rect 284588 299946 284616 306206
rect 284680 300286 284708 306274
rect 284772 300490 284800 310406
rect 285048 306134 285076 310420
rect 285140 310406 285338 310434
rect 285140 306338 285168 310406
rect 285508 306406 285536 310420
rect 285784 309134 285812 310420
rect 285692 309106 285812 309134
rect 285496 306400 285548 306406
rect 285496 306342 285548 306348
rect 285128 306332 285180 306338
rect 285128 306274 285180 306280
rect 285036 306128 285088 306134
rect 285036 306070 285088 306076
rect 284760 300484 284812 300490
rect 284760 300426 284812 300432
rect 285692 300422 285720 309106
rect 285968 306474 285996 310420
rect 286152 310406 286258 310434
rect 285956 306468 286008 306474
rect 285956 306410 286008 306416
rect 286048 306332 286100 306338
rect 286048 306274 286100 306280
rect 285772 306264 285824 306270
rect 285772 306206 285824 306212
rect 285784 300762 285812 306206
rect 285864 306196 285916 306202
rect 285864 306138 285916 306144
rect 285876 300830 285904 306138
rect 285864 300824 285916 300830
rect 285864 300766 285916 300772
rect 285772 300756 285824 300762
rect 285772 300698 285824 300704
rect 285680 300416 285732 300422
rect 285680 300358 285732 300364
rect 284668 300280 284720 300286
rect 284668 300222 284720 300228
rect 284576 299940 284628 299946
rect 284576 299882 284628 299888
rect 274638 246256 274694 246265
rect 274638 246191 274694 246200
rect 257344 245132 257396 245138
rect 257344 245074 257396 245080
rect 233240 245064 233292 245070
rect 233240 245006 233292 245012
rect 232044 244996 232096 245002
rect 232044 244938 232096 244944
rect 231952 244928 232004 244934
rect 231952 244870 232004 244876
rect 286060 243710 286088 306274
rect 286152 306270 286180 310406
rect 286140 306264 286192 306270
rect 286140 306206 286192 306212
rect 286428 300082 286456 310420
rect 286520 310406 286718 310434
rect 286520 306202 286548 310406
rect 286888 306338 286916 310420
rect 286876 306332 286928 306338
rect 286876 306274 286928 306280
rect 286508 306196 286560 306202
rect 286508 306138 286560 306144
rect 287164 302234 287192 310420
rect 287348 308854 287376 310420
rect 287336 308848 287388 308854
rect 287336 308790 287388 308796
rect 287624 305726 287652 310420
rect 287612 305720 287664 305726
rect 287612 305662 287664 305668
rect 287808 302234 287836 310420
rect 288084 305794 288112 310420
rect 288072 305788 288124 305794
rect 288072 305730 288124 305736
rect 288268 303414 288296 310420
rect 288544 306542 288572 310420
rect 288532 306536 288584 306542
rect 288532 306478 288584 306484
rect 288728 306354 288756 310420
rect 288820 310406 289018 310434
rect 288820 306474 288848 310406
rect 288808 306468 288860 306474
rect 288808 306410 288860 306416
rect 288452 306326 288756 306354
rect 288256 303408 288308 303414
rect 288256 303350 288308 303356
rect 287164 302206 287376 302234
rect 286416 300076 286468 300082
rect 286416 300018 286468 300024
rect 287348 243778 287376 302206
rect 287440 302206 287836 302234
rect 287336 243772 287388 243778
rect 287336 243714 287388 243720
rect 286048 243704 286100 243710
rect 286048 243646 286100 243652
rect 287440 243574 287468 302206
rect 288452 300150 288480 306326
rect 288624 306264 288676 306270
rect 288624 306206 288676 306212
rect 288900 306264 288952 306270
rect 288900 306206 288952 306212
rect 288532 306128 288584 306134
rect 288532 306070 288584 306076
rect 288440 300144 288492 300150
rect 288440 300086 288492 300092
rect 288544 245274 288572 306070
rect 288636 245342 288664 306206
rect 288716 306196 288768 306202
rect 288716 306138 288768 306144
rect 288728 247722 288756 306138
rect 288808 306060 288860 306066
rect 288808 306002 288860 306008
rect 288820 247790 288848 306002
rect 288808 247784 288860 247790
rect 288808 247726 288860 247732
rect 288716 247716 288768 247722
rect 288716 247658 288768 247664
rect 288624 245336 288676 245342
rect 288624 245278 288676 245284
rect 288532 245268 288584 245274
rect 288532 245210 288584 245216
rect 288912 243642 288940 306206
rect 289188 306134 289216 310420
rect 289280 310406 289478 310434
rect 289176 306128 289228 306134
rect 289176 306070 289228 306076
rect 289280 306066 289308 310406
rect 289648 306202 289676 310420
rect 289924 308242 289952 310420
rect 289912 308236 289964 308242
rect 289912 308178 289964 308184
rect 289820 306400 289872 306406
rect 289820 306342 289872 306348
rect 289636 306196 289688 306202
rect 289636 306138 289688 306144
rect 289268 306060 289320 306066
rect 289268 306002 289320 306008
rect 289832 243710 289860 306342
rect 289912 306332 289964 306338
rect 289912 306274 289964 306280
rect 289820 243704 289872 243710
rect 289820 243646 289872 243652
rect 289924 243642 289952 306274
rect 290108 296714 290136 310420
rect 290200 310406 290398 310434
rect 290200 306338 290228 310406
rect 290568 308582 290596 310420
rect 290556 308576 290608 308582
rect 290556 308518 290608 308524
rect 290844 308514 290872 310420
rect 290832 308508 290884 308514
rect 290832 308450 290884 308456
rect 291028 306406 291056 310420
rect 291304 308718 291332 310420
rect 291292 308712 291344 308718
rect 291292 308654 291344 308660
rect 291488 306490 291516 310420
rect 291212 306462 291516 306490
rect 291580 310406 291778 310434
rect 291016 306400 291068 306406
rect 291016 306342 291068 306348
rect 290188 306332 290240 306338
rect 290188 306274 290240 306280
rect 290016 296686 290136 296714
rect 290016 243778 290044 296686
rect 290004 243772 290056 243778
rect 290004 243714 290056 243720
rect 288900 243636 288952 243642
rect 288900 243578 288952 243584
rect 289912 243636 289964 243642
rect 289912 243578 289964 243584
rect 291212 243574 291240 306462
rect 291580 306354 291608 310406
rect 291292 306332 291344 306338
rect 291292 306274 291344 306280
rect 291396 306326 291608 306354
rect 291948 306338 291976 310420
rect 292040 310406 292238 310434
rect 291936 306332 291988 306338
rect 291304 245206 291332 306274
rect 291396 246702 291424 306326
rect 291936 306274 291988 306280
rect 291476 306264 291528 306270
rect 291476 306206 291528 306212
rect 291488 247586 291516 306206
rect 292040 296714 292068 310406
rect 292408 306270 292436 310420
rect 292684 308650 292712 310420
rect 292672 308644 292724 308650
rect 292672 308586 292724 308592
rect 292868 306490 292896 310420
rect 292592 306462 292896 306490
rect 292960 310406 293158 310434
rect 292960 306474 292988 310406
rect 292948 306468 293000 306474
rect 292396 306264 292448 306270
rect 292396 306206 292448 306212
rect 291580 296686 292068 296714
rect 291580 250646 291608 296686
rect 291568 250640 291620 250646
rect 291568 250582 291620 250588
rect 291476 247580 291528 247586
rect 291476 247522 291528 247528
rect 291384 246696 291436 246702
rect 291384 246638 291436 246644
rect 292592 245274 292620 306462
rect 292948 306410 293000 306416
rect 292672 306400 292724 306406
rect 293328 306354 293356 310420
rect 292672 306342 292724 306348
rect 292684 248198 292712 306342
rect 292776 306326 293356 306354
rect 293420 310406 293618 310434
rect 292672 248192 292724 248198
rect 292672 248134 292724 248140
rect 292776 247994 292804 306326
rect 292856 306264 292908 306270
rect 292856 306206 292908 306212
rect 292764 247988 292816 247994
rect 292764 247930 292816 247936
rect 292868 247926 292896 306206
rect 293420 296714 293448 310406
rect 293788 306270 293816 310420
rect 293960 306332 294012 306338
rect 294064 306320 294092 310420
rect 294248 308854 294276 310420
rect 294236 308848 294288 308854
rect 294236 308790 294288 308796
rect 294524 308786 294552 310420
rect 294512 308780 294564 308786
rect 294512 308722 294564 308728
rect 294064 306292 294184 306320
rect 293960 306274 294012 306280
rect 293776 306264 293828 306270
rect 293776 306206 293828 306212
rect 292960 296686 293448 296714
rect 292960 251054 292988 296686
rect 292948 251048 293000 251054
rect 292948 250990 293000 250996
rect 292856 247920 292908 247926
rect 292856 247862 292908 247868
rect 293972 247858 294000 306274
rect 294052 306196 294104 306202
rect 294052 306138 294104 306144
rect 294064 250714 294092 306138
rect 294156 250782 294184 306292
rect 294708 306202 294736 310420
rect 294984 308922 295012 310420
rect 294972 308916 295024 308922
rect 294972 308858 295024 308864
rect 295168 306338 295196 310420
rect 295352 310406 295458 310434
rect 295156 306332 295208 306338
rect 295156 306274 295208 306280
rect 294696 306196 294748 306202
rect 294696 306138 294748 306144
rect 295352 306134 295380 310406
rect 295628 306320 295656 310420
rect 295444 306292 295656 306320
rect 295720 310406 295918 310434
rect 295340 306128 295392 306134
rect 295340 306070 295392 306076
rect 295340 305992 295392 305998
rect 295340 305934 295392 305940
rect 294144 250776 294196 250782
rect 294144 250718 294196 250724
rect 294052 250708 294104 250714
rect 294052 250650 294104 250656
rect 293960 247852 294012 247858
rect 293960 247794 294012 247800
rect 295352 245342 295380 305934
rect 295340 245336 295392 245342
rect 295340 245278 295392 245284
rect 292580 245268 292632 245274
rect 292580 245210 292632 245216
rect 291292 245200 291344 245206
rect 291292 245142 291344 245148
rect 295444 245041 295472 306292
rect 295720 306252 295748 310406
rect 295536 306224 295748 306252
rect 295536 248169 295564 306224
rect 295708 306128 295760 306134
rect 295708 306070 295760 306076
rect 295616 306060 295668 306066
rect 295616 306002 295668 306008
rect 295628 248402 295656 306002
rect 295720 250306 295748 306070
rect 296088 296714 296116 310420
rect 296180 310406 296378 310434
rect 296180 305998 296208 310406
rect 296548 306066 296576 310420
rect 296824 306542 296852 310420
rect 296812 306536 296864 306542
rect 296812 306478 296864 306484
rect 297008 306388 297036 310420
rect 296732 306360 297036 306388
rect 297100 310406 297298 310434
rect 296536 306060 296588 306066
rect 296536 306002 296588 306008
rect 296168 305992 296220 305998
rect 296168 305934 296220 305940
rect 295812 296686 296116 296714
rect 295812 250374 295840 296686
rect 295800 250368 295852 250374
rect 295800 250310 295852 250316
rect 295708 250300 295760 250306
rect 295708 250242 295760 250248
rect 295616 248396 295668 248402
rect 295616 248338 295668 248344
rect 295522 248160 295578 248169
rect 295522 248095 295578 248104
rect 296732 245177 296760 306360
rect 297100 306320 297128 310406
rect 297180 306536 297232 306542
rect 297180 306478 297232 306484
rect 297008 306292 297128 306320
rect 296904 306264 296956 306270
rect 296904 306206 296956 306212
rect 296812 306196 296864 306202
rect 296812 306138 296864 306144
rect 296824 248062 296852 306138
rect 296812 248056 296864 248062
rect 296812 247998 296864 248004
rect 296718 245168 296774 245177
rect 296718 245103 296774 245112
rect 295430 245032 295486 245041
rect 295430 244967 295486 244976
rect 296916 244905 296944 306206
rect 297008 248130 297036 306292
rect 297192 302234 297220 306478
rect 297100 302206 297220 302234
rect 297100 248334 297128 302206
rect 297468 296714 297496 310420
rect 297560 310406 297758 310434
rect 297560 306270 297588 310406
rect 297548 306264 297600 306270
rect 297548 306206 297600 306212
rect 297928 306202 297956 310420
rect 298218 310406 298416 310434
rect 298100 306400 298152 306406
rect 298100 306342 298152 306348
rect 297916 306196 297968 306202
rect 297916 306138 297968 306144
rect 297192 296686 297496 296714
rect 297192 250850 297220 296686
rect 297180 250844 297232 250850
rect 297180 250786 297232 250792
rect 297088 248328 297140 248334
rect 297088 248270 297140 248276
rect 298112 248266 298140 306342
rect 298284 306332 298336 306338
rect 298284 306274 298336 306280
rect 298192 306264 298244 306270
rect 298192 306206 298244 306212
rect 298100 248260 298152 248266
rect 298100 248202 298152 248208
rect 296996 248124 297048 248130
rect 296996 248066 297048 248072
rect 298204 247654 298232 306206
rect 298296 250986 298324 306274
rect 298284 250980 298336 250986
rect 298284 250922 298336 250928
rect 298388 250918 298416 310406
rect 298480 308553 298508 310420
rect 298466 308544 298522 308553
rect 298466 308479 298522 308488
rect 298664 306406 298692 310420
rect 298756 310406 298954 310434
rect 298652 306400 298704 306406
rect 298652 306342 298704 306348
rect 298756 306338 298784 310406
rect 299124 308417 299152 310420
rect 299216 310406 299414 310434
rect 299110 308408 299166 308417
rect 299110 308343 299166 308352
rect 298744 306332 298796 306338
rect 298744 306274 298796 306280
rect 299216 306270 299244 310406
rect 299584 306610 299612 310420
rect 299676 310406 299874 310434
rect 299572 306604 299624 306610
rect 299572 306546 299624 306552
rect 299676 306490 299704 310406
rect 299492 306462 299704 306490
rect 299204 306264 299256 306270
rect 299204 306206 299256 306212
rect 298376 250912 298428 250918
rect 298376 250854 298428 250860
rect 298192 247648 298244 247654
rect 298192 247590 298244 247596
rect 299492 245449 299520 306462
rect 300044 306354 300072 310420
rect 299572 306332 299624 306338
rect 299572 306274 299624 306280
rect 299676 306326 300072 306354
rect 300136 310406 300334 310434
rect 299478 245440 299534 245449
rect 299584 245410 299612 306274
rect 299676 247518 299704 306326
rect 300136 306252 300164 310406
rect 300216 306604 300268 306610
rect 300216 306546 300268 306552
rect 299768 306224 300164 306252
rect 299768 251190 299796 306224
rect 299848 306128 299900 306134
rect 299848 306070 299900 306076
rect 299756 251184 299808 251190
rect 299756 251126 299808 251132
rect 299860 250442 299888 306070
rect 300228 296714 300256 306546
rect 300504 306338 300532 310420
rect 300596 310406 300794 310434
rect 300978 310406 301084 310434
rect 300492 306332 300544 306338
rect 300492 306274 300544 306280
rect 300596 306134 300624 310406
rect 301056 309134 301084 310406
rect 300964 309106 301084 309134
rect 301148 310406 301254 310434
rect 300860 307012 300912 307018
rect 300860 306954 300912 306960
rect 300584 306128 300636 306134
rect 300584 306070 300636 306076
rect 299952 296686 300256 296714
rect 299952 251122 299980 296686
rect 299940 251116 299992 251122
rect 299940 251058 299992 251064
rect 299848 250436 299900 250442
rect 299848 250378 299900 250384
rect 299664 247512 299716 247518
rect 299664 247454 299716 247460
rect 299478 245375 299534 245384
rect 299572 245404 299624 245410
rect 299572 245346 299624 245352
rect 300872 245313 300900 306954
rect 300964 306898 300992 309106
rect 301148 307018 301176 310406
rect 301424 309134 301452 310420
rect 301332 309106 301452 309134
rect 301516 310406 301714 310434
rect 301136 307012 301188 307018
rect 301136 306954 301188 306960
rect 300964 306870 301084 306898
rect 300952 306332 301004 306338
rect 300952 306274 301004 306280
rect 300964 245614 300992 306274
rect 301056 304366 301084 306870
rect 301332 304450 301360 309106
rect 301148 304422 301360 304450
rect 301044 304360 301096 304366
rect 301044 304302 301096 304308
rect 301044 303204 301096 303210
rect 301044 303146 301096 303152
rect 300952 245608 301004 245614
rect 300952 245550 301004 245556
rect 301056 245478 301084 303146
rect 301148 250753 301176 304422
rect 301228 304360 301280 304366
rect 301228 304302 301280 304308
rect 301240 253570 301268 304302
rect 301516 296714 301544 310406
rect 301884 303210 301912 310420
rect 301976 310406 302174 310434
rect 301976 306338 302004 310406
rect 302344 306354 302372 310420
rect 302528 310406 302634 310434
rect 301964 306332 302016 306338
rect 301964 306274 302016 306280
rect 302252 306326 302372 306354
rect 302424 306400 302476 306406
rect 302424 306342 302476 306348
rect 301872 303204 301924 303210
rect 301872 303146 301924 303152
rect 301332 296686 301544 296714
rect 301228 253564 301280 253570
rect 301228 253506 301280 253512
rect 301332 253502 301360 296686
rect 301320 253496 301372 253502
rect 301320 253438 301372 253444
rect 301134 250744 301190 250753
rect 301134 250679 301190 250688
rect 302252 245585 302280 306326
rect 302332 306264 302384 306270
rect 302332 306206 302384 306212
rect 302344 249121 302372 306206
rect 302436 254794 302464 306342
rect 302528 260137 302556 310406
rect 302608 306332 302660 306338
rect 302608 306274 302660 306280
rect 302620 267073 302648 306274
rect 302804 296714 302832 310420
rect 302896 310406 303094 310434
rect 302896 306406 302924 310406
rect 302884 306400 302936 306406
rect 302884 306342 302936 306348
rect 303264 306338 303292 310420
rect 303356 310406 303554 310434
rect 303252 306332 303304 306338
rect 303252 306274 303304 306280
rect 303356 306270 303384 310406
rect 303724 306456 303752 310420
rect 303632 306428 303752 306456
rect 303816 310406 304014 310434
rect 303632 306270 303660 306428
rect 303816 306354 303844 310406
rect 304184 306354 304212 310420
rect 303724 306326 303844 306354
rect 303908 306326 304212 306354
rect 304276 310406 304474 310434
rect 303344 306264 303396 306270
rect 303344 306206 303396 306212
rect 303620 306264 303672 306270
rect 303620 306206 303672 306212
rect 303620 306060 303672 306066
rect 303620 306002 303672 306008
rect 302712 296686 302832 296714
rect 302712 284889 302740 296686
rect 302698 284880 302754 284889
rect 302698 284815 302754 284824
rect 302606 267064 302662 267073
rect 302606 266999 302662 267008
rect 302514 260128 302570 260137
rect 302514 260063 302570 260072
rect 302424 254788 302476 254794
rect 302424 254730 302476 254736
rect 303632 254561 303660 306002
rect 303724 268666 303752 306326
rect 303804 306128 303856 306134
rect 303804 306070 303856 306076
rect 303816 269793 303844 306070
rect 303908 286385 303936 306326
rect 304080 306264 304132 306270
rect 304080 306206 304132 306212
rect 303988 306196 304040 306202
rect 303988 306138 304040 306144
rect 304000 287910 304028 306138
rect 304092 298761 304120 306206
rect 304276 306066 304304 310406
rect 304644 306134 304672 310420
rect 304736 310406 304934 310434
rect 304736 306202 304764 310406
rect 304724 306196 304776 306202
rect 304724 306138 304776 306144
rect 304632 306128 304684 306134
rect 304632 306070 304684 306076
rect 304264 306060 304316 306066
rect 304264 306002 304316 306008
rect 304078 298752 304134 298761
rect 304078 298687 304134 298696
rect 303988 287904 304040 287910
rect 303988 287846 304040 287852
rect 303894 286376 303950 286385
rect 303894 286311 303950 286320
rect 305012 270026 305040 310490
rect 305118 310406 305316 310434
rect 305092 306400 305144 306406
rect 305092 306342 305144 306348
rect 305288 306354 305316 310406
rect 305104 271386 305132 306342
rect 305184 306332 305236 306338
rect 305288 306326 305408 306354
rect 305184 306274 305236 306280
rect 305196 287774 305224 306274
rect 305276 302388 305328 302394
rect 305276 302330 305328 302336
rect 305288 287842 305316 302330
rect 305380 300490 305408 306326
rect 305564 302394 305592 310420
rect 305656 310406 305854 310434
rect 305552 302388 305604 302394
rect 305552 302330 305604 302336
rect 305656 301850 305684 310406
rect 306024 306406 306052 310420
rect 306116 310406 306314 310434
rect 306012 306400 306064 306406
rect 306012 306342 306064 306348
rect 306116 306338 306144 310406
rect 306104 306332 306156 306338
rect 306104 306274 306156 306280
rect 306380 306332 306432 306338
rect 306380 306274 306432 306280
rect 305644 301844 305696 301850
rect 305644 301786 305696 301792
rect 305368 300484 305420 300490
rect 305368 300426 305420 300432
rect 305276 287836 305328 287842
rect 305276 287778 305328 287784
rect 305184 287768 305236 287774
rect 305184 287710 305236 287716
rect 305092 271380 305144 271386
rect 305092 271322 305144 271328
rect 305000 270020 305052 270026
rect 305000 269962 305052 269968
rect 303802 269784 303858 269793
rect 303802 269719 303858 269728
rect 303712 268660 303764 268666
rect 303712 268602 303764 268608
rect 303618 254552 303674 254561
rect 303618 254487 303674 254496
rect 306392 250578 306420 306274
rect 306668 303346 306696 310542
rect 309416 310490 309468 310496
rect 309784 310548 309836 310554
rect 310638 310548 310848 310554
rect 310638 310542 310796 310548
rect 309784 310490 309836 310496
rect 310796 310490 310848 310496
rect 311164 310548 311216 310554
rect 312018 310548 312228 310554
rect 312018 310542 312176 310548
rect 311164 310490 311216 310496
rect 312176 310490 312228 310496
rect 312544 310548 312596 310554
rect 362986 310542 363184 310570
rect 312544 310490 312596 310496
rect 306656 303340 306708 303346
rect 306656 303282 306708 303288
rect 306760 303226 306788 310420
rect 306484 303198 306788 303226
rect 306484 271318 306512 303198
rect 306564 303068 306616 303074
rect 306564 303010 306616 303016
rect 306472 271312 306524 271318
rect 306472 271254 306524 271260
rect 306576 271250 306604 303010
rect 306944 302234 306972 310420
rect 307220 303278 307248 310420
rect 307208 303272 307260 303278
rect 307208 303214 307260 303220
rect 307404 303074 307432 310420
rect 307496 310406 307694 310434
rect 307496 306338 307524 310406
rect 307864 306490 307892 310420
rect 307864 306462 308076 306490
rect 307852 306400 307904 306406
rect 307852 306342 307904 306348
rect 307484 306332 307536 306338
rect 307484 306274 307536 306280
rect 307760 306332 307812 306338
rect 307760 306274 307812 306280
rect 307392 303068 307444 303074
rect 307392 303010 307444 303016
rect 306668 302206 306972 302234
rect 306668 289338 306696 302206
rect 306656 289332 306708 289338
rect 306656 289274 306708 289280
rect 306564 271244 306616 271250
rect 306564 271186 306616 271192
rect 306380 250572 306432 250578
rect 306380 250514 306432 250520
rect 307772 250510 307800 306274
rect 307864 272610 307892 306342
rect 308048 303210 308076 306462
rect 308036 303204 308088 303210
rect 308036 303146 308088 303152
rect 308140 303090 308168 310420
rect 308324 306338 308352 310420
rect 308312 306332 308364 306338
rect 308312 306274 308364 306280
rect 308600 304434 308628 310420
rect 308784 306406 308812 310420
rect 308876 310406 309074 310434
rect 309336 310406 309534 310434
rect 308772 306400 308824 306406
rect 308772 306342 308824 306348
rect 308588 304428 308640 304434
rect 308588 304370 308640 304376
rect 307956 303062 308168 303090
rect 307956 272678 307984 303062
rect 308876 302234 308904 310406
rect 309336 306456 309364 310406
rect 308048 302206 308904 302234
rect 309152 306428 309364 306456
rect 308048 289270 308076 302206
rect 308036 289264 308088 289270
rect 308036 289206 308088 289212
rect 307944 272672 307996 272678
rect 307944 272614 307996 272620
rect 307852 272604 307904 272610
rect 307852 272546 307904 272552
rect 309152 272542 309180 306428
rect 309704 306354 309732 310420
rect 309232 306332 309284 306338
rect 309232 306274 309284 306280
rect 309336 306326 309732 306354
rect 309244 274174 309272 306274
rect 309336 289202 309364 306326
rect 309796 304337 309824 310490
rect 309782 304328 309838 304337
rect 309782 304263 309838 304272
rect 309980 304201 310008 310420
rect 310164 306338 310192 310420
rect 310256 310406 310454 310434
rect 310716 310406 310914 310434
rect 310152 306332 310204 306338
rect 310152 306274 310204 306280
rect 309966 304192 310022 304201
rect 309966 304127 310022 304136
rect 310256 302234 310284 310406
rect 310716 306456 310744 310406
rect 310624 306428 310744 306456
rect 310520 306332 310572 306338
rect 310520 306274 310572 306280
rect 309428 302206 310284 302234
rect 309428 290698 309456 302206
rect 309416 290692 309468 290698
rect 309416 290634 309468 290640
rect 309324 289196 309376 289202
rect 309324 289138 309376 289144
rect 309232 274168 309284 274174
rect 309232 274110 309284 274116
rect 309140 272536 309192 272542
rect 309140 272478 309192 272484
rect 307760 250504 307812 250510
rect 307760 250446 307812 250452
rect 302330 249112 302386 249121
rect 302330 249047 302386 249056
rect 310532 246634 310560 306274
rect 310624 274106 310652 306428
rect 311084 306354 311112 310420
rect 310716 306326 311112 306354
rect 310716 290630 310744 306326
rect 311176 306105 311204 310490
rect 311162 306096 311218 306105
rect 311162 306031 311218 306040
rect 311360 305969 311388 310420
rect 311544 306338 311572 310420
rect 311636 310406 311834 310434
rect 312096 310406 312294 310434
rect 311532 306332 311584 306338
rect 311532 306274 311584 306280
rect 311346 305960 311402 305969
rect 311346 305895 311402 305904
rect 311636 302234 311664 310406
rect 312096 306490 312124 310406
rect 310808 302206 311664 302234
rect 311912 306462 312124 306490
rect 310704 290624 310756 290630
rect 310704 290566 310756 290572
rect 310808 290562 310836 302206
rect 310796 290556 310848 290562
rect 310796 290498 310848 290504
rect 310612 274100 310664 274106
rect 310612 274042 310664 274048
rect 311912 265878 311940 306462
rect 312464 306354 312492 310420
rect 311992 306332 312044 306338
rect 311992 306274 312044 306280
rect 312096 306326 312492 306354
rect 312004 274038 312032 306274
rect 312096 292058 312124 306326
rect 312556 305833 312584 310490
rect 312740 307057 312768 310420
rect 312726 307048 312782 307057
rect 312726 306983 312782 306992
rect 312924 306338 312952 310420
rect 313016 310406 313214 310434
rect 312912 306332 312964 306338
rect 312912 306274 312964 306280
rect 312542 305824 312598 305833
rect 312542 305759 312598 305768
rect 313016 302234 313044 310406
rect 313384 306320 313412 310420
rect 312188 302206 313044 302234
rect 313292 306292 313412 306320
rect 313476 310406 313674 310434
rect 312084 292052 312136 292058
rect 312084 291994 312136 292000
rect 312188 291990 312216 302206
rect 312176 291984 312228 291990
rect 312176 291926 312228 291932
rect 311992 274032 312044 274038
rect 311992 273974 312044 273980
rect 311900 265872 311952 265878
rect 311900 265814 311952 265820
rect 313292 254726 313320 306292
rect 313476 306252 313504 310406
rect 313844 306354 313872 310420
rect 313384 306224 313504 306252
rect 313568 306326 313872 306354
rect 313384 275466 313412 306224
rect 313464 306128 313516 306134
rect 313464 306070 313516 306076
rect 313372 275460 313424 275466
rect 313372 275402 313424 275408
rect 313476 275398 313504 306070
rect 313568 282402 313596 306326
rect 314120 304366 314148 310420
rect 314304 306134 314332 310420
rect 314396 310406 314594 310434
rect 314292 306128 314344 306134
rect 314292 306070 314344 306076
rect 314108 304360 314160 304366
rect 314108 304302 314160 304308
rect 314396 302234 314424 310406
rect 314856 307222 314884 310420
rect 314844 307216 314896 307222
rect 314844 307158 314896 307164
rect 315040 306490 315068 310420
rect 313660 302206 314424 302234
rect 314672 306462 315068 306490
rect 315132 310406 315330 310434
rect 313660 290494 313688 302206
rect 313648 290488 313700 290494
rect 313648 290430 313700 290436
rect 313556 282396 313608 282402
rect 313556 282338 313608 282344
rect 313464 275392 313516 275398
rect 313464 275334 313516 275340
rect 313280 254720 313332 254726
rect 313280 254662 313332 254668
rect 310520 246628 310572 246634
rect 310520 246570 310572 246576
rect 314672 246498 314700 306462
rect 315132 306354 315160 310406
rect 314752 306332 314804 306338
rect 314752 306274 314804 306280
rect 314856 306326 315160 306354
rect 314764 273970 314792 306274
rect 314856 291922 314884 306326
rect 315500 302841 315528 310420
rect 315592 310406 315790 310434
rect 315592 306338 315620 310406
rect 315580 306332 315632 306338
rect 315580 306274 315632 306280
rect 315486 302832 315542 302841
rect 315486 302767 315542 302776
rect 315960 302234 315988 310420
rect 316132 306400 316184 306406
rect 316236 306388 316264 310420
rect 316420 308990 316448 310420
rect 316512 310406 316710 310434
rect 316408 308984 316460 308990
rect 316408 308926 316460 308932
rect 316236 306360 316356 306388
rect 316132 306342 316184 306348
rect 316040 306332 316092 306338
rect 316040 306274 316092 306280
rect 314948 302206 315988 302234
rect 314948 293486 314976 302206
rect 314936 293480 314988 293486
rect 314936 293422 314988 293428
rect 314844 291916 314896 291922
rect 314844 291858 314896 291864
rect 314752 273964 314804 273970
rect 314752 273906 314804 273912
rect 316052 263022 316080 306274
rect 316144 276894 316172 306342
rect 316328 305697 316356 306360
rect 316314 305688 316370 305697
rect 316314 305623 316370 305632
rect 316512 305538 316540 310406
rect 316880 306338 316908 310420
rect 316972 310406 317170 310434
rect 316972 306406 317000 310406
rect 316960 306400 317012 306406
rect 316960 306342 317012 306348
rect 316868 306332 316920 306338
rect 316868 306274 316920 306280
rect 316236 305510 316540 305538
rect 316236 283830 316264 305510
rect 317340 302234 317368 310420
rect 317524 310406 317630 310434
rect 317420 304564 317472 304570
rect 317420 304506 317472 304512
rect 316328 302206 317368 302234
rect 316328 291854 316356 302206
rect 316316 291848 316368 291854
rect 316316 291790 316368 291796
rect 316224 283824 316276 283830
rect 316224 283766 316276 283772
rect 316132 276888 316184 276894
rect 316132 276830 316184 276836
rect 316040 263016 316092 263022
rect 316040 262958 316092 262964
rect 314660 246492 314712 246498
rect 314660 246434 314712 246440
rect 317432 246430 317460 304506
rect 317524 249286 317552 310406
rect 317800 307018 317828 310420
rect 317892 310406 318090 310434
rect 317788 307012 317840 307018
rect 317788 306954 317840 306960
rect 317788 306808 317840 306814
rect 317788 306750 317840 306756
rect 317696 306332 317748 306338
rect 317696 306274 317748 306280
rect 317604 304224 317656 304230
rect 317604 304166 317656 304172
rect 317616 250617 317644 304166
rect 317708 264382 317736 306274
rect 317800 276826 317828 306750
rect 317892 304230 317920 310406
rect 318260 306338 318288 310420
rect 318352 310406 318550 310434
rect 318248 306332 318300 306338
rect 318248 306274 318300 306280
rect 318352 304570 318380 310406
rect 318340 304564 318392 304570
rect 318340 304506 318392 304512
rect 317880 304224 317932 304230
rect 317880 304166 317932 304172
rect 318720 296714 318748 310420
rect 318904 310406 319010 310434
rect 318800 306332 318852 306338
rect 318800 306274 318852 306280
rect 317892 296686 318748 296714
rect 317892 293418 317920 296686
rect 317880 293412 317932 293418
rect 317880 293354 317932 293360
rect 317788 276820 317840 276826
rect 317788 276762 317840 276768
rect 317696 264376 317748 264382
rect 317696 264318 317748 264324
rect 318812 252074 318840 306274
rect 318904 254658 318932 310406
rect 319180 306320 319208 310420
rect 318996 306292 319208 306320
rect 319272 310406 319470 310434
rect 318996 271182 319024 306292
rect 319168 306196 319220 306202
rect 319168 306138 319220 306144
rect 319076 306128 319128 306134
rect 319076 306070 319128 306076
rect 319088 275330 319116 306070
rect 319180 286550 319208 306138
rect 319272 287706 319300 310406
rect 319640 306202 319668 310420
rect 319732 310406 319930 310434
rect 319628 306196 319680 306202
rect 319628 306138 319680 306144
rect 319732 306134 319760 310406
rect 320100 306338 320128 310420
rect 320088 306332 320140 306338
rect 320088 306274 320140 306280
rect 320180 306332 320232 306338
rect 320180 306274 320232 306280
rect 319720 306128 319772 306134
rect 319720 306070 319772 306076
rect 319260 287700 319312 287706
rect 319260 287642 319312 287648
rect 319168 286544 319220 286550
rect 319168 286486 319220 286492
rect 319076 275324 319128 275330
rect 319076 275266 319128 275272
rect 318984 271176 319036 271182
rect 318984 271118 319036 271124
rect 318892 254652 318944 254658
rect 318892 254594 318944 254600
rect 318800 252068 318852 252074
rect 318800 252010 318852 252016
rect 320192 251938 320220 306274
rect 320272 303748 320324 303754
rect 320272 303690 320324 303696
rect 320284 252006 320312 303690
rect 320376 269958 320404 310420
rect 320560 306320 320588 310420
rect 320468 306292 320588 306320
rect 320652 310406 320850 310434
rect 320468 276758 320496 306292
rect 320548 306196 320600 306202
rect 320548 306138 320600 306144
rect 320560 278254 320588 306138
rect 320652 303754 320680 310406
rect 320640 303748 320692 303754
rect 320640 303690 320692 303696
rect 321020 298994 321048 310420
rect 321112 310406 321310 310434
rect 321112 306202 321140 310406
rect 321480 306338 321508 310420
rect 321652 306400 321704 306406
rect 321652 306342 321704 306348
rect 321756 306354 321784 310420
rect 321940 307154 321968 310420
rect 322032 310406 322230 310434
rect 321928 307148 321980 307154
rect 321928 307090 321980 307096
rect 321468 306332 321520 306338
rect 321468 306274 321520 306280
rect 321560 306332 321612 306338
rect 321560 306274 321612 306280
rect 321100 306196 321152 306202
rect 321100 306138 321152 306144
rect 321008 298988 321060 298994
rect 321008 298930 321060 298936
rect 320548 278248 320600 278254
rect 320548 278190 320600 278196
rect 320456 276752 320508 276758
rect 320456 276694 320508 276700
rect 320364 269952 320416 269958
rect 320364 269894 320416 269900
rect 321572 256222 321600 306274
rect 321664 278186 321692 306342
rect 321756 306326 321968 306354
rect 321744 306264 321796 306270
rect 321744 306206 321796 306212
rect 321756 293350 321784 306206
rect 321836 306196 321888 306202
rect 321836 306138 321888 306144
rect 321848 294846 321876 306138
rect 321940 300422 321968 306326
rect 322032 306270 322060 310406
rect 322400 306338 322428 310420
rect 322492 310406 322690 310434
rect 322492 306406 322520 310406
rect 322480 306400 322532 306406
rect 322480 306342 322532 306348
rect 322388 306332 322440 306338
rect 322388 306274 322440 306280
rect 322020 306264 322072 306270
rect 322020 306206 322072 306212
rect 322860 306202 322888 310420
rect 323136 309134 323164 310420
rect 323136 309106 323256 309134
rect 323032 306332 323084 306338
rect 323032 306274 323084 306280
rect 322848 306196 322900 306202
rect 322848 306138 322900 306144
rect 322940 304224 322992 304230
rect 322940 304166 322992 304172
rect 321928 300416 321980 300422
rect 321928 300358 321980 300364
rect 321836 294840 321888 294846
rect 321836 294782 321888 294788
rect 321744 293344 321796 293350
rect 321744 293286 321796 293292
rect 321652 278180 321704 278186
rect 321652 278122 321704 278128
rect 321560 256216 321612 256222
rect 321560 256158 321612 256164
rect 320272 252000 320324 252006
rect 320272 251942 320324 251948
rect 320180 251932 320232 251938
rect 320180 251874 320232 251880
rect 317602 250608 317658 250617
rect 317602 250543 317658 250552
rect 317512 249280 317564 249286
rect 317512 249222 317564 249228
rect 322952 248033 322980 304166
rect 323044 251870 323072 306274
rect 323124 306264 323176 306270
rect 323124 306206 323176 306212
rect 323032 251864 323084 251870
rect 323032 251806 323084 251812
rect 322938 248024 322994 248033
rect 322938 247959 322994 247968
rect 323136 247897 323164 306206
rect 323228 256154 323256 309106
rect 323320 304230 323348 310420
rect 323412 310406 323610 310434
rect 323412 306338 323440 310406
rect 323780 309126 323808 310420
rect 323872 310406 324070 310434
rect 323768 309120 323820 309126
rect 323768 309062 323820 309068
rect 323400 306332 323452 306338
rect 323400 306274 323452 306280
rect 323872 306270 323900 310406
rect 323860 306264 323912 306270
rect 323860 306206 323912 306212
rect 323308 304224 323360 304230
rect 323308 304166 323360 304172
rect 324240 296714 324268 310420
rect 324516 309058 324544 310420
rect 324504 309052 324556 309058
rect 324504 308994 324556 309000
rect 324320 306400 324372 306406
rect 324320 306342 324372 306348
rect 323320 296686 324268 296714
rect 323320 289134 323348 296686
rect 323308 289128 323360 289134
rect 323308 289070 323360 289076
rect 323216 256148 323268 256154
rect 323216 256090 323268 256096
rect 323122 247888 323178 247897
rect 323122 247823 323178 247832
rect 324332 247625 324360 306342
rect 324412 306332 324464 306338
rect 324412 306274 324464 306280
rect 324424 256086 324452 306274
rect 324700 304314 324728 310420
rect 324516 304286 324728 304314
rect 324792 310406 324990 310434
rect 324412 256080 324464 256086
rect 324412 256022 324464 256028
rect 324516 247761 324544 304286
rect 324596 304224 324648 304230
rect 324596 304166 324648 304172
rect 324608 293282 324636 304166
rect 324792 296714 324820 310406
rect 325160 306338 325188 310420
rect 325252 310406 325450 310434
rect 325252 306406 325280 310406
rect 325240 306400 325292 306406
rect 325240 306342 325292 306348
rect 325148 306332 325200 306338
rect 325148 306274 325200 306280
rect 325620 304230 325648 310420
rect 325712 310406 325910 310434
rect 325608 304224 325660 304230
rect 325608 304166 325660 304172
rect 324700 296686 324820 296714
rect 324700 294778 324728 296686
rect 324688 294772 324740 294778
rect 324688 294714 324740 294720
rect 324596 293276 324648 293282
rect 324596 293218 324648 293224
rect 325712 256018 325740 310406
rect 326080 307018 326108 310420
rect 326172 310406 326370 310434
rect 326068 307012 326120 307018
rect 326068 306954 326120 306960
rect 326172 306354 326200 310406
rect 326344 308984 326396 308990
rect 326344 308926 326396 308932
rect 326356 308106 326384 308926
rect 326344 308100 326396 308106
rect 326344 308042 326396 308048
rect 325792 306332 325844 306338
rect 325792 306274 325844 306280
rect 325896 306326 326200 306354
rect 325804 260234 325832 306274
rect 325896 278118 325924 306326
rect 325976 306264 326028 306270
rect 325976 306206 326028 306212
rect 325988 279682 326016 306206
rect 326540 296714 326568 310420
rect 326632 310406 326830 310434
rect 326632 306338 326660 310406
rect 326620 306332 326672 306338
rect 326620 306274 326672 306280
rect 327000 306270 327028 310420
rect 327080 306468 327132 306474
rect 327080 306410 327132 306416
rect 326988 306264 327040 306270
rect 326988 306206 327040 306212
rect 326080 296686 326568 296714
rect 326080 294710 326108 296686
rect 326068 294704 326120 294710
rect 326068 294646 326120 294652
rect 325976 279676 326028 279682
rect 325976 279618 326028 279624
rect 325884 278112 325936 278118
rect 325884 278054 325936 278060
rect 327092 261730 327120 306410
rect 327276 306354 327304 310420
rect 327460 306474 327488 310420
rect 327552 310406 327750 310434
rect 327448 306468 327500 306474
rect 327448 306410 327500 306416
rect 327172 306332 327224 306338
rect 327276 306326 327488 306354
rect 327172 306274 327224 306280
rect 327080 261724 327132 261730
rect 327080 261666 327132 261672
rect 327184 261662 327212 306274
rect 327264 306264 327316 306270
rect 327264 306206 327316 306212
rect 327276 278050 327304 306206
rect 327356 306196 327408 306202
rect 327356 306138 327408 306144
rect 327368 279614 327396 306138
rect 327460 285190 327488 306326
rect 327552 306270 327580 310406
rect 327540 306264 327592 306270
rect 327540 306206 327592 306212
rect 327920 296714 327948 310420
rect 328012 310406 328210 310434
rect 328012 306338 328040 310406
rect 328000 306332 328052 306338
rect 328000 306274 328052 306280
rect 328380 306202 328408 310420
rect 328656 306610 328684 310420
rect 328644 306604 328696 306610
rect 328644 306546 328696 306552
rect 328840 306490 328868 310420
rect 328564 306462 328868 306490
rect 328932 310406 329130 310434
rect 328460 306400 328512 306406
rect 328460 306342 328512 306348
rect 328368 306196 328420 306202
rect 328368 306138 328420 306144
rect 327552 296686 327948 296714
rect 327552 296206 327580 296686
rect 327540 296200 327592 296206
rect 327540 296142 327592 296148
rect 327448 285184 327500 285190
rect 327448 285126 327500 285132
rect 327356 279608 327408 279614
rect 327356 279550 327408 279556
rect 327264 278044 327316 278050
rect 327264 277986 327316 277992
rect 327172 261656 327224 261662
rect 327172 261598 327224 261604
rect 325792 260228 325844 260234
rect 325792 260170 325844 260176
rect 325700 256012 325752 256018
rect 325700 255954 325752 255960
rect 324502 247752 324558 247761
rect 324502 247687 324558 247696
rect 324318 247616 324374 247625
rect 324318 247551 324374 247560
rect 317420 246424 317472 246430
rect 317420 246366 317472 246372
rect 328472 246362 328500 306342
rect 328564 261594 328592 306462
rect 328932 306354 328960 310406
rect 329012 306604 329064 306610
rect 329012 306546 329064 306552
rect 328644 306332 328696 306338
rect 328644 306274 328696 306280
rect 328748 306326 328960 306354
rect 328656 262954 328684 306274
rect 328748 279546 328776 306326
rect 328828 306264 328880 306270
rect 328828 306206 328880 306212
rect 328840 281042 328868 306206
rect 329024 296714 329052 306546
rect 329300 306406 329328 310420
rect 329392 310406 329590 310434
rect 329288 306400 329340 306406
rect 329288 306342 329340 306348
rect 329392 306338 329420 310406
rect 329380 306332 329432 306338
rect 329380 306274 329432 306280
rect 329760 306270 329788 310420
rect 329932 306400 329984 306406
rect 329932 306342 329984 306348
rect 329840 306332 329892 306338
rect 329840 306274 329892 306280
rect 329748 306264 329800 306270
rect 329748 306206 329800 306212
rect 328932 296686 329052 296714
rect 328932 296138 328960 296686
rect 328920 296132 328972 296138
rect 328920 296074 328972 296080
rect 328828 281036 328880 281042
rect 328828 280978 328880 280984
rect 328736 279540 328788 279546
rect 328736 279482 328788 279488
rect 328644 262948 328696 262954
rect 328644 262890 328696 262896
rect 328552 261588 328604 261594
rect 328552 261530 328604 261536
rect 328460 246356 328512 246362
rect 328460 246298 328512 246304
rect 302238 245576 302294 245585
rect 302238 245511 302294 245520
rect 301044 245472 301096 245478
rect 301044 245414 301096 245420
rect 300858 245304 300914 245313
rect 300858 245239 300914 245248
rect 329852 245138 329880 306274
rect 329944 262857 329972 306342
rect 330036 306218 330064 310420
rect 330220 306406 330248 310420
rect 330312 310406 330510 310434
rect 330208 306400 330260 306406
rect 330208 306342 330260 306348
rect 330312 306338 330340 310406
rect 330300 306332 330352 306338
rect 330300 306274 330352 306280
rect 330036 306190 330156 306218
rect 330024 306128 330076 306134
rect 330024 306070 330076 306076
rect 330036 263090 330064 306070
rect 330128 296070 330156 306190
rect 330680 297634 330708 310420
rect 330772 310406 330970 310434
rect 330772 306134 330800 310406
rect 331128 308984 331180 308990
rect 331128 308926 331180 308932
rect 331140 308258 331168 308926
rect 331232 308394 331260 310420
rect 331416 308530 331444 310420
rect 331508 310406 331706 310434
rect 331508 308990 331536 310406
rect 331496 308984 331548 308990
rect 331496 308926 331548 308932
rect 331416 308502 331720 308530
rect 331232 308366 331444 308394
rect 331140 308230 331260 308258
rect 330760 306128 330812 306134
rect 330760 306070 330812 306076
rect 330668 297628 330720 297634
rect 330668 297570 330720 297576
rect 330116 296064 330168 296070
rect 330116 296006 330168 296012
rect 331232 264314 331260 308230
rect 331312 306264 331364 306270
rect 331312 306206 331364 306212
rect 331220 264308 331272 264314
rect 331220 264250 331272 264256
rect 331324 264246 331352 306206
rect 331416 280974 331444 308366
rect 331588 306400 331640 306406
rect 331588 306342 331640 306348
rect 331496 306332 331548 306338
rect 331496 306274 331548 306280
rect 331404 280968 331456 280974
rect 331404 280910 331456 280916
rect 331508 280906 331536 306274
rect 331600 297498 331628 306342
rect 331692 297566 331720 308502
rect 331772 308100 331824 308106
rect 331772 308042 331824 308048
rect 331784 302234 331812 308042
rect 331876 306338 331904 310420
rect 331968 310406 332166 310434
rect 331968 306406 331996 310406
rect 331956 306400 332008 306406
rect 331956 306342 332008 306348
rect 331864 306332 331916 306338
rect 331864 306274 331916 306280
rect 332336 306270 332364 310420
rect 332612 306270 332640 310420
rect 332692 306604 332744 306610
rect 332692 306546 332744 306552
rect 332324 306264 332376 306270
rect 332324 306206 332376 306212
rect 332600 306264 332652 306270
rect 332600 306206 332652 306212
rect 332600 306128 332652 306134
rect 332600 306070 332652 306076
rect 331784 302206 331904 302234
rect 331680 297560 331732 297566
rect 331680 297502 331732 297508
rect 331588 297492 331640 297498
rect 331588 297434 331640 297440
rect 331496 280900 331548 280906
rect 331496 280842 331548 280848
rect 331312 264240 331364 264246
rect 331312 264182 331364 264188
rect 330024 263084 330076 263090
rect 330024 263026 330076 263032
rect 329930 262848 329986 262857
rect 329930 262783 329986 262792
rect 331876 246566 331904 302206
rect 332612 253434 332640 306070
rect 332704 264450 332732 306546
rect 332796 306252 332824 310420
rect 332888 310406 333086 310434
rect 332888 306610 332916 310406
rect 332876 306604 332928 306610
rect 332876 306546 332928 306552
rect 332968 306264 333020 306270
rect 332796 306224 332916 306252
rect 332784 306060 332836 306066
rect 332784 306002 332836 306008
rect 332796 265810 332824 306002
rect 332888 268462 332916 306224
rect 332968 306206 333020 306212
rect 332980 276690 333008 306206
rect 333256 296714 333284 310420
rect 333348 310406 333546 310434
rect 333348 306134 333376 310406
rect 333336 306128 333388 306134
rect 333336 306070 333388 306076
rect 333716 306066 333744 310420
rect 333992 306202 334020 310420
rect 334176 306320 334204 310420
rect 334084 306292 334204 306320
rect 334268 310406 334466 310434
rect 333980 306196 334032 306202
rect 333980 306138 334032 306144
rect 333704 306060 333756 306066
rect 333704 306002 333756 306008
rect 333980 306060 334032 306066
rect 333980 306002 334032 306008
rect 333072 296686 333284 296714
rect 333072 282334 333100 296686
rect 333060 282328 333112 282334
rect 333060 282270 333112 282276
rect 332968 276684 333020 276690
rect 332968 276626 333020 276632
rect 332876 268456 332928 268462
rect 332876 268398 332928 268404
rect 332784 265804 332836 265810
rect 332784 265746 332836 265752
rect 332692 264444 332744 264450
rect 332692 264386 332744 264392
rect 332600 253428 332652 253434
rect 332600 253370 332652 253376
rect 333992 253298 334020 306002
rect 334084 253366 334112 306292
rect 334164 306128 334216 306134
rect 334164 306070 334216 306076
rect 334176 265674 334204 306070
rect 334268 265742 334296 310406
rect 334636 306320 334664 310420
rect 334360 306292 334664 306320
rect 334728 310406 334926 310434
rect 334360 267102 334388 306292
rect 334440 306196 334492 306202
rect 334440 306138 334492 306144
rect 334452 282266 334480 306138
rect 334728 306066 334756 310406
rect 335096 306134 335124 310420
rect 335372 306320 335400 310420
rect 335570 310406 335768 310434
rect 335636 306332 335688 306338
rect 335372 306292 335584 306320
rect 335360 306196 335412 306202
rect 335360 306138 335412 306144
rect 335084 306128 335136 306134
rect 335084 306070 335136 306076
rect 334716 306060 334768 306066
rect 334716 306002 334768 306008
rect 334440 282260 334492 282266
rect 334440 282202 334492 282208
rect 334348 267096 334400 267102
rect 334348 267038 334400 267044
rect 334256 265736 334308 265742
rect 334256 265678 334308 265684
rect 334164 265668 334216 265674
rect 334164 265610 334216 265616
rect 335372 260166 335400 306138
rect 335452 304700 335504 304706
rect 335452 304642 335504 304648
rect 335464 267238 335492 304642
rect 335556 282198 335584 306292
rect 335636 306274 335688 306280
rect 335648 283762 335676 306274
rect 335740 294642 335768 310406
rect 335832 306202 335860 310420
rect 336016 306338 336044 310420
rect 336108 310406 336306 310434
rect 336004 306332 336056 306338
rect 336004 306274 336056 306280
rect 335820 306196 335872 306202
rect 335820 306138 335872 306144
rect 336108 298926 336136 310406
rect 336476 304706 336504 310420
rect 336752 306320 336780 310420
rect 336832 307012 336884 307018
rect 336832 306954 336884 306960
rect 336844 306388 336872 306954
rect 336936 306490 336964 310420
rect 337028 310406 337226 310434
rect 337028 307018 337056 310406
rect 337016 307012 337068 307018
rect 337016 306954 337068 306960
rect 336936 306462 337240 306490
rect 336844 306360 336964 306388
rect 336752 306292 336872 306320
rect 336740 306128 336792 306134
rect 336740 306070 336792 306076
rect 336464 304700 336516 304706
rect 336464 304642 336516 304648
rect 336096 298920 336148 298926
rect 336096 298862 336148 298868
rect 335728 294636 335780 294642
rect 335728 294578 335780 294584
rect 335636 283756 335688 283762
rect 335636 283698 335688 283704
rect 335544 282192 335596 282198
rect 335544 282134 335596 282140
rect 335452 267232 335504 267238
rect 335452 267174 335504 267180
rect 335360 260160 335412 260166
rect 335360 260102 335412 260108
rect 334072 253360 334124 253366
rect 334072 253302 334124 253308
rect 333980 253292 334032 253298
rect 333980 253234 334032 253240
rect 336752 249082 336780 306070
rect 336844 249150 336872 306292
rect 336936 267170 336964 306360
rect 337108 306332 337160 306338
rect 337108 306274 337160 306280
rect 337016 306196 337068 306202
rect 337016 306138 337068 306144
rect 336924 267164 336976 267170
rect 336924 267106 336976 267112
rect 337028 267034 337056 306138
rect 337120 298790 337148 306274
rect 337212 298858 337240 306462
rect 337396 306134 337424 310420
rect 337488 310406 337686 310434
rect 337488 306338 337516 310406
rect 337476 306332 337528 306338
rect 337476 306274 337528 306280
rect 337856 306202 337884 310420
rect 337844 306196 337896 306202
rect 337844 306138 337896 306144
rect 337384 306128 337436 306134
rect 337384 306070 337436 306076
rect 337200 298852 337252 298858
rect 337200 298794 337252 298800
rect 337108 298784 337160 298790
rect 337108 298726 337160 298732
rect 337016 267028 337068 267034
rect 337016 266970 337068 266976
rect 338132 249218 338160 310420
rect 338316 306490 338344 310420
rect 338224 306462 338344 306490
rect 338408 310406 338606 310434
rect 338224 306202 338252 306462
rect 338408 306320 338436 310406
rect 338776 306320 338804 310420
rect 338316 306292 338436 306320
rect 338500 306292 338804 306320
rect 338868 310406 339066 310434
rect 338212 306196 338264 306202
rect 338212 306138 338264 306144
rect 338212 306060 338264 306066
rect 338212 306002 338264 306008
rect 338224 250481 338252 306002
rect 338316 261526 338344 306292
rect 338396 306128 338448 306134
rect 338396 306070 338448 306076
rect 338408 268394 338436 306070
rect 338500 279478 338528 306292
rect 338580 306196 338632 306202
rect 338580 306138 338632 306144
rect 338592 300286 338620 306138
rect 338868 306066 338896 310406
rect 339236 306134 339264 310420
rect 339512 306320 339540 310420
rect 339710 310406 339816 310434
rect 339512 306292 339724 306320
rect 339500 306196 339552 306202
rect 339500 306138 339552 306144
rect 339224 306128 339276 306134
rect 339224 306070 339276 306076
rect 338856 306060 338908 306066
rect 338856 306002 338908 306008
rect 338580 300280 338632 300286
rect 338580 300222 338632 300228
rect 338488 279472 338540 279478
rect 338488 279414 338540 279420
rect 339512 268598 339540 306138
rect 339592 306128 339644 306134
rect 339592 306070 339644 306076
rect 339500 268592 339552 268598
rect 339500 268534 339552 268540
rect 339604 268530 339632 306070
rect 339696 283694 339724 306292
rect 339788 300218 339816 310406
rect 339972 306202 340000 310420
rect 339960 306196 340012 306202
rect 339960 306138 340012 306144
rect 339776 300212 339828 300218
rect 339776 300154 339828 300160
rect 340156 299474 340184 310420
rect 340248 310406 340446 310434
rect 340248 300150 340276 310406
rect 340616 306134 340644 310420
rect 340892 306354 340920 310420
rect 341090 310406 341288 310434
rect 340892 306326 341104 306354
rect 340972 306264 341024 306270
rect 340972 306206 341024 306212
rect 340880 306196 340932 306202
rect 340880 306138 340932 306144
rect 340604 306128 340656 306134
rect 340604 306070 340656 306076
rect 340236 300144 340288 300150
rect 340236 300086 340288 300092
rect 339788 299446 340184 299474
rect 339684 283688 339736 283694
rect 339684 283630 339736 283636
rect 339788 283626 339816 299446
rect 339776 283620 339828 283626
rect 339776 283562 339828 283568
rect 339592 268524 339644 268530
rect 339592 268466 339644 268472
rect 338396 268388 338448 268394
rect 338396 268330 338448 268336
rect 338304 261520 338356 261526
rect 338304 261462 338356 261468
rect 338210 250472 338266 250481
rect 338210 250407 338266 250416
rect 338120 249212 338172 249218
rect 338120 249154 338172 249160
rect 336832 249144 336884 249150
rect 336832 249086 336884 249092
rect 336740 249076 336792 249082
rect 336740 249018 336792 249024
rect 331864 246560 331916 246566
rect 331864 246502 331916 246508
rect 329840 245132 329892 245138
rect 329840 245074 329892 245080
rect 340892 245002 340920 306138
rect 340984 245070 341012 306206
rect 341076 280838 341104 306326
rect 341156 306332 341208 306338
rect 341156 306274 341208 306280
rect 341168 285122 341196 306274
rect 341260 296002 341288 310406
rect 341352 306270 341380 310420
rect 341536 306338 341564 310420
rect 341628 310406 341826 310434
rect 341524 306332 341576 306338
rect 341524 306274 341576 306280
rect 341340 306264 341392 306270
rect 341340 306206 341392 306212
rect 341628 301646 341656 310406
rect 341996 306202 342024 310420
rect 342272 306354 342300 310420
rect 342470 310406 342668 310434
rect 342640 306474 342668 310406
rect 342732 306542 342760 310420
rect 342720 306536 342772 306542
rect 342720 306478 342772 306484
rect 342628 306468 342680 306474
rect 342628 306410 342680 306416
rect 342916 306354 342944 310420
rect 342272 306326 342484 306354
rect 342260 306264 342312 306270
rect 342260 306206 342312 306212
rect 341984 306196 342036 306202
rect 341984 306138 342036 306144
rect 341616 301640 341668 301646
rect 341616 301582 341668 301588
rect 341248 295996 341300 296002
rect 341248 295938 341300 295944
rect 341156 285116 341208 285122
rect 341156 285058 341208 285064
rect 341064 280832 341116 280838
rect 341064 280774 341116 280780
rect 340972 245064 341024 245070
rect 340972 245006 341024 245012
rect 340880 244996 340932 245002
rect 340880 244938 340932 244944
rect 342272 244934 342300 306206
rect 342352 306060 342404 306066
rect 342352 306002 342404 306008
rect 342364 269890 342392 306002
rect 342456 285054 342484 306326
rect 342548 306326 342944 306354
rect 343008 310406 343206 310434
rect 342444 285048 342496 285054
rect 342444 284990 342496 284996
rect 342548 284986 342576 306326
rect 343008 306218 343036 310406
rect 342640 306190 343036 306218
rect 342640 297430 342668 306190
rect 342812 306128 342864 306134
rect 342812 306070 342864 306076
rect 342824 301578 342852 306070
rect 343376 306066 343404 310420
rect 343652 306474 343680 310420
rect 343640 306468 343692 306474
rect 343640 306410 343692 306416
rect 343836 306354 343864 310420
rect 343652 306326 343864 306354
rect 343928 310406 344126 310434
rect 343364 306060 343416 306066
rect 343364 306002 343416 306008
rect 342812 301572 342864 301578
rect 342812 301514 342864 301520
rect 342628 297424 342680 297430
rect 342628 297366 342680 297372
rect 342536 284980 342588 284986
rect 342536 284922 342588 284928
rect 342352 269884 342404 269890
rect 342352 269826 342404 269832
rect 343652 253230 343680 306326
rect 343732 306264 343784 306270
rect 343928 306218 343956 310406
rect 344008 306468 344060 306474
rect 344008 306410 344060 306416
rect 343732 306206 343784 306212
rect 343744 262886 343772 306206
rect 343836 306190 343956 306218
rect 343836 269822 343864 306190
rect 344020 306082 344048 306410
rect 343928 306054 344048 306082
rect 343928 286346 343956 306054
rect 344296 302234 344324 310420
rect 344020 302206 344324 302234
rect 344388 310406 344586 310434
rect 344020 286482 344048 302206
rect 344388 301510 344416 310406
rect 344756 306270 344784 310420
rect 345032 306354 345060 310420
rect 345230 310406 345428 310434
rect 345032 306326 345244 306354
rect 344744 306264 344796 306270
rect 344744 306206 344796 306212
rect 345020 306264 345072 306270
rect 345020 306206 345072 306212
rect 345032 301782 345060 306206
rect 345020 301776 345072 301782
rect 345020 301718 345072 301724
rect 344376 301504 344428 301510
rect 344376 301446 344428 301452
rect 344008 286476 344060 286482
rect 344008 286418 344060 286424
rect 345216 286414 345244 306326
rect 345204 286408 345256 286414
rect 345204 286350 345256 286356
rect 343916 286340 343968 286346
rect 343916 286282 343968 286288
rect 343824 269816 343876 269822
rect 343824 269758 343876 269764
rect 343732 262880 343784 262886
rect 343732 262822 343784 262828
rect 345400 254590 345428 310406
rect 345492 306270 345520 310420
rect 345480 306264 345532 306270
rect 345480 306206 345532 306212
rect 345676 305658 345704 310420
rect 345768 310406 345966 310434
rect 345664 305652 345716 305658
rect 345664 305594 345716 305600
rect 345768 296714 345796 310406
rect 346136 309097 346164 310420
rect 346122 309088 346178 309097
rect 346122 309023 346178 309032
rect 346412 308961 346440 310420
rect 346398 308952 346454 308961
rect 346398 308887 346454 308896
rect 346596 305658 346624 310420
rect 346584 305652 346636 305658
rect 346584 305594 346636 305600
rect 346872 303142 346900 310420
rect 347056 308825 347084 310420
rect 347042 308816 347098 308825
rect 347042 308751 347098 308760
rect 347332 308689 347360 310420
rect 347318 308680 347374 308689
rect 347318 308615 347374 308624
rect 347608 303414 347636 310420
rect 347596 303408 347648 303414
rect 347596 303350 347648 303356
rect 346860 303136 346912 303142
rect 346860 303078 346912 303084
rect 347792 303006 347820 310420
rect 347780 303000 347832 303006
rect 347780 302942 347832 302948
rect 348068 302938 348096 310420
rect 348252 305590 348280 310420
rect 348240 305584 348292 305590
rect 348240 305526 348292 305532
rect 348528 303142 348556 310420
rect 348516 303136 348568 303142
rect 348516 303078 348568 303084
rect 348712 302938 348740 310420
rect 348804 310406 349002 310434
rect 348056 302932 348108 302938
rect 348056 302874 348108 302880
rect 348700 302932 348752 302938
rect 348700 302874 348752 302880
rect 348804 296714 348832 310406
rect 349172 306241 349200 310420
rect 349158 306232 349214 306241
rect 349158 306167 349214 306176
rect 349448 302870 349476 310420
rect 349632 303006 349660 310420
rect 349724 310406 349922 310434
rect 349620 303000 349672 303006
rect 349620 302942 349672 302948
rect 349436 302864 349488 302870
rect 349436 302806 349488 302812
rect 349724 302234 349752 310406
rect 350092 305794 350120 310420
rect 350080 305788 350132 305794
rect 350080 305730 350132 305736
rect 350368 302802 350396 310420
rect 350356 302796 350408 302802
rect 350356 302738 350408 302744
rect 345492 296686 345796 296714
rect 348252 296686 348832 296714
rect 349172 302206 349752 302234
rect 345492 257378 345520 296686
rect 348252 294914 348280 296686
rect 349172 296274 349200 302206
rect 350552 300354 350580 310420
rect 350828 305318 350856 310420
rect 351012 308106 351040 310420
rect 351104 310406 351302 310434
rect 351000 308100 351052 308106
rect 351000 308042 351052 308048
rect 350816 305312 350868 305318
rect 350816 305254 350868 305260
rect 351104 302234 351132 310406
rect 351472 305454 351500 310420
rect 351460 305448 351512 305454
rect 351460 305390 351512 305396
rect 351748 303482 351776 310420
rect 351736 303476 351788 303482
rect 351736 303418 351788 303424
rect 351932 302666 351960 310420
rect 352208 305726 352236 310420
rect 352196 305720 352248 305726
rect 352196 305662 352248 305668
rect 352392 303550 352420 310420
rect 352668 304298 352696 310420
rect 352852 305930 352880 310420
rect 352840 305924 352892 305930
rect 352840 305866 352892 305872
rect 352656 304292 352708 304298
rect 352656 304234 352708 304240
rect 352380 303544 352432 303550
rect 352380 303486 352432 303492
rect 353128 303074 353156 310420
rect 353312 305386 353340 310420
rect 353300 305380 353352 305386
rect 353300 305322 353352 305328
rect 353588 303618 353616 310420
rect 353772 308281 353800 310420
rect 353758 308272 353814 308281
rect 353758 308207 353814 308216
rect 354048 305998 354076 310420
rect 354232 308990 354260 310420
rect 354220 308984 354272 308990
rect 354220 308926 354272 308932
rect 354036 305992 354088 305998
rect 354036 305934 354088 305940
rect 354508 305862 354536 310420
rect 354692 307970 354720 310420
rect 354680 307964 354732 307970
rect 354680 307906 354732 307912
rect 354968 306202 354996 310420
rect 355152 308242 355180 310420
rect 355324 308712 355376 308718
rect 355324 308654 355376 308660
rect 355428 308666 355456 310420
rect 355140 308236 355192 308242
rect 355140 308178 355192 308184
rect 354956 306196 355008 306202
rect 354956 306138 355008 306144
rect 354496 305856 354548 305862
rect 354496 305798 354548 305804
rect 353576 303612 353628 303618
rect 353576 303554 353628 303560
rect 353116 303068 353168 303074
rect 353116 303010 353168 303016
rect 351920 302660 351972 302666
rect 351920 302602 351972 302608
rect 350644 302206 351132 302234
rect 350644 301714 350672 302206
rect 350632 301708 350684 301714
rect 350632 301650 350684 301656
rect 350540 300348 350592 300354
rect 350540 300290 350592 300296
rect 349160 296268 349212 296274
rect 349160 296210 349212 296216
rect 348240 294908 348292 294914
rect 348240 294850 348292 294856
rect 345480 257372 345532 257378
rect 345480 257314 345532 257320
rect 345388 254584 345440 254590
rect 345388 254526 345440 254532
rect 343640 253224 343692 253230
rect 343640 253166 343692 253172
rect 342260 244928 342312 244934
rect 296902 244896 296958 244905
rect 342260 244870 342312 244876
rect 296902 244831 296958 244840
rect 355336 244118 355364 308654
rect 355428 308638 355548 308666
rect 355416 308576 355468 308582
rect 355416 308518 355468 308524
rect 355324 244112 355376 244118
rect 355324 244054 355376 244060
rect 355428 244050 355456 308518
rect 355520 306066 355548 308638
rect 355612 308310 355640 310420
rect 355600 308304 355652 308310
rect 355600 308246 355652 308252
rect 355888 306338 355916 310420
rect 356072 308038 356100 310420
rect 356152 308848 356204 308854
rect 356152 308790 356204 308796
rect 356164 308378 356192 308790
rect 356152 308372 356204 308378
rect 356152 308314 356204 308320
rect 356060 308032 356112 308038
rect 356060 307974 356112 307980
rect 355876 306332 355928 306338
rect 355876 306274 355928 306280
rect 355508 306060 355560 306066
rect 355508 306002 355560 306008
rect 356348 302734 356376 310420
rect 356532 308718 356560 310420
rect 356520 308712 356572 308718
rect 356520 308654 356572 308660
rect 356336 302728 356388 302734
rect 356336 302670 356388 302676
rect 356704 247580 356756 247586
rect 356704 247522 356756 247528
rect 356610 245304 356666 245313
rect 356610 245239 356666 245248
rect 356624 244633 356652 245239
rect 356610 244624 356666 244633
rect 356610 244559 356666 244568
rect 355416 244044 355468 244050
rect 355416 243986 355468 243992
rect 287428 243568 287480 243574
rect 287428 243510 287480 243516
rect 291200 243568 291252 243574
rect 291200 243510 291252 243516
rect 273350 159896 273406 159905
rect 273350 159831 273406 159840
rect 278134 159896 278190 159905
rect 278134 159831 278190 159840
rect 261114 159760 261170 159769
rect 261114 159695 261170 159704
rect 256700 159656 256752 159662
rect 256700 159598 256752 159604
rect 239588 158772 239640 158778
rect 239588 158714 239640 158720
rect 238116 158704 238168 158710
rect 220818 158672 220874 158681
rect 238114 158672 238116 158681
rect 239600 158681 239628 158714
rect 238168 158672 238170 158681
rect 220818 158607 220874 158616
rect 233240 158636 233292 158642
rect 219438 158400 219494 158409
rect 219438 158335 219494 158344
rect 219452 16574 219480 158335
rect 220832 16574 220860 158607
rect 238114 158607 238170 158616
rect 239586 158672 239642 158681
rect 239586 158607 239642 158616
rect 242438 158672 242494 158681
rect 242438 158607 242494 158616
rect 244646 158672 244702 158681
rect 244646 158607 244702 158616
rect 245566 158672 245622 158681
rect 245566 158607 245622 158616
rect 248326 158672 248382 158681
rect 248326 158607 248382 158616
rect 252374 158672 252430 158681
rect 252374 158607 252430 158616
rect 255870 158672 255926 158681
rect 255870 158607 255926 158616
rect 233240 158578 233292 158584
rect 224958 158536 225014 158545
rect 224958 158471 225014 158480
rect 223578 157992 223634 158001
rect 223578 157927 223634 157936
rect 219452 16546 220032 16574
rect 220832 16546 221136 16574
rect 219348 4004 219400 4010
rect 219348 3946 219400 3952
rect 219346 3632 219402 3641
rect 218058 3567 218114 3576
rect 219256 3596 219308 3602
rect 217508 3528 217560 3534
rect 216862 3496 216918 3505
rect 217508 3470 217560 3476
rect 216862 3431 216918 3440
rect 216586 3088 216642 3097
rect 216586 3023 216642 3032
rect 216876 480 216904 3431
rect 218072 480 218100 3567
rect 219346 3567 219402 3576
rect 219256 3538 219308 3544
rect 219254 3496 219310 3505
rect 219254 3431 219310 3440
rect 219268 480 219296 3431
rect 219360 3097 219388 3567
rect 219346 3088 219402 3097
rect 219346 3023 219402 3032
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 220452 4140 220504 4146
rect 220452 4082 220504 4088
rect 220464 4026 220492 4082
rect 220820 4072 220872 4078
rect 220464 4020 220820 4026
rect 220464 4014 220872 4020
rect 220464 3998 220860 4014
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 16546
rect 222750 3904 222806 3913
rect 222750 3839 222806 3848
rect 222764 480 222792 3839
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 157927
rect 224972 16574 225000 158471
rect 227718 158264 227774 158273
rect 227718 158199 227774 158208
rect 227732 16574 227760 158199
rect 230480 157956 230532 157962
rect 230480 157898 230532 157904
rect 229100 157888 229152 157894
rect 229100 157830 229152 157836
rect 229112 16574 229140 157830
rect 230492 16574 230520 157898
rect 231860 157820 231912 157826
rect 231860 157762 231912 157768
rect 224972 16546 225184 16574
rect 227732 16546 228312 16574
rect 229112 16546 229416 16574
rect 230492 16546 231072 16574
rect 225156 480 225184 16546
rect 227534 3768 227590 3777
rect 227534 3703 227590 3712
rect 226338 3224 226394 3233
rect 226338 3159 226394 3168
rect 226352 480 226380 3159
rect 227548 480 227576 3703
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 16546
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 16546
rect 231044 480 231072 16546
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 231872 354 231900 157762
rect 233252 16574 233280 158578
rect 238760 158568 238812 158574
rect 238760 158510 238812 158516
rect 237380 158500 237432 158506
rect 237380 158442 237432 158448
rect 234618 158128 234674 158137
rect 234618 158063 234674 158072
rect 233252 16546 233464 16574
rect 233436 480 233464 16546
rect 234632 11762 234660 158063
rect 234710 157992 234766 158001
rect 234710 157927 234766 157936
rect 234620 11756 234672 11762
rect 234620 11698 234672 11704
rect 234724 6914 234752 157927
rect 237392 16574 237420 158442
rect 238772 16574 238800 158510
rect 241520 158364 241572 158370
rect 241520 158306 241572 158312
rect 241426 158264 241482 158273
rect 241426 158199 241482 158208
rect 241440 155922 241468 158199
rect 241428 155916 241480 155922
rect 241428 155858 241480 155864
rect 241532 16574 241560 158306
rect 242452 157350 242480 158607
rect 242992 158432 243044 158438
rect 242992 158374 243044 158380
rect 242440 157344 242492 157350
rect 242440 157286 242492 157292
rect 243004 16574 243032 158374
rect 244660 157282 244688 158607
rect 244648 157276 244700 157282
rect 244648 157218 244700 157224
rect 245580 157146 245608 158607
rect 245660 158296 245712 158302
rect 245660 158238 245712 158244
rect 245568 157140 245620 157146
rect 245568 157082 245620 157088
rect 245672 16574 245700 158238
rect 247040 158228 247092 158234
rect 247040 158170 247092 158176
rect 246670 157992 246726 158001
rect 246670 157927 246726 157936
rect 246684 155854 246712 157927
rect 246672 155848 246724 155854
rect 246672 155790 246724 155796
rect 247052 16574 247080 158170
rect 247958 157992 248014 158001
rect 247958 157927 248014 157936
rect 247972 155718 248000 157927
rect 248340 157214 248368 158607
rect 248420 158160 248472 158166
rect 248420 158102 248472 158108
rect 248328 157208 248380 157214
rect 248328 157150 248380 157156
rect 247960 155712 248012 155718
rect 247960 155654 248012 155660
rect 237392 16546 237696 16574
rect 238772 16546 239352 16574
rect 241532 16546 241744 16574
rect 243004 16546 244136 16574
rect 245672 16546 245976 16574
rect 247052 16546 247632 16574
rect 235816 11756 235868 11762
rect 235816 11698 235868 11704
rect 234632 6886 234752 6914
rect 234632 480 234660 6886
rect 235828 480 235856 11698
rect 237010 3496 237066 3505
rect 237010 3431 237066 3440
rect 237024 480 237052 3431
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 237668 354 237696 16546
rect 239324 480 239352 16546
rect 240508 3256 240560 3262
rect 240508 3198 240560 3204
rect 240520 480 240548 3198
rect 241716 480 241744 16546
rect 242900 3324 242952 3330
rect 242900 3266 242952 3272
rect 242912 480 242940 3266
rect 244108 480 244136 16546
rect 245200 3392 245252 3398
rect 245200 3334 245252 3340
rect 245212 480 245240 3334
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 16546
rect 247604 480 247632 16546
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248432 354 248460 158102
rect 249800 158092 249852 158098
rect 249800 158034 249852 158040
rect 248694 157856 248750 157865
rect 248694 157791 248750 157800
rect 248708 155650 248736 157791
rect 248696 155644 248748 155650
rect 248696 155586 248748 155592
rect 249812 16574 249840 158034
rect 251086 157992 251142 158001
rect 251086 157927 251142 157936
rect 250442 157856 250498 157865
rect 250442 157791 250498 157800
rect 250456 155582 250484 157791
rect 251100 155786 251128 157927
rect 252388 157078 252416 158607
rect 252560 158024 252612 158030
rect 252560 157966 252612 157972
rect 252466 157856 252522 157865
rect 252466 157791 252522 157800
rect 252376 157072 252428 157078
rect 252376 157014 252428 157020
rect 251088 155780 251140 155786
rect 251088 155722 251140 155728
rect 250444 155576 250496 155582
rect 250444 155518 250496 155524
rect 252480 155514 252508 157791
rect 252468 155508 252520 155514
rect 252468 155450 252520 155456
rect 251180 155440 251232 155446
rect 251180 155382 251232 155388
rect 249812 16546 250024 16574
rect 249996 480 250024 16546
rect 251192 3398 251220 155382
rect 252572 16574 252600 157966
rect 253478 157856 253534 157865
rect 253478 157791 253534 157800
rect 253492 155446 253520 157791
rect 255884 157010 255912 158607
rect 256238 157584 256294 157593
rect 256238 157519 256294 157528
rect 255872 157004 255924 157010
rect 255872 156946 255924 156952
rect 253938 155952 253994 155961
rect 253938 155887 253994 155896
rect 253480 155440 253532 155446
rect 253480 155382 253532 155388
rect 253952 16574 253980 155887
rect 255318 155816 255374 155825
rect 255318 155751 255374 155760
rect 255332 16574 255360 155751
rect 256252 154562 256280 157519
rect 256240 154556 256292 154562
rect 256240 154498 256292 154504
rect 252572 16546 253520 16574
rect 253952 16546 254256 16574
rect 255332 16546 255912 16574
rect 251180 3392 251232 3398
rect 251180 3334 251232 3340
rect 252376 3392 252428 3398
rect 252376 3334 252428 3340
rect 251178 3224 251234 3233
rect 251178 3159 251234 3168
rect 251192 480 251220 3159
rect 252388 480 252416 3334
rect 253492 480 253520 16546
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 16546
rect 255884 480 255912 16546
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 256712 354 256740 159598
rect 260840 159520 260892 159526
rect 260840 159462 260892 159468
rect 257250 158672 257306 158681
rect 257250 158607 257306 158616
rect 257264 156942 257292 158607
rect 257252 156936 257304 156942
rect 257252 156878 257304 156884
rect 259550 155680 259606 155689
rect 259550 155615 259606 155624
rect 259564 6914 259592 155615
rect 260852 16574 260880 159462
rect 261128 158778 261156 159695
rect 263600 159588 263652 159594
rect 263600 159530 263652 159536
rect 261116 158772 261168 158778
rect 261116 158714 261168 158720
rect 261758 158672 261814 158681
rect 261758 158607 261814 158616
rect 261772 156874 261800 158607
rect 261760 156868 261812 156874
rect 261760 156810 261812 156816
rect 263612 16574 263640 159530
rect 264980 159452 265032 159458
rect 264980 159394 265032 159400
rect 263690 157584 263746 157593
rect 263690 157519 263746 157528
rect 263704 154494 263732 157519
rect 263692 154488 263744 154494
rect 263692 154430 263744 154436
rect 260852 16546 261800 16574
rect 263612 16546 264192 16574
rect 259472 6886 259592 6914
rect 258264 4140 258316 4146
rect 258264 4082 258316 4088
rect 258276 480 258304 4082
rect 259472 480 259500 6886
rect 260656 4072 260708 4078
rect 260656 4014 260708 4020
rect 260668 480 260696 4014
rect 261772 480 261800 16546
rect 262956 3936 263008 3942
rect 262956 3878 263008 3884
rect 262968 480 262996 3878
rect 264164 480 264192 16546
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 264992 354 265020 159394
rect 273364 158982 273392 159831
rect 275834 159624 275890 159633
rect 275834 159559 275890 159568
rect 277030 159624 277086 159633
rect 277030 159559 277086 159568
rect 273352 158976 273404 158982
rect 273352 158918 273404 158924
rect 275848 158914 275876 159559
rect 277044 159050 277072 159559
rect 278148 159118 278176 159831
rect 355322 159760 355378 159769
rect 351920 159724 351972 159730
rect 355322 159695 355378 159704
rect 351920 159666 351972 159672
rect 325884 159656 325936 159662
rect 279238 159624 279294 159633
rect 325884 159598 325936 159604
rect 279238 159559 279294 159568
rect 313280 159588 313332 159594
rect 279252 159186 279280 159559
rect 313280 159530 313332 159536
rect 310980 159520 311032 159526
rect 310980 159462 311032 159468
rect 291108 159452 291160 159458
rect 291108 159394 291160 159400
rect 284392 159384 284444 159390
rect 284392 159326 284444 159332
rect 285680 159384 285732 159390
rect 285680 159326 285732 159332
rect 279240 159180 279292 159186
rect 279240 159122 279292 159128
rect 278136 159112 278188 159118
rect 278136 159054 278188 159060
rect 277032 159044 277084 159050
rect 277032 158986 277084 158992
rect 275836 158908 275888 158914
rect 275836 158850 275888 158856
rect 274456 158840 274508 158846
rect 274456 158782 274508 158788
rect 269948 158704 270000 158710
rect 265438 158672 265494 158681
rect 265438 158607 265494 158616
rect 265990 158672 266046 158681
rect 265990 158607 266046 158616
rect 266542 158672 266598 158681
rect 266542 158607 266598 158616
rect 268750 158672 268806 158681
rect 268750 158607 268806 158616
rect 269946 158672 269948 158681
rect 274468 158681 274496 158782
rect 270000 158672 270002 158681
rect 269946 158607 270002 158616
rect 270958 158672 271014 158681
rect 270958 158607 271014 158616
rect 272246 158672 272302 158681
rect 272246 158607 272302 158616
rect 274454 158672 274510 158681
rect 274454 158607 274510 158616
rect 276110 158672 276166 158681
rect 276110 158607 276166 158616
rect 281078 158672 281134 158681
rect 281078 158607 281134 158616
rect 265452 157826 265480 158607
rect 265440 157820 265492 157826
rect 265440 157762 265492 157768
rect 266004 156806 266032 158607
rect 265992 156800 266044 156806
rect 265992 156742 266044 156748
rect 266556 156738 266584 158607
rect 268764 158166 268792 158607
rect 268752 158160 268804 158166
rect 268752 158102 268804 158108
rect 268382 157720 268438 157729
rect 268382 157655 268438 157664
rect 266544 156732 266596 156738
rect 266544 156674 266596 156680
rect 267830 155544 267886 155553
rect 267830 155479 267886 155488
rect 267740 155372 267792 155378
rect 267740 155314 267792 155320
rect 266544 4004 266596 4010
rect 266544 3946 266596 3952
rect 266556 480 266584 3946
rect 267752 480 267780 155314
rect 267844 16574 267872 155479
rect 268396 155378 268424 157655
rect 270972 156670 271000 158607
rect 272260 158574 272288 158607
rect 272248 158568 272300 158574
rect 272248 158510 272300 158516
rect 271326 157720 271382 157729
rect 271326 157655 271382 157664
rect 273718 157720 273774 157729
rect 273718 157655 273774 157664
rect 270960 156664 271012 156670
rect 270960 156606 271012 156612
rect 269118 155408 269174 155417
rect 268384 155372 268436 155378
rect 269118 155343 269174 155352
rect 268384 155314 268436 155320
rect 269132 16574 269160 155343
rect 271340 155242 271368 157655
rect 273732 155310 273760 157655
rect 276124 156602 276152 158607
rect 278502 157720 278558 157729
rect 278502 157655 278558 157664
rect 276112 156596 276164 156602
rect 276112 156538 276164 156544
rect 271880 155304 271932 155310
rect 271880 155246 271932 155252
rect 273720 155304 273772 155310
rect 273720 155246 273772 155252
rect 274638 155272 274694 155281
rect 270500 155236 270552 155242
rect 270500 155178 270552 155184
rect 271328 155236 271380 155242
rect 271328 155178 271380 155184
rect 270512 16574 270540 155178
rect 271892 16574 271920 155246
rect 274638 155207 274694 155216
rect 273260 152584 273312 152590
rect 273260 152526 273312 152532
rect 267844 16546 268424 16574
rect 269132 16546 270080 16574
rect 270512 16546 270816 16574
rect 271892 16546 272472 16574
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 16546
rect 270052 480 270080 16546
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 270788 354 270816 16546
rect 272444 480 272472 16546
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273272 354 273300 152526
rect 274652 16574 274680 155207
rect 278516 155174 278544 157655
rect 281092 156534 281120 158607
rect 283654 157584 283710 157593
rect 283654 157519 283710 157528
rect 281080 156528 281132 156534
rect 281080 156470 281132 156476
rect 277400 155168 277452 155174
rect 277400 155110 277452 155116
rect 278504 155168 278556 155174
rect 278504 155110 278556 155116
rect 276112 152652 276164 152658
rect 276112 152594 276164 152600
rect 276124 16574 276152 152594
rect 277412 16574 277440 155110
rect 283668 155106 283696 157519
rect 282920 155100 282972 155106
rect 282920 155042 282972 155048
rect 283656 155100 283708 155106
rect 283656 155042 283708 155048
rect 278780 155032 278832 155038
rect 278780 154974 278832 154980
rect 278792 16574 278820 154974
rect 282932 16574 282960 155042
rect 284404 16574 284432 159326
rect 285692 158574 285720 159326
rect 291120 158710 291148 159394
rect 291108 158704 291160 158710
rect 288254 158672 288310 158681
rect 288254 158607 288310 158616
rect 291014 158672 291070 158681
rect 295984 158704 296036 158710
rect 291108 158646 291160 158652
rect 293590 158672 293646 158681
rect 291014 158607 291070 158616
rect 293590 158607 293646 158616
rect 295982 158672 295984 158681
rect 296036 158672 296038 158681
rect 295982 158607 296038 158616
rect 298558 158672 298614 158681
rect 298558 158607 298614 158616
rect 300950 158672 301006 158681
rect 300950 158607 301006 158616
rect 303526 158672 303582 158681
rect 303526 158607 303582 158616
rect 306102 158672 306158 158681
rect 306102 158607 306158 158616
rect 308678 158672 308734 158681
rect 308678 158607 308734 158616
rect 285680 158568 285732 158574
rect 285680 158510 285732 158516
rect 288268 158098 288296 158607
rect 288256 158092 288308 158098
rect 288256 158034 288308 158040
rect 286046 157584 286102 157593
rect 286046 157519 286102 157528
rect 285680 156460 285732 156466
rect 285680 156402 285732 156408
rect 285692 16574 285720 156402
rect 286060 154426 286088 157519
rect 291028 156466 291056 158607
rect 293604 158574 293632 158607
rect 293592 158568 293644 158574
rect 293592 158510 293644 158516
rect 298572 158506 298600 158607
rect 298560 158500 298612 158506
rect 298560 158442 298612 158448
rect 300964 158438 300992 158607
rect 300952 158432 301004 158438
rect 300952 158374 301004 158380
rect 303540 158370 303568 158607
rect 303528 158364 303580 158370
rect 303528 158306 303580 158312
rect 306116 158302 306144 158607
rect 306104 158296 306156 158302
rect 306104 158238 306156 158244
rect 308692 158234 308720 158607
rect 308680 158228 308732 158234
rect 308680 158170 308732 158176
rect 310992 158166 311020 159462
rect 311070 158672 311126 158681
rect 311070 158607 311126 158616
rect 311084 158166 311112 158607
rect 310980 158160 311032 158166
rect 310980 158102 311032 158108
rect 311072 158160 311124 158166
rect 311072 158102 311124 158108
rect 313292 158098 313320 159530
rect 313462 158672 313518 158681
rect 313462 158607 313518 158616
rect 315854 158672 315910 158681
rect 315854 158607 315856 158616
rect 313476 158098 313504 158607
rect 315908 158607 315910 158616
rect 318614 158672 318670 158681
rect 318614 158607 318670 158616
rect 321006 158672 321062 158681
rect 321006 158607 321062 158616
rect 323398 158672 323454 158681
rect 323398 158607 323454 158616
rect 315856 158578 315908 158584
rect 313280 158092 313332 158098
rect 313280 158034 313332 158040
rect 313464 158092 313516 158098
rect 313464 158034 313516 158040
rect 318628 158030 318656 158607
rect 318616 158024 318668 158030
rect 318616 157966 318668 157972
rect 321020 157894 321048 158607
rect 323412 157962 323440 158607
rect 323400 157956 323452 157962
rect 323400 157898 323452 157904
rect 321008 157888 321060 157894
rect 321008 157830 321060 157836
rect 325896 157826 325924 159598
rect 325974 158672 326030 158681
rect 325974 158607 326030 158616
rect 325988 157826 326016 158607
rect 351932 158574 351960 159666
rect 355232 159112 355284 159118
rect 355232 159054 355284 159060
rect 355244 158914 355272 159054
rect 355232 158908 355284 158914
rect 355232 158850 355284 158856
rect 351920 158568 351972 158574
rect 351920 158510 351972 158516
rect 355336 157865 355364 159695
rect 355322 157856 355378 157865
rect 325884 157820 325936 157826
rect 325884 157762 325936 157768
rect 325976 157820 326028 157826
rect 355322 157791 355378 157800
rect 325976 157762 326028 157768
rect 291016 156460 291068 156466
rect 291016 156402 291068 156408
rect 286048 154420 286100 154426
rect 286048 154362 286100 154368
rect 288440 152516 288492 152522
rect 288440 152458 288492 152464
rect 288452 16574 288480 152458
rect 274652 16546 274864 16574
rect 276124 16546 276704 16574
rect 277412 16546 278360 16574
rect 278792 16546 279096 16574
rect 282932 16546 283144 16574
rect 284404 16546 284984 16574
rect 285692 16546 286640 16574
rect 288452 16546 289032 16574
rect 274836 480 274864 16546
rect 276020 3868 276072 3874
rect 276020 3810 276072 3816
rect 276032 480 276060 3810
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276676 354 276704 16546
rect 278332 480 278360 16546
rect 277094 354 277206 480
rect 276676 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 280712 3800 280764 3806
rect 280712 3742 280764 3748
rect 280724 480 280752 3742
rect 281908 3664 281960 3670
rect 281908 3606 281960 3612
rect 281920 480 281948 3606
rect 283116 480 283144 16546
rect 284300 3732 284352 3738
rect 284300 3674 284352 3680
rect 284312 480 284340 3674
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 284956 354 284984 16546
rect 286612 480 286640 16546
rect 287796 3596 287848 3602
rect 287796 3538 287848 3544
rect 287808 480 287836 3538
rect 289004 480 289032 16546
rect 300768 9648 300820 9654
rect 300768 9590 300820 9596
rect 296076 9172 296128 9178
rect 296076 9114 296128 9120
rect 294880 9036 294932 9042
rect 294880 8978 294932 8984
rect 293684 8968 293736 8974
rect 293684 8910 293736 8916
rect 292580 6180 292632 6186
rect 292580 6122 292632 6128
rect 291384 3528 291436 3534
rect 291384 3470 291436 3476
rect 290188 3460 290240 3466
rect 290188 3402 290240 3408
rect 290200 480 290228 3402
rect 291396 480 291424 3470
rect 292592 480 292620 6122
rect 293696 480 293724 8910
rect 294892 480 294920 8978
rect 296088 480 296116 9114
rect 299664 9104 299716 9110
rect 299664 9046 299716 9052
rect 298468 8900 298520 8906
rect 298468 8842 298520 8848
rect 297272 3460 297324 3466
rect 297272 3402 297324 3408
rect 297284 480 297312 3402
rect 298480 480 298508 8842
rect 299676 480 299704 9046
rect 300780 480 300808 9590
rect 301964 9580 302016 9586
rect 301964 9522 302016 9528
rect 301976 480 302004 9522
rect 309048 9512 309100 9518
rect 309048 9454 309100 9460
rect 306748 9444 306800 9450
rect 306748 9386 306800 9392
rect 305552 9376 305604 9382
rect 305552 9318 305604 9324
rect 304356 9308 304408 9314
rect 304356 9250 304408 9256
rect 303160 9240 303212 9246
rect 303160 9182 303212 9188
rect 303172 480 303200 9182
rect 304368 480 304396 9250
rect 305564 480 305592 9318
rect 306760 480 306788 9386
rect 307944 3528 307996 3534
rect 307944 3470 307996 3476
rect 307956 480 307984 3470
rect 309060 480 309088 9454
rect 322110 8936 322166 8945
rect 322110 8871 322166 8880
rect 312636 8832 312688 8838
rect 312636 8774 312688 8780
rect 311440 6316 311492 6322
rect 311440 6258 311492 6264
rect 310244 6248 310296 6254
rect 310244 6190 310296 6196
rect 310256 480 310284 6190
rect 311452 480 311480 6258
rect 312648 480 312676 8774
rect 316224 8764 316276 8770
rect 316224 8706 316276 8712
rect 313832 6656 313884 6662
rect 313832 6598 313884 6604
rect 313844 480 313872 6598
rect 315028 6384 315080 6390
rect 315028 6326 315080 6332
rect 315040 480 315068 6326
rect 316236 480 316264 8706
rect 319720 6588 319772 6594
rect 319720 6530 319772 6536
rect 318524 6520 318576 6526
rect 318524 6462 318576 6468
rect 317328 6452 317380 6458
rect 317328 6394 317380 6400
rect 317340 480 317368 6394
rect 318536 480 318564 6462
rect 319732 480 319760 6530
rect 320914 6216 320970 6225
rect 320914 6151 320970 6160
rect 320928 480 320956 6151
rect 322124 480 322152 8871
rect 330392 6860 330444 6866
rect 330392 6802 330444 6808
rect 323308 6724 323360 6730
rect 323308 6666 323360 6672
rect 323320 480 323348 6666
rect 326804 6112 326856 6118
rect 326804 6054 326856 6060
rect 325606 3496 325662 3505
rect 325606 3431 325662 3440
rect 324410 3360 324466 3369
rect 324410 3295 324466 3304
rect 324424 480 324452 3295
rect 325620 480 325648 3431
rect 326816 480 326844 6054
rect 329196 3664 329248 3670
rect 329196 3606 329248 3612
rect 328000 3596 328052 3602
rect 328000 3538 328052 3544
rect 328012 480 328040 3538
rect 329208 480 329236 3606
rect 330404 480 330432 6802
rect 333888 6792 333940 6798
rect 333888 6734 333940 6740
rect 351642 6760 351698 6769
rect 332692 3732 332744 3738
rect 332692 3674 332744 3680
rect 331586 3632 331642 3641
rect 331586 3567 331642 3576
rect 331600 480 331628 3567
rect 332704 480 332732 3674
rect 333900 480 333928 6734
rect 351642 6695 351698 6704
rect 348054 6624 348110 6633
rect 348054 6559 348110 6568
rect 346950 6488 347006 6497
rect 346950 6423 347006 6432
rect 344558 6352 344614 6361
rect 344558 6287 344614 6296
rect 337476 6044 337528 6050
rect 337476 5986 337528 5992
rect 336280 3800 336332 3806
rect 335082 3768 335138 3777
rect 336280 3742 336332 3748
rect 335082 3703 335138 3712
rect 335096 480 335124 3703
rect 336292 480 336320 3742
rect 337488 480 337516 5986
rect 340972 5976 341024 5982
rect 340972 5918 341024 5924
rect 338670 3904 338726 3913
rect 338670 3839 338726 3848
rect 339868 3868 339920 3874
rect 338684 480 338712 3839
rect 339868 3810 339920 3816
rect 339880 480 339908 3810
rect 340984 480 341012 5918
rect 342166 4040 342222 4049
rect 342166 3975 342222 3984
rect 342180 480 342208 3975
rect 343364 3936 343416 3942
rect 343364 3878 343416 3884
rect 343376 480 343404 3878
rect 344572 480 344600 6287
rect 345754 3224 345810 3233
rect 345754 3159 345810 3168
rect 345768 480 345796 3159
rect 346964 480 346992 6423
rect 348068 480 348096 6559
rect 350448 4072 350500 4078
rect 350448 4014 350500 4020
rect 349252 4004 349304 4010
rect 349252 3946 349304 3952
rect 349264 480 349292 3946
rect 350460 480 350488 4014
rect 351656 480 351684 6695
rect 355232 4140 355284 4146
rect 355232 4082 355284 4088
rect 352840 3392 352892 3398
rect 352840 3334 352892 3340
rect 352852 480 352880 3334
rect 354036 3324 354088 3330
rect 354036 3266 354088 3272
rect 354048 480 354076 3266
rect 355244 480 355272 4082
rect 356716 3534 356744 247522
rect 356808 159594 356836 310420
rect 356992 308922 357020 310420
rect 356888 308916 356940 308922
rect 356888 308858 356940 308864
rect 356980 308916 357032 308922
rect 356980 308858 357032 308864
rect 356900 244769 356928 308858
rect 357268 308802 357296 310420
rect 357466 310406 357664 310434
rect 357072 308780 357124 308786
rect 357268 308774 357388 308802
rect 357072 308722 357124 308728
rect 356980 308372 357032 308378
rect 356980 308314 357032 308320
rect 356886 244760 356942 244769
rect 356886 244695 356942 244704
rect 356992 244662 357020 308314
rect 357084 244866 357112 308722
rect 357256 308644 357308 308650
rect 357256 308586 357308 308592
rect 357164 308508 357216 308514
rect 357164 308450 357216 308456
rect 357072 244860 357124 244866
rect 357072 244802 357124 244808
rect 356980 244656 357032 244662
rect 356980 244598 357032 244604
rect 357176 244526 357204 308450
rect 357268 245546 357296 308586
rect 357360 305522 357388 308774
rect 357636 306354 357664 310406
rect 357728 306474 357756 310420
rect 357808 308440 357860 308446
rect 357808 308382 357860 308388
rect 357716 306468 357768 306474
rect 357716 306410 357768 306416
rect 357636 306326 357756 306354
rect 357624 306264 357676 306270
rect 357624 306206 357676 306212
rect 357348 305516 357400 305522
rect 357348 305458 357400 305464
rect 357440 250300 357492 250306
rect 357440 250242 357492 250248
rect 357452 248414 357480 250242
rect 357452 248386 357572 248414
rect 357440 245608 357492 245614
rect 357440 245550 357492 245556
rect 357256 245540 357308 245546
rect 357256 245482 357308 245488
rect 357452 245177 357480 245550
rect 357438 245168 357494 245177
rect 357438 245103 357494 245112
rect 357164 244520 357216 244526
rect 357164 244462 357216 244468
rect 356796 159588 356848 159594
rect 356796 159530 356848 159536
rect 357438 159352 357494 159361
rect 357438 159287 357494 159296
rect 356704 3528 356756 3534
rect 356704 3470 356756 3476
rect 357452 3482 357480 159287
rect 357544 6730 357572 248386
rect 357636 158778 357664 306206
rect 357728 159769 357756 306326
rect 357820 306134 357848 308382
rect 357808 306128 357860 306134
rect 357808 306070 357860 306076
rect 357912 302234 357940 310420
rect 358096 310406 358202 310434
rect 357992 306468 358044 306474
rect 357992 306410 358044 306416
rect 357820 302206 357940 302234
rect 357714 159760 357770 159769
rect 357714 159695 357770 159704
rect 357820 159662 357848 302206
rect 358004 296714 358032 306410
rect 358096 306270 358124 310406
rect 358372 308582 358400 310420
rect 358464 310406 358662 310434
rect 358360 308576 358412 308582
rect 358360 308518 358412 308524
rect 358268 308372 358320 308378
rect 358268 308314 358320 308320
rect 358176 307828 358228 307834
rect 358176 307770 358228 307776
rect 358084 306264 358136 306270
rect 358084 306206 358136 306212
rect 358084 306128 358136 306134
rect 358084 306070 358136 306076
rect 357912 296686 358032 296714
rect 357912 159730 357940 296686
rect 358096 245274 358124 306070
rect 357992 245268 358044 245274
rect 357992 245210 358044 245216
rect 358084 245268 358136 245274
rect 358084 245210 358136 245216
rect 357900 159724 357952 159730
rect 357900 159666 357952 159672
rect 357808 159656 357860 159662
rect 357808 159598 357860 159604
rect 357624 158772 357676 158778
rect 357624 158714 357676 158720
rect 357532 6724 357584 6730
rect 357532 6666 357584 6672
rect 358004 6254 358032 245210
rect 358084 243772 358136 243778
rect 358084 243714 358136 243720
rect 358096 9178 358124 243714
rect 358188 158370 358216 307770
rect 358176 158364 358228 158370
rect 358176 158306 358228 158312
rect 358280 158302 358308 308314
rect 358360 306468 358412 306474
rect 358360 306410 358412 306416
rect 358372 305998 358400 306410
rect 358360 305992 358412 305998
rect 358360 305934 358412 305940
rect 358464 296714 358492 310406
rect 358832 308446 358860 310420
rect 358924 310406 359122 310434
rect 358820 308440 358872 308446
rect 358820 308382 358872 308388
rect 358820 305992 358872 305998
rect 358820 305934 358872 305940
rect 358544 305924 358596 305930
rect 358544 305866 358596 305872
rect 358556 305726 358584 305866
rect 358544 305720 358596 305726
rect 358544 305662 358596 305668
rect 358728 305720 358780 305726
rect 358728 305662 358780 305668
rect 358740 305318 358768 305662
rect 358832 305454 358860 305934
rect 358820 305448 358872 305454
rect 358820 305390 358872 305396
rect 358728 305312 358780 305318
rect 358728 305254 358780 305260
rect 358372 296686 358492 296714
rect 358372 158506 358400 296686
rect 358820 250368 358872 250374
rect 358820 250310 358872 250316
rect 358360 158500 358412 158506
rect 358360 158442 358412 158448
rect 358268 158296 358320 158302
rect 358268 158238 358320 158244
rect 358084 9172 358136 9178
rect 358084 9114 358136 9120
rect 357992 6248 358044 6254
rect 357992 6190 358044 6196
rect 358832 6118 358860 250310
rect 358924 158438 358952 310406
rect 359004 309120 359056 309126
rect 359004 309062 359056 309068
rect 359016 308009 359044 309062
rect 359002 308000 359058 308009
rect 359002 307935 359058 307944
rect 359292 306354 359320 310420
rect 359464 308100 359516 308106
rect 359464 308042 359516 308048
rect 359016 306326 359320 306354
rect 359016 159526 359044 306326
rect 359476 306082 359504 308042
rect 359568 307834 359596 310420
rect 359648 308168 359700 308174
rect 359648 308110 359700 308116
rect 359556 307828 359608 307834
rect 359556 307770 359608 307776
rect 359384 306054 359504 306082
rect 359096 305448 359148 305454
rect 359096 305390 359148 305396
rect 359004 159520 359056 159526
rect 359004 159462 359056 159468
rect 359108 159458 359136 305390
rect 359188 248192 359240 248198
rect 359188 248134 359240 248140
rect 359096 159452 359148 159458
rect 359096 159394 359148 159400
rect 358912 158432 358964 158438
rect 358912 158374 358964 158380
rect 359200 6322 359228 248134
rect 359280 244044 359332 244050
rect 359280 243986 359332 243992
rect 359292 8906 359320 243986
rect 359384 158846 359412 306054
rect 359660 305130 359688 308110
rect 359752 305454 359780 310420
rect 360028 308378 360056 310420
rect 360016 308372 360068 308378
rect 360016 308314 360068 308320
rect 360212 308106 360240 310420
rect 360396 310406 360502 310434
rect 360200 308100 360252 308106
rect 360200 308042 360252 308048
rect 360108 307964 360160 307970
rect 360108 307906 360160 307912
rect 359832 307692 359884 307698
rect 359832 307634 359884 307640
rect 359740 305448 359792 305454
rect 359740 305390 359792 305396
rect 359464 305108 359516 305114
rect 359464 305050 359516 305056
rect 359568 305102 359688 305130
rect 359372 158840 359424 158846
rect 359372 158782 359424 158788
rect 359476 157894 359504 305050
rect 359568 158030 359596 305102
rect 359844 302234 359872 307634
rect 360016 306468 360068 306474
rect 360016 306410 360068 306416
rect 359924 306264 359976 306270
rect 359924 306206 359976 306212
rect 359936 306134 359964 306206
rect 359924 306128 359976 306134
rect 359924 306070 359976 306076
rect 360028 306066 360056 306410
rect 360016 306060 360068 306066
rect 360016 306002 360068 306008
rect 360120 305114 360148 307906
rect 360292 306468 360344 306474
rect 360292 306410 360344 306416
rect 360200 306400 360252 306406
rect 360200 306342 360252 306348
rect 360212 306270 360240 306342
rect 360200 306264 360252 306270
rect 360200 306206 360252 306212
rect 360108 305108 360160 305114
rect 360108 305050 360160 305056
rect 359660 302206 359872 302234
rect 359660 158098 359688 302206
rect 360200 251048 360252 251054
rect 360200 250990 360252 250996
rect 359648 158092 359700 158098
rect 359648 158034 359700 158040
rect 359556 158024 359608 158030
rect 359556 157966 359608 157972
rect 359464 157888 359516 157894
rect 359464 157830 359516 157836
rect 359280 8900 359332 8906
rect 359280 8842 359332 8848
rect 360212 6662 360240 250990
rect 360304 158166 360332 306410
rect 360396 158234 360424 310406
rect 360476 306400 360528 306406
rect 360476 306342 360528 306348
rect 360488 158982 360516 306342
rect 360672 296714 360700 310420
rect 360764 310406 360962 310434
rect 360764 306474 360792 310406
rect 360936 307896 360988 307902
rect 360936 307838 360988 307844
rect 360752 306468 360804 306474
rect 360752 306410 360804 306416
rect 360580 296686 360700 296714
rect 360580 159390 360608 296686
rect 360752 247988 360804 247994
rect 360752 247930 360804 247936
rect 360660 245336 360712 245342
rect 360660 245278 360712 245284
rect 360568 159384 360620 159390
rect 360568 159326 360620 159332
rect 360476 158976 360528 158982
rect 360476 158918 360528 158924
rect 360384 158228 360436 158234
rect 360384 158170 360436 158176
rect 360292 158160 360344 158166
rect 360292 158102 360344 158108
rect 360200 6656 360252 6662
rect 360200 6598 360252 6604
rect 359188 6316 359240 6322
rect 359188 6258 359240 6264
rect 358820 6112 358872 6118
rect 358820 6054 358872 6060
rect 360672 3602 360700 245278
rect 360764 8838 360792 247930
rect 360844 243704 360896 243710
rect 360844 243646 360896 243652
rect 360856 9654 360884 243646
rect 360948 157826 360976 307838
rect 361028 307828 361080 307834
rect 361028 307770 361080 307776
rect 361040 158914 361068 307770
rect 361132 306406 361160 310420
rect 361408 307698 361436 310420
rect 361488 309052 361540 309058
rect 361488 308994 361540 309000
rect 361500 307873 361528 308994
rect 361486 307864 361542 307873
rect 361592 307834 361620 310420
rect 361486 307799 361542 307808
rect 361580 307828 361632 307834
rect 361580 307770 361632 307776
rect 361396 307692 361448 307698
rect 361396 307634 361448 307640
rect 361120 306400 361172 306406
rect 361120 306342 361172 306348
rect 361580 254788 361632 254794
rect 361580 254730 361632 254736
rect 361118 159352 361174 159361
rect 361118 159287 361174 159296
rect 361028 158908 361080 158914
rect 361028 158850 361080 158856
rect 360936 157820 360988 157826
rect 360936 157762 360988 157768
rect 360844 9648 360896 9654
rect 360844 9590 360896 9596
rect 360752 8832 360804 8838
rect 360752 8774 360804 8780
rect 361132 6914 361160 159287
rect 361040 6886 361160 6914
rect 360660 3596 360712 3602
rect 360660 3538 360712 3544
rect 358726 3496 358782 3505
rect 357452 3454 357572 3482
rect 356336 3052 356388 3058
rect 356336 2994 356388 3000
rect 356348 480 356376 2994
rect 357544 480 357572 3454
rect 358726 3431 358782 3440
rect 359922 3496 359978 3505
rect 359922 3431 359978 3440
rect 358740 480 358768 3431
rect 359936 480 359964 3431
rect 361040 3330 361068 6886
rect 361118 3496 361174 3505
rect 361118 3431 361174 3440
rect 361028 3324 361080 3330
rect 361028 3266 361080 3272
rect 361132 480 361160 3431
rect 285374 354 285486 480
rect 284956 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 361592 354 361620 254730
rect 361672 253564 361724 253570
rect 361672 253506 361724 253512
rect 361684 6769 361712 253506
rect 361764 248396 361816 248402
rect 361764 248338 361816 248344
rect 361670 6760 361726 6769
rect 361670 6695 361726 6704
rect 361776 3670 361804 248338
rect 361868 158642 361896 310420
rect 362052 302234 362080 310420
rect 362328 308174 362356 310420
rect 362316 308168 362368 308174
rect 362316 308110 362368 308116
rect 361960 302206 362080 302234
rect 361960 159118 361988 302206
rect 362512 296714 362540 310420
rect 362788 307970 362816 310420
rect 362776 307964 362828 307970
rect 362776 307906 362828 307912
rect 363052 306400 363104 306406
rect 363052 306342 363104 306348
rect 362052 296686 362540 296714
rect 361948 159112 362000 159118
rect 361948 159054 362000 159060
rect 362052 159050 362080 296686
rect 362960 250436 363012 250442
rect 362960 250378 363012 250384
rect 362224 247920 362276 247926
rect 362224 247862 362276 247868
rect 362132 245472 362184 245478
rect 362132 245414 362184 245420
rect 362040 159044 362092 159050
rect 362040 158986 362092 158992
rect 361856 158636 361908 158642
rect 361856 158578 361908 158584
rect 361764 3664 361816 3670
rect 361764 3606 361816 3612
rect 362144 3058 362172 245414
rect 362236 6390 362264 247862
rect 362316 244520 362368 244526
rect 362316 244462 362368 244468
rect 362328 9110 362356 244462
rect 362408 244112 362460 244118
rect 362408 244054 362460 244060
rect 362420 9586 362448 244054
rect 362408 9580 362460 9586
rect 362408 9522 362460 9528
rect 362316 9104 362368 9110
rect 362316 9046 362368 9052
rect 362224 6384 362276 6390
rect 362224 6326 362276 6332
rect 362972 4078 363000 250378
rect 363064 157962 363092 306342
rect 363156 159186 363184 310542
rect 363248 306406 363276 310420
rect 363236 306400 363288 306406
rect 363236 306342 363288 306348
rect 363432 296714 363460 310420
rect 363708 307902 363736 310420
rect 365166 309088 365222 309097
rect 365166 309023 365222 309032
rect 363696 307896 363748 307902
rect 363696 307838 363748 307844
rect 363788 305584 363840 305590
rect 363788 305526 363840 305532
rect 363248 296686 363460 296714
rect 363248 159254 363276 296686
rect 363512 250776 363564 250782
rect 363512 250718 363564 250724
rect 363420 248328 363472 248334
rect 363420 248270 363472 248276
rect 363328 245404 363380 245410
rect 363328 245346 363380 245352
rect 363236 159248 363288 159254
rect 363236 159190 363288 159196
rect 363144 159180 363196 159186
rect 363144 159122 363196 159128
rect 363052 157956 363104 157962
rect 363052 157898 363104 157904
rect 362960 4072 363012 4078
rect 362960 4014 363012 4020
rect 363340 4010 363368 245346
rect 363432 6866 363460 248270
rect 363524 8770 363552 250718
rect 363696 244656 363748 244662
rect 363696 244598 363748 244604
rect 363604 243636 363656 243642
rect 363604 243578 363656 243584
rect 363512 8764 363564 8770
rect 363512 8706 363564 8712
rect 363420 6860 363472 6866
rect 363420 6802 363472 6808
rect 363328 4004 363380 4010
rect 363328 3946 363380 3952
rect 363510 3496 363566 3505
rect 363616 3466 363644 243578
rect 363708 6458 363736 244598
rect 363800 157146 363828 305526
rect 365076 305448 365128 305454
rect 365076 305390 365128 305396
rect 364708 251184 364760 251190
rect 364708 251126 364760 251132
rect 364616 248260 364668 248266
rect 364616 248202 364668 248208
rect 364432 248124 364484 248130
rect 364432 248066 364484 248072
rect 364340 247648 364392 247654
rect 364340 247590 364392 247596
rect 363878 159352 363934 159361
rect 363878 159287 363934 159296
rect 363788 157140 363840 157146
rect 363788 157082 363840 157088
rect 363696 6452 363748 6458
rect 363696 6394 363748 6400
rect 363510 3431 363566 3440
rect 363604 3460 363656 3466
rect 362132 3052 362184 3058
rect 362132 2994 362184 3000
rect 363524 480 363552 3431
rect 363604 3402 363656 3408
rect 363892 3398 363920 159287
rect 364352 3942 364380 247590
rect 364340 3936 364392 3942
rect 364340 3878 364392 3884
rect 364444 3738 364472 248066
rect 364524 248056 364576 248062
rect 364524 247998 364576 248004
rect 364536 3806 364564 247998
rect 364628 3874 364656 248202
rect 364720 6633 364748 251126
rect 364800 247512 364852 247518
rect 364800 247454 364852 247460
rect 364706 6624 364762 6633
rect 364706 6559 364762 6568
rect 364812 6497 364840 247454
rect 364892 244860 364944 244866
rect 364892 244802 364944 244808
rect 364904 6526 364932 244802
rect 364984 243568 365036 243574
rect 364984 243510 365036 243516
rect 364996 9246 365024 243510
rect 365088 155446 365116 305390
rect 365180 158545 365208 309023
rect 367284 308984 367336 308990
rect 367284 308926 367336 308932
rect 366456 308032 366508 308038
rect 366456 307974 366508 307980
rect 365720 268660 365772 268666
rect 365720 268602 365772 268608
rect 365166 158536 365222 158545
rect 365166 158471 365222 158480
rect 365076 155440 365128 155446
rect 365076 155382 365128 155388
rect 364984 9240 365036 9246
rect 364984 9182 365036 9188
rect 364892 6520 364944 6526
rect 364798 6488 364854 6497
rect 364892 6462 364944 6468
rect 364798 6423 364854 6432
rect 364616 3868 364668 3874
rect 364616 3810 364668 3816
rect 364524 3800 364576 3806
rect 364524 3742 364576 3748
rect 364432 3732 364484 3738
rect 364432 3674 364484 3680
rect 365732 3534 365760 268602
rect 365812 253496 365864 253502
rect 365812 253438 365864 253444
rect 365824 4146 365852 253438
rect 366180 251116 366232 251122
rect 366180 251058 366232 251064
rect 365904 250980 365956 250986
rect 365904 250922 365956 250928
rect 365916 5982 365944 250922
rect 366088 250912 366140 250918
rect 366088 250854 366140 250860
rect 365996 250708 366048 250714
rect 365996 250650 366048 250656
rect 366008 6594 366036 250650
rect 365996 6588 366048 6594
rect 365996 6530 366048 6536
rect 366100 6050 366128 250854
rect 366192 6361 366220 251058
rect 366272 250844 366324 250850
rect 366272 250786 366324 250792
rect 366284 6798 366312 250786
rect 366364 246696 366416 246702
rect 366364 246638 366416 246644
rect 366376 9314 366404 246638
rect 366468 159497 366496 307974
rect 366548 302796 366600 302802
rect 366548 302738 366600 302744
rect 366454 159488 366510 159497
rect 366454 159423 366510 159432
rect 366560 158273 366588 302738
rect 367100 247784 367152 247790
rect 367100 247726 367152 247732
rect 366546 158264 366602 158273
rect 366546 158199 366602 158208
rect 366364 9308 366416 9314
rect 366364 9250 366416 9256
rect 366272 6792 366324 6798
rect 366272 6734 366324 6740
rect 366178 6352 366234 6361
rect 366178 6287 366234 6296
rect 367112 6186 367140 247726
rect 367192 245200 367244 245206
rect 367192 245142 367244 245148
rect 367204 9382 367232 245142
rect 367296 157010 367324 308926
rect 367466 308816 367522 308825
rect 367466 308751 367522 308760
rect 367376 307828 367428 307834
rect 367376 307770 367428 307776
rect 367284 157004 367336 157010
rect 367284 156946 367336 156952
rect 367388 156942 367416 307770
rect 367480 157457 367508 308751
rect 367560 308236 367612 308242
rect 367560 308178 367612 308184
rect 367572 158409 367600 308178
rect 367652 302864 367704 302870
rect 367652 302806 367704 302812
rect 367558 158400 367614 158409
rect 367558 158335 367614 158344
rect 367466 157448 367522 157457
rect 367466 157383 367522 157392
rect 367376 156936 367428 156942
rect 367376 156878 367428 156884
rect 367664 154562 367692 302806
rect 367756 273222 367784 444926
rect 367834 308952 367890 308961
rect 367834 308887 367890 308896
rect 369124 308916 369176 308922
rect 367744 273216 367796 273222
rect 367744 273158 367796 273164
rect 367848 158817 367876 308887
rect 369124 308858 369176 308864
rect 368848 308576 368900 308582
rect 368848 308518 368900 308524
rect 367928 308304 367980 308310
rect 367928 308246 367980 308252
rect 368018 308272 368074 308281
rect 367940 159225 367968 308246
rect 368018 308207 368074 308216
rect 367926 159216 367982 159225
rect 367926 159151 367982 159160
rect 368032 159089 368060 308207
rect 368756 308100 368808 308106
rect 368756 308042 368808 308048
rect 368480 250640 368532 250646
rect 368480 250582 368532 250588
rect 368018 159080 368074 159089
rect 368018 159015 368074 159024
rect 367834 158808 367890 158817
rect 367834 158743 367890 158752
rect 367652 154556 367704 154562
rect 367652 154498 367704 154504
rect 368492 9450 368520 250582
rect 368664 247852 368716 247858
rect 368664 247794 368716 247800
rect 368572 247716 368624 247722
rect 368572 247658 368624 247664
rect 368480 9444 368532 9450
rect 368480 9386 368532 9392
rect 367192 9376 367244 9382
rect 367192 9318 367244 9324
rect 368584 8974 368612 247658
rect 368572 8968 368624 8974
rect 368676 8945 368704 247794
rect 368768 155242 368796 308042
rect 368860 156738 368888 308518
rect 369032 305992 369084 305998
rect 369032 305934 369084 305940
rect 368940 305788 368992 305794
rect 368940 305730 368992 305736
rect 368848 156732 368900 156738
rect 368848 156674 368900 156680
rect 368952 155718 368980 305730
rect 368940 155712 368992 155718
rect 368940 155654 368992 155660
rect 369044 155582 369072 305934
rect 369136 158137 369164 308858
rect 370042 308680 370098 308689
rect 370042 308615 370098 308624
rect 369216 306196 369268 306202
rect 369216 306138 369268 306144
rect 369122 158128 369178 158137
rect 369122 158063 369178 158072
rect 369228 157078 369256 306138
rect 369308 305652 369360 305658
rect 369308 305594 369360 305600
rect 369320 157214 369348 305594
rect 369860 245540 369912 245546
rect 369860 245482 369912 245488
rect 369308 157208 369360 157214
rect 369308 157150 369360 157156
rect 369216 157072 369268 157078
rect 369216 157014 369268 157020
rect 369032 155576 369084 155582
rect 369032 155518 369084 155524
rect 368756 155236 368808 155242
rect 368756 155178 368808 155184
rect 369872 9518 369900 245482
rect 369952 245268 370004 245274
rect 369952 245210 370004 245216
rect 369860 9512 369912 9518
rect 369860 9454 369912 9460
rect 369964 9042 369992 245210
rect 370056 157282 370084 308615
rect 370136 308576 370188 308582
rect 370136 308518 370188 308524
rect 370044 157276 370096 157282
rect 370044 157218 370096 157224
rect 370148 156874 370176 308518
rect 370504 308440 370556 308446
rect 370504 308382 370556 308388
rect 370226 306232 370282 306241
rect 370226 306167 370282 306176
rect 370136 156868 370188 156874
rect 370136 156810 370188 156816
rect 370240 155854 370268 306167
rect 370412 305924 370464 305930
rect 370412 305866 370464 305872
rect 370320 305720 370372 305726
rect 370320 305662 370372 305668
rect 370228 155848 370280 155854
rect 370228 155790 370280 155796
rect 370332 155650 370360 305662
rect 370320 155644 370372 155650
rect 370320 155586 370372 155592
rect 370424 155514 370452 305866
rect 370516 158001 370544 308382
rect 467838 308000 467894 308009
rect 467838 307935 467894 307944
rect 422300 307216 422352 307222
rect 422300 307158 422352 307164
rect 371424 306332 371476 306338
rect 371424 306274 371476 306280
rect 371332 306264 371384 306270
rect 371332 306206 371384 306212
rect 370688 303136 370740 303142
rect 370688 303078 370740 303084
rect 370596 302728 370648 302734
rect 370596 302670 370648 302676
rect 370502 157992 370558 158001
rect 370502 157927 370558 157936
rect 370412 155508 370464 155514
rect 370412 155450 370464 155456
rect 370608 154426 370636 302670
rect 370700 158953 370728 303078
rect 371240 287904 371292 287910
rect 371240 287846 371292 287852
rect 370686 158944 370742 158953
rect 370686 158879 370742 158888
rect 370596 154420 370648 154426
rect 370596 154362 370648 154368
rect 369952 9036 370004 9042
rect 369952 8978 370004 8984
rect 368572 8910 368624 8916
rect 368662 8936 368718 8945
rect 368662 8871 368718 8880
rect 367100 6180 367152 6186
rect 367100 6122 367152 6128
rect 366088 6044 366140 6050
rect 366088 5986 366140 5992
rect 365904 5976 365956 5982
rect 365904 5918 365956 5924
rect 365812 4140 365864 4146
rect 365812 4082 365864 4088
rect 365720 3528 365772 3534
rect 364614 3496 364670 3505
rect 367008 3528 367060 3534
rect 365720 3470 365772 3476
rect 365810 3496 365866 3505
rect 364614 3431 364670 3440
rect 367008 3470 367060 3476
rect 368202 3496 368258 3505
rect 365810 3431 365866 3440
rect 363880 3392 363932 3398
rect 363880 3334 363932 3340
rect 364628 480 364656 3431
rect 365824 480 365852 3431
rect 367020 480 367048 3470
rect 368202 3431 368258 3440
rect 369398 3496 369454 3505
rect 369398 3431 369454 3440
rect 370594 3496 370650 3505
rect 370594 3431 370650 3440
rect 368216 480 368244 3431
rect 369412 480 369440 3431
rect 370608 480 370636 3431
rect 362286 354 362398 480
rect 361592 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371252 354 371280 287846
rect 371344 155106 371372 306206
rect 371436 155174 371464 306274
rect 371884 306128 371936 306134
rect 371884 306070 371936 306076
rect 400218 306096 400274 306105
rect 371516 306060 371568 306066
rect 371516 306002 371568 306008
rect 371528 155310 371556 306002
rect 371792 305856 371844 305862
rect 371792 305798 371844 305804
rect 371700 305516 371752 305522
rect 371700 305458 371752 305464
rect 371608 303476 371660 303482
rect 371608 303418 371660 303424
rect 371516 155304 371568 155310
rect 371516 155246 371568 155252
rect 371424 155168 371476 155174
rect 371424 155110 371476 155116
rect 371332 155100 371384 155106
rect 371332 155042 371384 155048
rect 371620 154494 371648 303418
rect 371712 156466 371740 305458
rect 371804 156602 371832 305798
rect 371792 156596 371844 156602
rect 371792 156538 371844 156544
rect 371896 156534 371924 306070
rect 400218 306031 400274 306040
rect 390560 304428 390612 304434
rect 390560 304370 390612 304376
rect 372804 303612 372856 303618
rect 372804 303554 372856 303560
rect 371976 303408 372028 303414
rect 371976 303350 372028 303356
rect 371884 156528 371936 156534
rect 371884 156470 371936 156476
rect 371700 156460 371752 156466
rect 371700 156402 371752 156408
rect 371988 155786 372016 303350
rect 372712 303000 372764 303006
rect 372712 302942 372764 302948
rect 372620 300484 372672 300490
rect 372620 300426 372672 300432
rect 371976 155780 372028 155786
rect 371976 155722 372028 155728
rect 371608 154488 371660 154494
rect 371608 154430 371660 154436
rect 372632 16574 372660 300426
rect 372724 157350 372752 302942
rect 372712 157344 372764 157350
rect 372712 157286 372764 157292
rect 372816 156670 372844 303554
rect 372896 303544 372948 303550
rect 372896 303486 372948 303492
rect 372908 156806 372936 303486
rect 379520 303340 379572 303346
rect 379520 303282 379572 303288
rect 374276 303068 374328 303074
rect 374276 303010 374328 303016
rect 374184 302932 374236 302938
rect 374184 302874 374236 302880
rect 374000 287836 374052 287842
rect 374000 287778 374052 287784
rect 372896 156800 372948 156806
rect 372896 156742 372948 156748
rect 372804 156664 372856 156670
rect 372804 156606 372856 156612
rect 372632 16546 372936 16574
rect 372908 480 372936 16546
rect 374012 3534 374040 287778
rect 374092 270020 374144 270026
rect 374092 269962 374144 269968
rect 374000 3528 374052 3534
rect 374000 3470 374052 3476
rect 374104 480 374132 269962
rect 374196 155922 374224 302874
rect 374184 155916 374236 155922
rect 374184 155858 374236 155864
rect 374288 155378 374316 303010
rect 375380 301844 375432 301850
rect 375380 301786 375432 301792
rect 374276 155372 374328 155378
rect 374276 155314 374328 155320
rect 375392 16574 375420 301786
rect 378140 287768 378192 287774
rect 378140 287710 378192 287716
rect 376760 271380 376812 271386
rect 376760 271322 376812 271328
rect 376772 16574 376800 271322
rect 378152 16574 378180 287710
rect 375392 16546 376064 16574
rect 376772 16546 377720 16574
rect 378152 16546 378456 16574
rect 375288 3528 375340 3534
rect 375288 3470 375340 3476
rect 375300 480 375328 3470
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 16546
rect 377692 480 377720 16546
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378428 354 378456 16546
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 379532 354 379560 303282
rect 382280 303272 382332 303278
rect 382280 303214 382332 303220
rect 380900 271312 380952 271318
rect 380900 271254 380952 271260
rect 380912 16574 380940 271254
rect 380912 16546 381216 16574
rect 381188 480 381216 16546
rect 382292 3534 382320 303214
rect 386420 303204 386472 303210
rect 386420 303146 386472 303152
rect 382372 289332 382424 289338
rect 382372 289274 382424 289280
rect 382280 3528 382332 3534
rect 382280 3470 382332 3476
rect 382384 480 382412 289274
rect 383660 271244 383712 271250
rect 383660 271186 383712 271192
rect 383672 16574 383700 271186
rect 385684 254720 385736 254726
rect 385684 254662 385736 254668
rect 385040 250572 385092 250578
rect 385040 250514 385092 250520
rect 385052 16574 385080 250514
rect 383672 16546 384344 16574
rect 385052 16546 385632 16574
rect 383568 3528 383620 3534
rect 383568 3470 383620 3476
rect 383580 480 383608 3470
rect 379950 354 380062 480
rect 379532 326 380062 354
rect 378846 -960 378958 326
rect 379950 -960 380062 326
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 354 384344 16546
rect 385604 3482 385632 16546
rect 385696 3602 385724 254662
rect 386432 16574 386460 303146
rect 387800 272672 387852 272678
rect 387800 272614 387852 272620
rect 386432 16546 386736 16574
rect 385684 3596 385736 3602
rect 385684 3538 385736 3544
rect 385604 3454 386000 3482
rect 385972 480 386000 3454
rect 384734 354 384846 480
rect 384316 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 386708 354 386736 16546
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387812 354 387840 272614
rect 389180 250504 389232 250510
rect 389180 250446 389232 250452
rect 389192 16574 389220 250446
rect 389192 16546 389496 16574
rect 389468 480 389496 16546
rect 390572 3346 390600 304370
rect 392582 302832 392638 302841
rect 392582 302767 392638 302776
rect 391940 289264 391992 289270
rect 391940 289206 391992 289212
rect 390652 272604 390704 272610
rect 390652 272546 390704 272552
rect 390664 3534 390692 272546
rect 391952 6914 391980 289206
rect 392596 16574 392624 302767
rect 398840 290692 398892 290698
rect 398840 290634 398892 290640
rect 396080 289196 396132 289202
rect 396080 289138 396132 289144
rect 394700 272536 394752 272542
rect 394700 272478 394752 272484
rect 394712 16574 394740 272478
rect 392596 16546 392716 16574
rect 394712 16546 395384 16574
rect 391952 6886 392624 6914
rect 390652 3528 390704 3534
rect 390652 3470 390704 3476
rect 391848 3528 391900 3534
rect 391848 3470 391900 3476
rect 390572 3318 390692 3346
rect 390664 480 390692 3318
rect 391860 480 391888 3470
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 387126 -960 387238 326
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 6886
rect 392688 3534 392716 16546
rect 394238 3768 394294 3777
rect 394238 3703 394294 3712
rect 392676 3528 392728 3534
rect 392676 3470 392728 3476
rect 394252 480 394280 3703
rect 395356 480 395384 16546
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 289138
rect 397734 3632 397790 3641
rect 398852 3602 398880 290634
rect 398932 274168 398984 274174
rect 398932 274110 398984 274116
rect 397734 3567 397790 3576
rect 398840 3596 398892 3602
rect 397748 480 397776 3567
rect 398840 3538 398892 3544
rect 398944 480 398972 274110
rect 400232 16574 400260 306031
rect 404358 305960 404414 305969
rect 404358 305895 404414 305904
rect 402980 290624 403032 290630
rect 402980 290566 403032 290572
rect 401600 274100 401652 274106
rect 401600 274042 401652 274048
rect 401612 16574 401640 274042
rect 402992 16574 403020 290566
rect 400232 16546 400904 16574
rect 401612 16546 402560 16574
rect 402992 16546 403664 16574
rect 400128 3596 400180 3602
rect 400128 3538 400180 3544
rect 400140 480 400168 3538
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 16546
rect 402532 480 402560 16546
rect 403636 480 403664 16546
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 305895
rect 407118 305824 407174 305833
rect 407118 305759 407174 305768
rect 405740 246628 405792 246634
rect 405740 246570 405792 246576
rect 405752 16574 405780 246570
rect 405752 16546 406056 16574
rect 406028 480 406056 16546
rect 407132 2242 407160 305759
rect 418160 304360 418212 304366
rect 418160 304302 418212 304308
rect 409880 292052 409932 292058
rect 409880 291994 409932 292000
rect 407212 290556 407264 290562
rect 407212 290498 407264 290504
rect 407120 2236 407172 2242
rect 407120 2178 407172 2184
rect 407224 480 407252 290498
rect 408500 265872 408552 265878
rect 408500 265814 408552 265820
rect 408512 16574 408540 265814
rect 409892 16574 409920 291994
rect 414020 291984 414072 291990
rect 414020 291926 414072 291932
rect 412640 274032 412692 274038
rect 412640 273974 412692 273980
rect 408512 16546 409184 16574
rect 409892 16546 410840 16574
rect 408408 2236 408460 2242
rect 408408 2178 408460 2184
rect 408420 480 408448 2178
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 410812 480 410840 16546
rect 411902 3496 411958 3505
rect 411902 3431 411958 3440
rect 411916 480 411944 3431
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 273974
rect 414032 16574 414060 291926
rect 416780 282396 416832 282402
rect 416780 282338 416832 282344
rect 415492 275460 415544 275466
rect 415492 275402 415544 275408
rect 414032 16546 414336 16574
rect 414308 480 414336 16546
rect 415504 3534 415532 275402
rect 416792 6914 416820 282338
rect 417424 263084 417476 263090
rect 417424 263026 417476 263032
rect 417436 16574 417464 263026
rect 418172 16574 418200 304302
rect 420920 290488 420972 290494
rect 420920 290430 420972 290436
rect 419540 275392 419592 275398
rect 419540 275334 419592 275340
rect 419552 16574 419580 275334
rect 417436 16546 417556 16574
rect 418172 16546 418568 16574
rect 419552 16546 420224 16574
rect 416792 6886 417464 6914
rect 415492 3528 415544 3534
rect 415492 3470 415544 3476
rect 416688 3528 416740 3534
rect 416688 3470 416740 3476
rect 415492 3392 415544 3398
rect 415492 3334 415544 3340
rect 415504 480 415532 3334
rect 416700 480 416728 3470
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 6886
rect 417528 3466 417556 16546
rect 417516 3460 417568 3466
rect 417516 3402 417568 3408
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 418540 354 418568 16546
rect 420196 480 420224 16546
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 290430
rect 422312 16574 422340 307158
rect 458180 307148 458232 307154
rect 458180 307090 458232 307096
rect 429198 305688 429254 305697
rect 429198 305623 429254 305632
rect 427820 293480 427872 293486
rect 427820 293422 427872 293428
rect 423680 291916 423732 291922
rect 423680 291858 423732 291864
rect 422312 16546 422616 16574
rect 422588 480 422616 16546
rect 423692 3534 423720 291858
rect 426440 273964 426492 273970
rect 426440 273906 426492 273912
rect 423772 246492 423824 246498
rect 423772 246434 423824 246440
rect 423680 3528 423732 3534
rect 423680 3470 423732 3476
rect 423784 480 423812 246434
rect 426452 16574 426480 273906
rect 427832 16574 427860 293422
rect 426452 16546 426848 16574
rect 427832 16546 428504 16574
rect 426164 3596 426216 3602
rect 426164 3538 426216 3544
rect 424968 3528 425020 3534
rect 424968 3470 425020 3476
rect 424980 480 425008 3470
rect 426176 480 426204 3538
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 426820 354 426848 16546
rect 428476 480 428504 16546
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429212 354 429240 305623
rect 456800 300416 456852 300422
rect 456800 300358 456852 300364
rect 454040 298988 454092 298994
rect 454040 298930 454092 298936
rect 441620 293412 441672 293418
rect 441620 293354 441672 293360
rect 434720 291848 434772 291854
rect 434720 291790 434772 291796
rect 431960 283824 432012 283830
rect 431960 283766 432012 283772
rect 430580 246560 430632 246566
rect 430580 246502 430632 246508
rect 430592 16574 430620 246502
rect 430592 16546 430896 16574
rect 430868 480 430896 16546
rect 431972 3346 432000 283766
rect 433340 276888 433392 276894
rect 433340 276830 433392 276836
rect 432604 264444 432656 264450
rect 432604 264386 432656 264392
rect 432052 263016 432104 263022
rect 432052 262958 432104 262964
rect 432064 3534 432092 262958
rect 432616 3602 432644 264386
rect 433352 16574 433380 276830
rect 434732 16574 434760 291790
rect 437480 276820 437532 276826
rect 437480 276762 437532 276768
rect 436100 249280 436152 249286
rect 436100 249222 436152 249228
rect 436112 16574 436140 249222
rect 433352 16546 434024 16574
rect 434732 16546 435128 16574
rect 436112 16546 436784 16574
rect 432604 3596 432656 3602
rect 432604 3538 432656 3544
rect 432052 3528 432104 3534
rect 432052 3470 432104 3476
rect 433248 3528 433300 3534
rect 433248 3470 433300 3476
rect 431972 3318 432092 3346
rect 432064 480 432092 3318
rect 433260 480 433288 3470
rect 429630 354 429742 480
rect 429212 326 429742 354
rect 429630 -960 429742 326
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 16546
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 16546
rect 436756 480 436784 16546
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437492 354 437520 276762
rect 440884 265804 440936 265810
rect 440884 265746 440936 265752
rect 440240 264376 440292 264382
rect 440240 264318 440292 264324
rect 438858 250608 438914 250617
rect 438858 250543 438914 250552
rect 438872 16574 438900 250543
rect 438872 16546 439176 16574
rect 439148 480 439176 16546
rect 440252 3210 440280 264318
rect 440332 246424 440384 246430
rect 440332 246366 440384 246372
rect 440344 3398 440372 246366
rect 440896 3602 440924 265746
rect 441632 16574 441660 293354
rect 445760 287700 445812 287706
rect 445760 287642 445812 287648
rect 444380 271176 444432 271182
rect 444380 271118 444432 271124
rect 443000 254652 443052 254658
rect 443000 254594 443052 254600
rect 443012 16574 443040 254594
rect 444392 16574 444420 271118
rect 441632 16546 442672 16574
rect 443012 16546 443408 16574
rect 444392 16546 445064 16574
rect 440884 3596 440936 3602
rect 440884 3538 440936 3544
rect 440332 3392 440384 3398
rect 440332 3334 440384 3340
rect 441528 3392 441580 3398
rect 441528 3334 441580 3340
rect 440252 3182 440372 3210
rect 440344 480 440372 3182
rect 441540 480 441568 3334
rect 442644 480 442672 16546
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 354 443408 16546
rect 445036 480 445064 16546
rect 443798 354 443910 480
rect 443380 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 445772 354 445800 287642
rect 447140 286544 447192 286550
rect 447140 286486 447192 286492
rect 446404 265736 446456 265742
rect 446404 265678 446456 265684
rect 446416 3670 446444 265678
rect 447152 16574 447180 286486
rect 451280 276752 451332 276758
rect 451280 276694 451332 276700
rect 448520 275324 448572 275330
rect 448520 275266 448572 275272
rect 447152 16546 447456 16574
rect 446404 3664 446456 3670
rect 446404 3606 446456 3612
rect 447428 480 447456 16546
rect 448532 3210 448560 275266
rect 449900 269952 449952 269958
rect 449900 269894 449952 269900
rect 448612 252068 448664 252074
rect 448612 252010 448664 252016
rect 448624 3398 448652 252010
rect 449912 16574 449940 269894
rect 451292 16574 451320 276694
rect 452660 252000 452712 252006
rect 452660 251942 452712 251948
rect 452672 16574 452700 251942
rect 449912 16546 450952 16574
rect 451292 16546 451688 16574
rect 452672 16546 453344 16574
rect 448612 3392 448664 3398
rect 448612 3334 448664 3340
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 448532 3182 448652 3210
rect 448624 480 448652 3182
rect 449820 480 449848 3334
rect 450924 480 450952 16546
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 453316 480 453344 16546
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454052 354 454080 298930
rect 455420 278248 455472 278254
rect 455420 278190 455472 278196
rect 455432 16574 455460 278190
rect 455432 16546 455736 16574
rect 455708 480 455736 16546
rect 456812 3398 456840 300358
rect 456892 251932 456944 251938
rect 456892 251874 456944 251880
rect 456800 3392 456852 3398
rect 456800 3334 456852 3340
rect 456904 480 456932 251874
rect 458192 16574 458220 307090
rect 463700 294840 463752 294846
rect 463700 294782 463752 294788
rect 459560 293344 459612 293350
rect 459560 293286 459612 293292
rect 459572 16574 459600 293286
rect 462320 278180 462372 278186
rect 462320 278122 462372 278128
rect 460940 256216 460992 256222
rect 460940 256158 460992 256164
rect 460952 16574 460980 256158
rect 458192 16546 459232 16574
rect 459572 16546 459968 16574
rect 460952 16546 461624 16574
rect 458088 3392 458140 3398
rect 458088 3334 458140 3340
rect 458100 480 458128 3334
rect 459204 480 459232 16546
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 461596 480 461624 16546
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462332 354 462360 278122
rect 463712 16574 463740 294782
rect 465080 256148 465132 256154
rect 465080 256090 465132 256096
rect 463712 16546 464016 16574
rect 463988 480 464016 16546
rect 465092 6914 465120 256090
rect 466460 251864 466512 251870
rect 466460 251806 466512 251812
rect 465170 248024 465226 248033
rect 465170 247959 465226 247968
rect 465184 16574 465212 247959
rect 466472 16574 466500 251806
rect 467852 16574 467880 307935
rect 471978 307864 472034 307873
rect 471978 307799 472034 307808
rect 470600 289128 470652 289134
rect 470600 289070 470652 289076
rect 469218 247888 469274 247897
rect 469218 247823 469274 247832
rect 469232 16574 469260 247823
rect 465184 16546 465856 16574
rect 466472 16546 467512 16574
rect 467852 16546 468248 16574
rect 469232 16546 469904 16574
rect 465092 6886 465212 6914
rect 465184 480 465212 6886
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 354 465856 16546
rect 467484 480 467512 16546
rect 466246 354 466358 480
rect 465828 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468220 354 468248 16546
rect 469876 480 469904 16546
rect 468638 354 468750 480
rect 468220 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 470612 354 470640 289070
rect 471992 16574 472020 307799
rect 480260 307080 480312 307086
rect 480260 307022 480312 307028
rect 473360 294772 473412 294778
rect 473360 294714 473412 294720
rect 471992 16546 472296 16574
rect 472268 480 472296 16546
rect 473372 3398 473400 294714
rect 477500 293276 477552 293282
rect 477500 293218 477552 293224
rect 474740 256080 474792 256086
rect 474740 256022 474792 256028
rect 473450 247752 473506 247761
rect 473450 247687 473506 247696
rect 473360 3392 473412 3398
rect 473360 3334 473412 3340
rect 473464 480 473492 247687
rect 474752 16574 474780 256022
rect 476118 247616 476174 247625
rect 476118 247551 476174 247560
rect 476132 16574 476160 247551
rect 477512 16574 477540 293218
rect 478880 256012 478932 256018
rect 478880 255954 478932 255960
rect 474752 16546 475792 16574
rect 476132 16546 476528 16574
rect 477512 16546 478184 16574
rect 474188 3392 474240 3398
rect 474188 3334 474240 3340
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474200 354 474228 3334
rect 475764 480 475792 16546
rect 474526 354 474638 480
rect 474200 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476500 354 476528 16546
rect 478156 480 478184 16546
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 478892 354 478920 255954
rect 480272 16574 480300 307022
rect 542360 300280 542412 300286
rect 542360 300222 542412 300228
rect 531320 298920 531372 298926
rect 531320 298862 531372 298868
rect 503720 297628 503772 297634
rect 503720 297570 503772 297576
rect 489920 296200 489972 296206
rect 489920 296142 489972 296148
rect 481640 294704 481692 294710
rect 481640 294646 481692 294652
rect 480272 16546 480576 16574
rect 480548 480 480576 16546
rect 481652 3398 481680 294646
rect 485780 285184 485832 285190
rect 485780 285126 485832 285132
rect 484400 279676 484452 279682
rect 484400 279618 484452 279624
rect 481732 278112 481784 278118
rect 481732 278054 481784 278060
rect 481640 3392 481692 3398
rect 481640 3334 481692 3340
rect 481744 480 481772 278054
rect 483020 260228 483072 260234
rect 483020 260170 483072 260176
rect 483032 16574 483060 260170
rect 484412 16574 484440 279618
rect 485792 16574 485820 285126
rect 488540 278044 488592 278050
rect 488540 277986 488592 277992
rect 487160 261724 487212 261730
rect 487160 261666 487212 261672
rect 483032 16546 484072 16574
rect 484412 16546 484808 16574
rect 485792 16546 486464 16574
rect 482468 3392 482520 3398
rect 482468 3334 482520 3340
rect 479310 354 479422 480
rect 478892 326 479422 354
rect 479310 -960 479422 326
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482480 354 482508 3334
rect 484044 480 484072 16546
rect 482806 354 482918 480
rect 482480 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 486436 480 486464 16546
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487172 354 487200 261666
rect 488552 16574 488580 277986
rect 488552 16546 488856 16574
rect 488828 480 488856 16546
rect 489932 480 489960 296142
rect 492680 296132 492732 296138
rect 492680 296074 492732 296080
rect 491300 279608 491352 279614
rect 491300 279550 491352 279556
rect 490012 261656 490064 261662
rect 490012 261598 490064 261604
rect 490024 16574 490052 261598
rect 491312 16574 491340 279550
rect 492692 16574 492720 296074
rect 499580 296064 499632 296070
rect 499580 296006 499632 296012
rect 498200 281036 498252 281042
rect 498200 280978 498252 280984
rect 495440 279540 495492 279546
rect 495440 279482 495492 279488
rect 494060 261588 494112 261594
rect 494060 261530 494112 261536
rect 494072 16574 494100 261530
rect 490024 16546 490696 16574
rect 491312 16546 492352 16574
rect 492692 16546 493088 16574
rect 494072 16546 494744 16574
rect 487590 354 487702 480
rect 487172 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490668 354 490696 16546
rect 492324 480 492352 16546
rect 491086 354 491198 480
rect 490668 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 494716 480 494744 16546
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 279482
rect 496084 267232 496136 267238
rect 496084 267174 496136 267180
rect 496096 3874 496124 267174
rect 496820 246356 496872 246362
rect 496820 246298 496872 246304
rect 496832 16574 496860 246298
rect 496832 16546 497136 16574
rect 496084 3868 496136 3874
rect 496084 3810 496136 3816
rect 497108 480 497136 16546
rect 498212 3398 498240 280978
rect 498292 262948 498344 262954
rect 498292 262890 498344 262896
rect 498200 3392 498252 3398
rect 498200 3334 498252 3340
rect 498304 3210 498332 262890
rect 499592 16574 499620 296006
rect 502984 267164 503036 267170
rect 502984 267106 503036 267112
rect 502340 245132 502392 245138
rect 502340 245074 502392 245080
rect 499592 16546 500632 16574
rect 499028 3392 499080 3398
rect 499028 3334 499080 3340
rect 498212 3182 498332 3210
rect 498212 480 498240 3182
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499040 354 499068 3334
rect 500604 480 500632 16546
rect 502352 6914 502380 245074
rect 502996 16574 503024 267106
rect 502996 16546 503116 16574
rect 502352 6886 503024 6914
rect 501786 3360 501842 3369
rect 501786 3295 501842 3304
rect 501800 480 501828 3295
rect 502996 480 503024 6886
rect 503088 3942 503116 16546
rect 503076 3936 503128 3942
rect 503076 3878 503128 3884
rect 499366 354 499478 480
rect 499040 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503732 354 503760 297570
rect 506480 297560 506532 297566
rect 506480 297502 506532 297508
rect 506492 3466 506520 297502
rect 510620 297492 510672 297498
rect 510620 297434 510672 297440
rect 506572 280968 506624 280974
rect 506572 280910 506624 280916
rect 505376 3460 505428 3466
rect 505376 3402 505428 3408
rect 506480 3460 506532 3466
rect 506480 3402 506532 3408
rect 505388 480 505416 3402
rect 506584 3346 506612 280910
rect 509240 280900 509292 280906
rect 509240 280842 509292 280848
rect 508504 268592 508556 268598
rect 508504 268534 508556 268540
rect 507860 264308 507912 264314
rect 507860 264250 507912 264256
rect 507872 16574 507900 264250
rect 507872 16546 508452 16574
rect 508424 3482 508452 16546
rect 508516 3738 508544 268534
rect 509252 16574 509280 280842
rect 510632 16574 510660 297434
rect 528560 294636 528612 294642
rect 528560 294578 528612 294584
rect 516140 282328 516192 282334
rect 516140 282270 516192 282276
rect 513380 276684 513432 276690
rect 513380 276626 513432 276632
rect 512000 264240 512052 264246
rect 512000 264182 512052 264188
rect 509252 16546 509648 16574
rect 510632 16546 511304 16574
rect 508504 3732 508556 3738
rect 508504 3674 508556 3680
rect 507308 3460 507360 3466
rect 508424 3454 508912 3482
rect 507308 3402 507360 3408
rect 506492 3318 506612 3346
rect 506492 480 506520 3318
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507320 354 507348 3402
rect 508884 480 508912 3454
rect 507646 354 507758 480
rect 507320 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 511276 480 511304 16546
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 264182
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 513392 354 513420 276626
rect 514852 268456 514904 268462
rect 514852 268398 514904 268404
rect 514864 6914 514892 268398
rect 516152 16574 516180 282270
rect 520280 282260 520332 282266
rect 520280 282202 520332 282208
rect 516784 268524 516836 268530
rect 516784 268466 516836 268472
rect 516152 16546 516732 16574
rect 514772 6886 514892 6914
rect 514772 480 514800 6886
rect 515956 3528 516008 3534
rect 515956 3470 516008 3476
rect 516704 3482 516732 16546
rect 516796 3806 516824 268466
rect 517520 253428 517572 253434
rect 517520 253370 517572 253376
rect 517532 16574 517560 253370
rect 517532 16546 517928 16574
rect 516784 3800 516836 3806
rect 516784 3742 516836 3748
rect 515968 480 515996 3470
rect 516704 3454 517192 3482
rect 517164 480 517192 3454
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512430 -960 512542 326
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 519544 3596 519596 3602
rect 519544 3538 519596 3544
rect 519556 480 519584 3538
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 282202
rect 527180 282192 527232 282198
rect 527180 282134 527232 282140
rect 520924 269884 520976 269890
rect 520924 269826 520976 269832
rect 520936 3466 520964 269826
rect 525064 269816 525116 269822
rect 525064 269758 525116 269764
rect 523132 267096 523184 267102
rect 523132 267038 523184 267044
rect 521660 253360 521712 253366
rect 521660 253302 521712 253308
rect 520924 3460 520976 3466
rect 520924 3402 520976 3408
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 253302
rect 523144 16574 523172 267038
rect 524420 253292 524472 253298
rect 524420 253234 524472 253240
rect 524432 16574 524460 253234
rect 523144 16546 523816 16574
rect 524432 16546 525012 16574
rect 523040 3664 523092 3670
rect 523040 3606 523092 3612
rect 523052 480 523080 3606
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523788 354 523816 16546
rect 524984 3482 525012 16546
rect 525076 3602 525104 269758
rect 525800 265668 525852 265674
rect 525800 265610 525852 265616
rect 525812 16574 525840 265610
rect 527192 16574 527220 282134
rect 525812 16546 526208 16574
rect 527192 16546 527864 16574
rect 525064 3596 525116 3602
rect 525064 3538 525116 3544
rect 524984 3454 525472 3482
rect 525444 480 525472 3454
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527836 480 527864 16546
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 294578
rect 529940 260160 529992 260166
rect 529940 260102 529992 260108
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 260102
rect 531332 3602 531360 298862
rect 535460 298852 535512 298858
rect 535460 298794 535512 298800
rect 531412 283756 531464 283762
rect 531412 283698 531464 283704
rect 531320 3596 531372 3602
rect 531320 3538 531372 3544
rect 531424 3482 531452 283698
rect 534724 249212 534776 249218
rect 534724 249154 534776 249160
rect 534080 249144 534132 249150
rect 534080 249086 534132 249092
rect 534092 16574 534120 249086
rect 534092 16546 534488 16574
rect 533712 3868 533764 3874
rect 533712 3810 533764 3816
rect 532148 3596 532200 3602
rect 532148 3538 532200 3544
rect 531332 3454 531452 3482
rect 531332 480 531360 3454
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532160 354 532188 3538
rect 533724 480 533752 3810
rect 532486 354 532598 480
rect 532160 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 534736 3602 534764 249154
rect 535472 16574 535500 298794
rect 539600 298784 539652 298790
rect 539600 298726 539652 298732
rect 538864 285116 538916 285122
rect 538864 285058 538916 285064
rect 538220 249076 538272 249082
rect 538220 249018 538272 249024
rect 535472 16546 536144 16574
rect 534724 3596 534776 3602
rect 534724 3538 534776 3544
rect 536116 480 536144 16546
rect 537208 3936 537260 3942
rect 537208 3878 537260 3884
rect 537220 480 537248 3878
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 249018
rect 538876 3874 538904 285058
rect 538864 3868 538916 3874
rect 538864 3810 538916 3816
rect 539612 480 539640 298726
rect 539692 267028 539744 267034
rect 539692 266970 539744 266976
rect 539704 16574 539732 266970
rect 542372 16574 542400 300222
rect 549260 300212 549312 300218
rect 549260 300154 549312 300160
rect 543004 286476 543056 286482
rect 543004 286418 543056 286424
rect 539704 16546 540376 16574
rect 542372 16546 542768 16574
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540348 354 540376 16546
rect 541992 3596 542044 3602
rect 541992 3538 542044 3544
rect 542004 480 542032 3538
rect 540766 354 540878 480
rect 540348 326 540878 354
rect 540766 -960 540878 326
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 543016 3670 543044 286418
rect 547880 283688 547932 283694
rect 547880 283630 547932 283636
rect 545120 279472 545172 279478
rect 545120 279414 545172 279420
rect 543740 261520 543792 261526
rect 543740 261462 543792 261468
rect 543752 16574 543780 261462
rect 545132 16574 545160 279414
rect 546498 250472 546554 250481
rect 546498 250407 546554 250416
rect 543752 16546 544424 16574
rect 545132 16546 545528 16574
rect 543004 3664 543056 3670
rect 543004 3606 543056 3612
rect 544396 480 544424 16546
rect 545500 480 545528 16546
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 250407
rect 547892 3602 547920 283630
rect 547972 268388 548024 268394
rect 547972 268330 548024 268336
rect 547880 3596 547932 3602
rect 547880 3538 547932 3544
rect 547984 3482 548012 268330
rect 549272 16574 549300 300154
rect 553400 300144 553452 300150
rect 553400 300086 553452 300092
rect 552664 286408 552716 286414
rect 552664 286350 552716 286356
rect 552020 283620 552072 283626
rect 552020 283562 552072 283568
rect 549272 16546 550312 16574
rect 548708 3596 548760 3602
rect 548708 3538 548760 3544
rect 547892 3454 548012 3482
rect 547892 480 547920 3454
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 548720 354 548748 3538
rect 550284 480 550312 16546
rect 552032 6914 552060 283562
rect 552676 16574 552704 286350
rect 553412 16574 553440 300086
rect 552676 16546 552796 16574
rect 553412 16546 553808 16574
rect 552032 6886 552704 6914
rect 551468 3732 551520 3738
rect 551468 3674 551520 3680
rect 551480 480 551508 3674
rect 552572 3664 552624 3670
rect 552572 3606 552624 3612
rect 552584 3398 552612 3606
rect 552572 3392 552624 3398
rect 552572 3334 552624 3340
rect 552676 480 552704 6886
rect 552768 3806 552796 16546
rect 552756 3800 552808 3806
rect 552756 3742 552808 3748
rect 553780 480 553808 16546
rect 554056 3738 554084 445839
rect 556160 295996 556212 296002
rect 556160 295938 556212 295944
rect 554044 3732 554096 3738
rect 554044 3674 554096 3680
rect 556172 3602 556200 295938
rect 556252 280832 556304 280838
rect 556252 280774 556304 280780
rect 554964 3596 555016 3602
rect 554964 3538 555016 3544
rect 556160 3596 556212 3602
rect 556160 3538 556212 3544
rect 554976 480 555004 3538
rect 556264 3482 556292 280774
rect 557540 245064 557592 245070
rect 557540 245006 557592 245012
rect 557552 16574 557580 245006
rect 557552 16546 558132 16574
rect 557172 3664 557224 3670
rect 557172 3606 557224 3612
rect 556988 3596 557040 3602
rect 556988 3538 557040 3544
rect 556172 3454 556292 3482
rect 556172 480 556200 3454
rect 549046 354 549158 480
rect 548720 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557000 354 557028 3538
rect 557184 3398 557212 3606
rect 558104 3482 558132 16546
rect 558196 3806 558224 446111
rect 580632 445188 580684 445194
rect 580632 445130 580684 445136
rect 580540 445120 580592 445126
rect 580540 445062 580592 445068
rect 580448 445052 580500 445058
rect 580448 444994 580500 445000
rect 580356 443080 580408 443086
rect 580356 443022 580408 443028
rect 580264 443012 580316 443018
rect 580264 442954 580316 442960
rect 580172 431928 580224 431934
rect 580172 431870 580224 431876
rect 580184 431633 580212 431870
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 579620 379500 579672 379506
rect 579620 379442 579672 379448
rect 579632 378457 579660 379442
rect 579618 378448 579674 378457
rect 579618 378383 579674 378392
rect 579988 325644 580040 325650
rect 579988 325586 580040 325592
rect 580000 325281 580028 325586
rect 579986 325272 580042 325281
rect 579986 325207 580042 325216
rect 560300 301640 560352 301646
rect 560300 301582 560352 301588
rect 560312 16574 560340 301582
rect 564440 301572 564492 301578
rect 564440 301514 564492 301520
rect 563060 285048 563112 285054
rect 563060 284990 563112 284996
rect 561680 244996 561732 245002
rect 561680 244938 561732 244944
rect 561692 16574 561720 244938
rect 560312 16546 560432 16574
rect 561692 16546 562088 16574
rect 559748 3868 559800 3874
rect 559748 3810 559800 3816
rect 558184 3800 558236 3806
rect 558184 3742 558236 3748
rect 558104 3454 558592 3482
rect 557172 3392 557224 3398
rect 557172 3334 557224 3340
rect 558564 480 558592 3454
rect 559760 480 559788 3810
rect 557326 354 557438 480
rect 557000 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560404 354 560432 16546
rect 562060 480 562088 16546
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563072 354 563100 284990
rect 564452 480 564480 301514
rect 574100 301504 574152 301510
rect 574100 301446 574152 301452
rect 567200 297424 567252 297430
rect 567200 297366 567252 297372
rect 565820 284980 565872 284986
rect 565820 284922 565872 284928
rect 564532 244928 564584 244934
rect 564532 244870 564584 244876
rect 564544 16574 564572 244870
rect 565832 16574 565860 284922
rect 567212 16574 567240 297366
rect 569960 286340 570012 286346
rect 569960 286282 570012 286288
rect 569972 16574 570000 286282
rect 571340 253224 571392 253230
rect 571340 253166 571392 253172
rect 564544 16546 565216 16574
rect 565832 16546 566872 16574
rect 567212 16546 567608 16574
rect 569972 16546 570368 16574
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565188 354 565216 16546
rect 566844 480 566872 16546
rect 565606 354 565718 480
rect 565188 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 569132 3460 569184 3466
rect 569132 3402 569184 3408
rect 569144 480 569172 3402
rect 570340 480 570368 16546
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 567998 -960 568110 326
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571352 354 571380 253166
rect 574112 16574 574140 301446
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 575480 262880 575532 262886
rect 575480 262822 575532 262828
rect 575492 16574 575520 262822
rect 578240 254584 578292 254590
rect 578240 254526 578292 254532
rect 578252 16574 578280 254526
rect 580276 33153 580304 442954
rect 580368 112849 580396 443022
rect 580460 152697 580488 444994
rect 580552 192545 580580 445062
rect 580644 232393 580672 445130
rect 580630 232384 580686 232393
rect 580630 232319 580686 232328
rect 580538 192536 580594 192545
rect 580538 192471 580594 192480
rect 581090 177304 581146 177313
rect 581090 177239 581146 177248
rect 580446 152688 580502 152697
rect 580446 152623 580502 152632
rect 580354 112840 580410 112849
rect 580354 112775 580410 112784
rect 580262 33144 580318 33153
rect 580262 33079 580318 33088
rect 574112 16546 575152 16574
rect 575492 16546 575888 16574
rect 578252 16546 578648 16574
rect 573916 3664 573968 3670
rect 573916 3606 573968 3612
rect 572720 3528 572772 3534
rect 572720 3470 572772 3476
rect 572732 480 572760 3470
rect 573928 480 573956 3606
rect 575124 480 575152 16546
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 575860 354 575888 16546
rect 577412 3732 577464 3738
rect 577412 3674 577464 3680
rect 577424 480 577452 3674
rect 578620 480 578648 16546
rect 581104 6914 581132 177239
rect 581012 6886 581132 6914
rect 581012 480 581040 6886
rect 583392 3800 583444 3806
rect 583392 3742 583444 3748
rect 582196 3596 582248 3602
rect 582196 3538 582248 3544
rect 582208 480 582236 3538
rect 583404 480 583432 3742
rect 576278 354 576390 480
rect 575860 326 576390 354
rect 576278 -960 576390 326
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 2778 684256 2834 684312
rect 3422 671200 3478 671256
rect 2778 632068 2780 632088
rect 2780 632068 2832 632088
rect 2832 632068 2834 632088
rect 2778 632032 2834 632068
rect 3330 606056 3386 606112
rect 2778 579964 2834 580000
rect 2778 579944 2780 579964
rect 2780 579944 2832 579964
rect 2832 579944 2834 579964
rect 3054 566888 3110 566944
rect 2778 553832 2834 553888
rect 3330 527856 3386 527912
rect 3330 475632 3386 475688
rect 3514 658144 3570 658200
rect 3514 619112 3570 619168
rect 3422 462576 3478 462632
rect 3606 514800 3662 514856
rect 3698 501744 3754 501800
rect 2870 449520 2926 449576
rect 217874 516840 217930 516896
rect 217598 515888 217654 515944
rect 217506 513712 217562 513768
rect 217414 488280 217470 488336
rect 217690 489912 217746 489968
rect 217782 488008 217838 488064
rect 3330 423580 3332 423600
rect 3332 423580 3384 423600
rect 3384 423580 3386 423600
rect 3330 423544 3386 423580
rect 3330 410488 3386 410544
rect 3330 371320 3386 371376
rect 3330 358400 3386 358456
rect 3330 319232 3386 319288
rect 3238 267144 3294 267200
rect 2778 254088 2834 254144
rect 3330 214920 3386 214976
rect 3974 397432 4030 397488
rect 3882 345344 3938 345400
rect 3790 306176 3846 306232
rect 3698 293120 3754 293176
rect 3606 241032 3662 241088
rect 3698 201864 3754 201920
rect 3514 188808 3570 188864
rect 3514 149776 3570 149832
rect 3514 136720 3570 136776
rect 3422 97552 3478 97608
rect 35162 308352 35218 308408
rect 75182 308488 75238 308544
rect 200302 3304 200358 3360
rect 219070 512760 219126 512816
rect 219162 510992 219218 511048
rect 219346 509904 219402 509960
rect 219254 508136 219310 508192
rect 264978 477264 265034 477320
rect 268014 477264 268070 477320
rect 255318 477128 255374 477184
rect 252558 476720 252614 476776
rect 210882 155488 210938 155544
rect 212078 303048 212134 303104
rect 211066 155760 211122 155816
rect 210974 155352 211030 155408
rect 211986 302776 212042 302832
rect 212354 155624 212410 155680
rect 213274 302912 213330 302968
rect 213182 155216 213238 155272
rect 213550 155896 213606 155952
rect 214930 300056 214986 300112
rect 213366 3440 213422 3496
rect 214470 3440 214526 3496
rect 215666 3440 215722 3496
rect 215114 3168 215170 3224
rect 217046 193704 217102 193760
rect 216678 192752 216734 192808
rect 216678 188128 216734 188184
rect 217138 169904 217194 169960
rect 217414 196832 217470 196888
rect 217506 195880 217562 195936
rect 217598 168272 217654 168328
rect 217690 168000 217746 168056
rect 218426 243344 218482 243400
rect 218610 190984 218666 191040
rect 218518 189896 218574 189952
rect 218886 158480 218942 158536
rect 218058 3576 218114 3632
rect 235906 476176 235962 476232
rect 237378 476312 237434 476368
rect 237470 476176 237526 476232
rect 240138 476176 240194 476232
rect 241426 476176 241482 476232
rect 244278 476584 244334 476640
rect 247038 476584 247094 476640
rect 249798 476584 249854 476640
rect 242898 476332 242954 476368
rect 242898 476312 242900 476332
rect 242900 476312 242952 476332
rect 242952 476312 242954 476332
rect 244278 476312 244334 476368
rect 242806 476196 242862 476232
rect 242806 476176 242808 476196
rect 242808 476176 242860 476196
rect 242860 476176 242862 476196
rect 245658 476176 245714 476232
rect 247222 476176 247278 476232
rect 249798 476176 249854 476232
rect 251086 476176 251142 476232
rect 252374 476312 252430 476368
rect 252466 476176 252522 476232
rect 259366 476856 259422 476912
rect 253846 476176 253902 476232
rect 255226 476176 255282 476232
rect 258262 476584 258318 476640
rect 256606 476176 256662 476232
rect 257986 476176 258042 476232
rect 263598 476584 263654 476640
rect 260838 476468 260894 476504
rect 260838 476448 260840 476468
rect 260840 476448 260892 476468
rect 260892 476448 260894 476468
rect 261482 476312 261538 476368
rect 263506 476312 263562 476368
rect 260746 476176 260802 476232
rect 262862 476176 262918 476232
rect 264886 476176 264942 476232
rect 280158 476992 280214 477048
rect 304998 476992 305054 477048
rect 307758 476992 307814 477048
rect 277858 476856 277914 476912
rect 270498 476720 270554 476776
rect 273258 476448 273314 476504
rect 267554 476312 267610 476368
rect 274546 476312 274602 476368
rect 276018 476312 276074 476368
rect 278042 476720 278098 476776
rect 266266 476176 266322 476232
rect 267646 476176 267702 476232
rect 269026 476176 269082 476232
rect 270406 476176 270462 476232
rect 271786 476176 271842 476232
rect 273166 476176 273222 476232
rect 275282 476176 275338 476232
rect 276662 476176 276718 476232
rect 302238 476740 302294 476776
rect 302238 476720 302240 476740
rect 302240 476720 302292 476740
rect 302292 476720 302294 476740
rect 278686 476176 278742 476232
rect 280066 476176 280122 476232
rect 310518 476856 310574 476912
rect 282918 476196 282974 476232
rect 282918 476176 282920 476196
rect 282920 476176 282972 476196
rect 282972 476176 282974 476196
rect 285770 476176 285826 476232
rect 287150 476176 287206 476232
rect 289910 476176 289966 476232
rect 292670 476176 292726 476232
rect 295338 476176 295394 476232
rect 298098 476176 298154 476232
rect 300858 476176 300914 476232
rect 322938 476720 322994 476776
rect 313278 476468 313334 476504
rect 313278 476448 313280 476468
rect 313280 476448 313332 476468
rect 313332 476448 313334 476468
rect 314658 476448 314714 476504
rect 317418 476332 317474 476368
rect 317418 476312 317420 476332
rect 317420 476312 317472 476332
rect 317472 476312 317474 476332
rect 320178 476312 320234 476368
rect 325790 476176 325846 476232
rect 296534 446120 296590 446176
rect 294970 445984 295026 446040
rect 295706 445848 295762 445904
rect 300398 444488 300454 444544
rect 350998 444352 351054 444408
rect 580170 697176 580226 697232
rect 580262 683848 580318 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579618 590960 579674 591016
rect 580170 564304 580226 564360
rect 580170 537784 580226 537840
rect 580170 484608 580226 484664
rect 580354 644000 580410 644056
rect 580446 577632 580502 577688
rect 362222 443400 362278 443456
rect 362774 443400 362830 443456
rect 363050 443400 363106 443456
rect 558182 446120 558238 446176
rect 554042 445848 554098 445904
rect 233422 308488 233478 308544
rect 234526 308352 234582 308408
rect 270498 262792 270554 262848
rect 274638 306992 274694 307048
rect 274914 306176 274970 306232
rect 275558 308896 275614 308952
rect 275374 306040 275430 306096
rect 275834 305904 275890 305960
rect 276018 305768 276074 305824
rect 276938 308760 276994 308816
rect 276754 303320 276810 303376
rect 278318 308624 278374 308680
rect 278134 303184 278190 303240
rect 277398 303048 277454 303104
rect 279514 302912 279570 302968
rect 278778 302776 278834 302832
rect 273718 275168 273774 275224
rect 273534 265512 273590 265568
rect 273350 249056 273406 249112
rect 281354 305632 281410 305688
rect 283194 300056 283250 300112
rect 274638 246200 274694 246256
rect 295522 248104 295578 248160
rect 296718 245112 296774 245168
rect 295430 244976 295486 245032
rect 298466 308488 298522 308544
rect 299110 308352 299166 308408
rect 299478 245384 299534 245440
rect 301134 250688 301190 250744
rect 302698 284824 302754 284880
rect 302606 267008 302662 267064
rect 302514 260072 302570 260128
rect 304078 298696 304134 298752
rect 303894 286320 303950 286376
rect 303802 269728 303858 269784
rect 303618 254496 303674 254552
rect 309782 304272 309838 304328
rect 309966 304136 310022 304192
rect 302330 249056 302386 249112
rect 311162 306040 311218 306096
rect 311346 305904 311402 305960
rect 312726 306992 312782 307048
rect 312542 305768 312598 305824
rect 315486 302776 315542 302832
rect 316314 305632 316370 305688
rect 317602 250552 317658 250608
rect 322938 247968 322994 248024
rect 323122 247832 323178 247888
rect 324502 247696 324558 247752
rect 324318 247560 324374 247616
rect 302238 245520 302294 245576
rect 300858 245248 300914 245304
rect 329930 262792 329986 262848
rect 338210 250416 338266 250472
rect 346122 309032 346178 309088
rect 346398 308896 346454 308952
rect 347042 308760 347098 308816
rect 347318 308624 347374 308680
rect 349158 306176 349214 306232
rect 353758 308216 353814 308272
rect 296902 244840 296958 244896
rect 356610 245248 356666 245304
rect 356610 244568 356666 244624
rect 273350 159840 273406 159896
rect 278134 159840 278190 159896
rect 261114 159704 261170 159760
rect 220818 158616 220874 158672
rect 238114 158652 238116 158672
rect 238116 158652 238168 158672
rect 238168 158652 238170 158672
rect 219438 158344 219494 158400
rect 238114 158616 238170 158652
rect 239586 158616 239642 158672
rect 242438 158616 242494 158672
rect 244646 158616 244702 158672
rect 245566 158616 245622 158672
rect 248326 158616 248382 158672
rect 252374 158616 252430 158672
rect 255870 158616 255926 158672
rect 224958 158480 225014 158536
rect 223578 157936 223634 157992
rect 216862 3440 216918 3496
rect 216586 3032 216642 3088
rect 219346 3576 219402 3632
rect 219254 3440 219310 3496
rect 219346 3032 219402 3088
rect 222750 3848 222806 3904
rect 227718 158208 227774 158264
rect 227534 3712 227590 3768
rect 226338 3168 226394 3224
rect 234618 158072 234674 158128
rect 234710 157936 234766 157992
rect 241426 158208 241482 158264
rect 246670 157936 246726 157992
rect 247958 157936 248014 157992
rect 237010 3440 237066 3496
rect 248694 157800 248750 157856
rect 251086 157936 251142 157992
rect 250442 157800 250498 157856
rect 252466 157800 252522 157856
rect 253478 157800 253534 157856
rect 256238 157528 256294 157584
rect 253938 155896 253994 155952
rect 255318 155760 255374 155816
rect 251178 3168 251234 3224
rect 257250 158616 257306 158672
rect 259550 155624 259606 155680
rect 261758 158616 261814 158672
rect 263690 157528 263746 157584
rect 275834 159568 275890 159624
rect 277030 159568 277086 159624
rect 355322 159704 355378 159760
rect 279238 159568 279294 159624
rect 265438 158616 265494 158672
rect 265990 158616 266046 158672
rect 266542 158616 266598 158672
rect 268750 158616 268806 158672
rect 269946 158652 269948 158672
rect 269948 158652 270000 158672
rect 270000 158652 270002 158672
rect 269946 158616 270002 158652
rect 270958 158616 271014 158672
rect 272246 158616 272302 158672
rect 274454 158616 274510 158672
rect 276110 158616 276166 158672
rect 281078 158616 281134 158672
rect 268382 157664 268438 157720
rect 267830 155488 267886 155544
rect 271326 157664 271382 157720
rect 273718 157664 273774 157720
rect 269118 155352 269174 155408
rect 278502 157664 278558 157720
rect 274638 155216 274694 155272
rect 283654 157528 283710 157584
rect 288254 158616 288310 158672
rect 291014 158616 291070 158672
rect 293590 158616 293646 158672
rect 295982 158652 295984 158672
rect 295984 158652 296036 158672
rect 296036 158652 296038 158672
rect 295982 158616 296038 158652
rect 298558 158616 298614 158672
rect 300950 158616 301006 158672
rect 303526 158616 303582 158672
rect 306102 158616 306158 158672
rect 308678 158616 308734 158672
rect 286046 157528 286102 157584
rect 311070 158616 311126 158672
rect 313462 158616 313518 158672
rect 315854 158636 315910 158672
rect 315854 158616 315856 158636
rect 315856 158616 315908 158636
rect 315908 158616 315910 158636
rect 318614 158616 318670 158672
rect 321006 158616 321062 158672
rect 323398 158616 323454 158672
rect 325974 158616 326030 158672
rect 355322 157800 355378 157856
rect 322110 8880 322166 8936
rect 320914 6160 320970 6216
rect 325606 3440 325662 3496
rect 324410 3304 324466 3360
rect 331586 3576 331642 3632
rect 351642 6704 351698 6760
rect 348054 6568 348110 6624
rect 346950 6432 347006 6488
rect 344558 6296 344614 6352
rect 335082 3712 335138 3768
rect 338670 3848 338726 3904
rect 342166 3984 342222 4040
rect 345754 3168 345810 3224
rect 356886 244704 356942 244760
rect 357438 245112 357494 245168
rect 357438 159296 357494 159352
rect 357714 159704 357770 159760
rect 359002 307944 359058 308000
rect 361486 307808 361542 307864
rect 361118 159296 361174 159352
rect 358726 3440 358782 3496
rect 359922 3440 359978 3496
rect 361118 3440 361174 3496
rect 361670 6704 361726 6760
rect 365166 309032 365222 309088
rect 363510 3440 363566 3496
rect 363878 159296 363934 159352
rect 364706 6568 364762 6624
rect 365166 158480 365222 158536
rect 364798 6432 364854 6488
rect 366454 159432 366510 159488
rect 366546 158208 366602 158264
rect 366178 6296 366234 6352
rect 367466 308760 367522 308816
rect 367558 158344 367614 158400
rect 367466 157392 367522 157448
rect 367834 308896 367890 308952
rect 368018 308216 368074 308272
rect 367926 159160 367982 159216
rect 368018 159024 368074 159080
rect 367834 158752 367890 158808
rect 370042 308624 370098 308680
rect 369122 158072 369178 158128
rect 370226 306176 370282 306232
rect 467838 307944 467894 308000
rect 370502 157936 370558 157992
rect 370686 158888 370742 158944
rect 368662 8880 368718 8936
rect 364614 3440 364670 3496
rect 365810 3440 365866 3496
rect 368202 3440 368258 3496
rect 369398 3440 369454 3496
rect 370594 3440 370650 3496
rect 400218 306040 400274 306096
rect 392582 302776 392638 302832
rect 394238 3712 394294 3768
rect 397734 3576 397790 3632
rect 404358 305904 404414 305960
rect 407118 305768 407174 305824
rect 411902 3440 411958 3496
rect 429198 305632 429254 305688
rect 438858 250552 438914 250608
rect 465170 247968 465226 248024
rect 471978 307808 472034 307864
rect 469218 247832 469274 247888
rect 473450 247696 473506 247752
rect 476118 247560 476174 247616
rect 501786 3304 501842 3360
rect 546498 250416 546554 250472
rect 580170 431568 580226 431624
rect 579618 378392 579674 378448
rect 579986 325216 580042 325272
rect 580170 272176 580226 272232
rect 580630 232328 580686 232384
rect 580538 192480 580594 192536
rect 581090 177248 581146 177304
rect 580446 152632 580502 152688
rect 580354 112784 580410 112840
rect 580262 33088 580318 33144
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 2773 684314 2839 684317
rect -960 684312 2839 684314
rect -960 684256 2778 684312
rect 2834 684256 2839 684312
rect -960 684254 2839 684256
rect -960 684164 480 684254
rect 2773 684251 2839 684254
rect 580257 683906 580323 683909
rect 583520 683906 584960 683996
rect 580257 683904 584960 683906
rect 580257 683848 580262 683904
rect 580318 683848 584960 683904
rect 580257 683846 584960 683848
rect 580257 683843 580323 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580349 644058 580415 644061
rect 583520 644058 584960 644148
rect 580349 644056 584960 644058
rect 580349 644000 580354 644056
rect 580410 644000 584960 644056
rect 580349 643998 584960 644000
rect 580349 643995 580415 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 2773 632090 2839 632093
rect -960 632088 2839 632090
rect -960 632032 2778 632088
rect 2834 632032 2839 632088
rect -960 632030 2839 632032
rect -960 631940 480 632030
rect 2773 632027 2839 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3325 606114 3391 606117
rect -960 606112 3391 606114
rect -960 606056 3330 606112
rect 3386 606056 3391 606112
rect -960 606054 3391 606056
rect -960 605964 480 606054
rect 3325 606051 3391 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579613 591018 579679 591021
rect 583520 591018 584960 591108
rect 579613 591016 584960 591018
rect 579613 590960 579618 591016
rect 579674 590960 584960 591016
rect 579613 590958 584960 590960
rect 579613 590955 579679 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 2773 580002 2839 580005
rect -960 580000 2839 580002
rect -960 579944 2778 580000
rect 2834 579944 2839 580000
rect -960 579942 2839 579944
rect -960 579852 480 579942
rect 2773 579939 2839 579942
rect 580441 577690 580507 577693
rect 583520 577690 584960 577780
rect 580441 577688 584960 577690
rect 580441 577632 580446 577688
rect 580502 577632 584960 577688
rect 580441 577630 584960 577632
rect 580441 577627 580507 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3049 566946 3115 566949
rect -960 566944 3115 566946
rect -960 566888 3054 566944
rect 3110 566888 3115 566944
rect -960 566886 3115 566888
rect -960 566796 480 566886
rect 3049 566883 3115 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 2773 553890 2839 553893
rect -960 553888 2839 553890
rect -960 553832 2778 553888
rect 2834 553832 2839 553888
rect -960 553830 2839 553832
rect -960 553740 480 553830
rect 2773 553827 2839 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3325 527914 3391 527917
rect -960 527912 3391 527914
rect -960 527856 3330 527912
rect 3386 527856 3391 527912
rect -960 527854 3391 527856
rect -960 527764 480 527854
rect 3325 527851 3391 527854
rect 583520 524364 584960 524604
rect 217869 516898 217935 516901
rect 219390 516898 220064 516924
rect 217869 516896 220064 516898
rect 217869 516840 217874 516896
rect 217930 516864 220064 516896
rect 217930 516840 219450 516864
rect 217869 516838 219450 516840
rect 217869 516835 217935 516838
rect 217593 515946 217659 515949
rect 219390 515946 220064 515972
rect 217593 515944 220064 515946
rect 217593 515888 217598 515944
rect 217654 515912 220064 515944
rect 217654 515888 219450 515912
rect 217593 515886 219450 515888
rect 217593 515883 217659 515886
rect -960 514858 480 514948
rect 3601 514858 3667 514861
rect -960 514856 3667 514858
rect -960 514800 3606 514856
rect 3662 514800 3667 514856
rect -960 514798 3667 514800
rect -960 514708 480 514798
rect 3601 514795 3667 514798
rect 217501 513770 217567 513773
rect 219390 513770 220064 513796
rect 217501 513768 220064 513770
rect 217501 513712 217506 513768
rect 217562 513736 220064 513768
rect 217562 513712 219450 513736
rect 217501 513710 219450 513712
rect 217501 513707 217567 513710
rect 219065 512818 219131 512821
rect 219390 512818 220064 512844
rect 219065 512816 220064 512818
rect 219065 512760 219070 512816
rect 219126 512784 220064 512816
rect 219126 512760 219450 512784
rect 219065 512758 219450 512760
rect 219065 512755 219131 512758
rect 583520 511172 584960 511412
rect 219157 511050 219223 511053
rect 219390 511050 220064 511076
rect 219157 511048 220064 511050
rect 219157 510992 219162 511048
rect 219218 511016 220064 511048
rect 219218 510992 219450 511016
rect 219157 510990 219450 510992
rect 219157 510987 219223 510990
rect 219390 509965 220064 509988
rect 219341 509960 220064 509965
rect 219341 509904 219346 509960
rect 219402 509928 220064 509960
rect 219402 509904 219450 509928
rect 219341 509902 219450 509904
rect 219341 509899 219407 509902
rect 219249 508194 219315 508197
rect 219390 508194 220064 508220
rect 219249 508192 220064 508194
rect 219249 508136 219254 508192
rect 219310 508160 220064 508192
rect 219310 508136 219450 508160
rect 219249 508134 219450 508136
rect 219249 508131 219315 508134
rect -960 501802 480 501892
rect 3693 501802 3759 501805
rect -960 501800 3759 501802
rect -960 501744 3698 501800
rect 3754 501744 3759 501800
rect -960 501742 3759 501744
rect -960 501652 480 501742
rect 3693 501739 3759 501742
rect 583520 497844 584960 498084
rect 217685 489970 217751 489973
rect 219390 489970 220064 489996
rect 217685 489968 220064 489970
rect 217685 489912 217690 489968
rect 217746 489936 220064 489968
rect 217746 489912 219450 489936
rect 217685 489910 219450 489912
rect 217685 489907 217751 489910
rect -960 488596 480 488836
rect 217409 488338 217475 488341
rect 219390 488338 220064 488364
rect 217409 488336 220064 488338
rect 217409 488280 217414 488336
rect 217470 488304 220064 488336
rect 217470 488280 219450 488304
rect 217409 488278 219450 488280
rect 217409 488275 217475 488278
rect 217777 488066 217843 488069
rect 219390 488066 220064 488092
rect 217777 488064 220064 488066
rect 217777 488008 217782 488064
rect 217838 488032 220064 488064
rect 217838 488008 219450 488032
rect 217777 488006 219450 488008
rect 217777 488003 217843 488006
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect 264973 477322 265039 477325
rect 265934 477322 265940 477324
rect 264973 477320 265940 477322
rect 264973 477264 264978 477320
rect 265034 477264 265940 477320
rect 264973 477262 265940 477264
rect 264973 477259 265039 477262
rect 265934 477260 265940 477262
rect 266004 477260 266010 477324
rect 268009 477322 268075 477325
rect 268326 477322 268332 477324
rect 268009 477320 268332 477322
rect 268009 477264 268014 477320
rect 268070 477264 268332 477320
rect 268009 477262 268332 477264
rect 268009 477259 268075 477262
rect 268326 477260 268332 477262
rect 268396 477260 268402 477324
rect 255313 477186 255379 477189
rect 256182 477186 256188 477188
rect 255313 477184 256188 477186
rect 255313 477128 255318 477184
rect 255374 477128 256188 477184
rect 255313 477126 256188 477128
rect 255313 477123 255379 477126
rect 256182 477124 256188 477126
rect 256252 477124 256258 477188
rect 280153 477050 280219 477053
rect 280838 477050 280844 477052
rect 280153 477048 280844 477050
rect 280153 476992 280158 477048
rect 280214 476992 280844 477048
rect 280153 476990 280844 476992
rect 280153 476987 280219 476990
rect 280838 476988 280844 476990
rect 280908 476988 280914 477052
rect 304993 477050 305059 477053
rect 305862 477050 305868 477052
rect 304993 477048 305868 477050
rect 304993 476992 304998 477048
rect 305054 476992 305868 477048
rect 304993 476990 305868 476992
rect 304993 476987 305059 476990
rect 305862 476988 305868 476990
rect 305932 476988 305938 477052
rect 307753 477050 307819 477053
rect 308438 477050 308444 477052
rect 307753 477048 308444 477050
rect 307753 476992 307758 477048
rect 307814 476992 308444 477048
rect 307753 476990 308444 476992
rect 307753 476987 307819 476990
rect 308438 476988 308444 476990
rect 308508 476988 308514 477052
rect 258022 476852 258028 476916
rect 258092 476914 258098 476916
rect 259361 476914 259427 476917
rect 258092 476912 259427 476914
rect 258092 476856 259366 476912
rect 259422 476856 259427 476912
rect 258092 476854 259427 476856
rect 258092 476852 258098 476854
rect 259361 476851 259427 476854
rect 277853 476914 277919 476917
rect 278446 476914 278452 476916
rect 277853 476912 278452 476914
rect 277853 476856 277858 476912
rect 277914 476856 278452 476912
rect 277853 476854 278452 476856
rect 277853 476851 277919 476854
rect 278446 476852 278452 476854
rect 278516 476852 278522 476916
rect 310513 476914 310579 476917
rect 311014 476914 311020 476916
rect 310513 476912 311020 476914
rect 310513 476856 310518 476912
rect 310574 476856 311020 476912
rect 310513 476854 311020 476856
rect 310513 476851 310579 476854
rect 311014 476852 311020 476854
rect 311084 476852 311090 476916
rect 252553 476778 252619 476781
rect 253606 476778 253612 476780
rect 252553 476776 253612 476778
rect 252553 476720 252558 476776
rect 252614 476720 253612 476776
rect 252553 476718 253612 476720
rect 252553 476715 252619 476718
rect 253606 476716 253612 476718
rect 253676 476716 253682 476780
rect 270493 476778 270559 476781
rect 270902 476778 270908 476780
rect 270493 476776 270908 476778
rect 270493 476720 270498 476776
rect 270554 476720 270908 476776
rect 270493 476718 270908 476720
rect 270493 476715 270559 476718
rect 270902 476716 270908 476718
rect 270972 476716 270978 476780
rect 276974 476716 276980 476780
rect 277044 476778 277050 476780
rect 278037 476778 278103 476781
rect 277044 476776 278103 476778
rect 277044 476720 278042 476776
rect 278098 476720 278103 476776
rect 277044 476718 278103 476720
rect 277044 476716 277050 476718
rect 278037 476715 278103 476718
rect 302233 476778 302299 476781
rect 303470 476778 303476 476780
rect 302233 476776 303476 476778
rect 302233 476720 302238 476776
rect 302294 476720 303476 476776
rect 302233 476718 303476 476720
rect 302233 476715 302299 476718
rect 303470 476716 303476 476718
rect 303540 476716 303546 476780
rect 322933 476778 322999 476781
rect 323342 476778 323348 476780
rect 322933 476776 323348 476778
rect 322933 476720 322938 476776
rect 322994 476720 323348 476776
rect 322933 476718 323348 476720
rect 322933 476715 322999 476718
rect 323342 476716 323348 476718
rect 323412 476716 323418 476780
rect 244273 476644 244339 476645
rect 244222 476580 244228 476644
rect 244292 476642 244339 476644
rect 247033 476642 247099 476645
rect 248270 476642 248276 476644
rect 244292 476640 244384 476642
rect 244334 476584 244384 476640
rect 244292 476582 244384 476584
rect 247033 476640 248276 476642
rect 247033 476584 247038 476640
rect 247094 476584 248276 476640
rect 247033 476582 248276 476584
rect 244292 476580 244339 476582
rect 244273 476579 244339 476580
rect 247033 476579 247099 476582
rect 248270 476580 248276 476582
rect 248340 476580 248346 476644
rect 249793 476642 249859 476645
rect 250662 476642 250668 476644
rect 249793 476640 250668 476642
rect 249793 476584 249798 476640
rect 249854 476584 250668 476640
rect 249793 476582 250668 476584
rect 249793 476579 249859 476582
rect 250662 476580 250668 476582
rect 250732 476580 250738 476644
rect 258257 476642 258323 476645
rect 263593 476644 263659 476645
rect 258390 476642 258396 476644
rect 258257 476640 258396 476642
rect 258257 476584 258262 476640
rect 258318 476584 258396 476640
rect 258257 476582 258396 476584
rect 258257 476579 258323 476582
rect 258390 476580 258396 476582
rect 258460 476580 258466 476644
rect 263542 476580 263548 476644
rect 263612 476642 263659 476644
rect 263612 476640 263704 476642
rect 263654 476584 263704 476640
rect 263612 476582 263704 476584
rect 263612 476580 263659 476582
rect 263593 476579 263659 476580
rect 260833 476506 260899 476509
rect 260966 476506 260972 476508
rect 260833 476504 260972 476506
rect 260833 476448 260838 476504
rect 260894 476448 260972 476504
rect 260833 476446 260972 476448
rect 260833 476443 260899 476446
rect 260966 476444 260972 476446
rect 261036 476444 261042 476508
rect 273253 476506 273319 476509
rect 273478 476506 273484 476508
rect 273253 476504 273484 476506
rect 273253 476448 273258 476504
rect 273314 476448 273484 476504
rect 273253 476446 273484 476448
rect 273253 476443 273319 476446
rect 273478 476444 273484 476446
rect 273548 476444 273554 476508
rect 313273 476506 313339 476509
rect 313406 476506 313412 476508
rect 313273 476504 313412 476506
rect 313273 476448 313278 476504
rect 313334 476448 313412 476504
rect 313273 476446 313412 476448
rect 313273 476443 313339 476446
rect 313406 476444 313412 476446
rect 313476 476444 313482 476508
rect 314653 476506 314719 476509
rect 315798 476506 315804 476508
rect 314653 476504 315804 476506
rect 314653 476448 314658 476504
rect 314714 476448 315804 476504
rect 314653 476446 315804 476448
rect 314653 476443 314719 476446
rect 315798 476444 315804 476446
rect 315868 476444 315874 476508
rect 237373 476370 237439 476373
rect 238150 476370 238156 476372
rect 237373 476368 238156 476370
rect 237373 476312 237378 476368
rect 237434 476312 238156 476368
rect 237373 476310 238156 476312
rect 237373 476307 237439 476310
rect 238150 476308 238156 476310
rect 238220 476308 238226 476372
rect 242893 476370 242959 476373
rect 243118 476370 243124 476372
rect 242893 476368 243124 476370
rect 242893 476312 242898 476368
rect 242954 476312 243124 476368
rect 242893 476310 243124 476312
rect 242893 476307 242959 476310
rect 243118 476308 243124 476310
rect 243188 476308 243194 476372
rect 244273 476370 244339 476373
rect 252369 476372 252435 476373
rect 245326 476370 245332 476372
rect 244273 476368 245332 476370
rect 244273 476312 244278 476368
rect 244334 476312 245332 476368
rect 244273 476310 245332 476312
rect 244273 476307 244339 476310
rect 245326 476308 245332 476310
rect 245396 476308 245402 476372
rect 252318 476308 252324 476372
rect 252388 476370 252435 476372
rect 252388 476368 252480 476370
rect 252430 476312 252480 476368
rect 252388 476310 252480 476312
rect 252388 476308 252435 476310
rect 260782 476308 260788 476372
rect 260852 476370 260858 476372
rect 261477 476370 261543 476373
rect 260852 476368 261543 476370
rect 260852 476312 261482 476368
rect 261538 476312 261543 476368
rect 260852 476310 261543 476312
rect 260852 476308 260858 476310
rect 252369 476307 252435 476308
rect 261477 476307 261543 476310
rect 262806 476308 262812 476372
rect 262876 476370 262882 476372
rect 263501 476370 263567 476373
rect 262876 476368 263567 476370
rect 262876 476312 263506 476368
rect 263562 476312 263567 476368
rect 262876 476310 263567 476312
rect 262876 476308 262882 476310
rect 263501 476307 263567 476310
rect 266486 476308 266492 476372
rect 266556 476370 266562 476372
rect 267549 476370 267615 476373
rect 266556 476368 267615 476370
rect 266556 476312 267554 476368
rect 267610 476312 267615 476368
rect 266556 476310 267615 476312
rect 266556 476308 266562 476310
rect 267549 476307 267615 476310
rect 273294 476308 273300 476372
rect 273364 476370 273370 476372
rect 274541 476370 274607 476373
rect 276013 476372 276079 476373
rect 276013 476370 276060 476372
rect 273364 476368 274607 476370
rect 273364 476312 274546 476368
rect 274602 476312 274607 476368
rect 273364 476310 274607 476312
rect 275968 476368 276060 476370
rect 275968 476312 276018 476368
rect 275968 476310 276060 476312
rect 273364 476308 273370 476310
rect 274541 476307 274607 476310
rect 276013 476308 276060 476310
rect 276124 476308 276130 476372
rect 317413 476370 317479 476373
rect 318374 476370 318380 476372
rect 317413 476368 318380 476370
rect 317413 476312 317418 476368
rect 317474 476312 318380 476368
rect 317413 476310 318380 476312
rect 276013 476307 276079 476308
rect 317413 476307 317479 476310
rect 318374 476308 318380 476310
rect 318444 476308 318450 476372
rect 320173 476370 320239 476373
rect 320950 476370 320956 476372
rect 320173 476368 320956 476370
rect 320173 476312 320178 476368
rect 320234 476312 320956 476368
rect 320173 476310 320956 476312
rect 320173 476307 320239 476310
rect 320950 476308 320956 476310
rect 321020 476308 321026 476372
rect 235901 476236 235967 476237
rect 235901 476234 235948 476236
rect 235856 476232 235948 476234
rect 235856 476176 235906 476232
rect 235856 476174 235948 476176
rect 235901 476172 235948 476174
rect 236012 476172 236018 476236
rect 237230 476172 237236 476236
rect 237300 476234 237306 476236
rect 237465 476234 237531 476237
rect 237300 476232 237531 476234
rect 237300 476176 237470 476232
rect 237526 476176 237531 476232
rect 237300 476174 237531 476176
rect 237300 476172 237306 476174
rect 235901 476171 235967 476172
rect 237465 476171 237531 476174
rect 239622 476172 239628 476236
rect 239692 476234 239698 476236
rect 240133 476234 240199 476237
rect 239692 476232 240199 476234
rect 239692 476176 240138 476232
rect 240194 476176 240199 476232
rect 239692 476174 240199 476176
rect 239692 476172 239698 476174
rect 240133 476171 240199 476174
rect 240542 476172 240548 476236
rect 240612 476234 240618 476236
rect 241421 476234 241487 476237
rect 240612 476232 241487 476234
rect 240612 476176 241426 476232
rect 241482 476176 241487 476232
rect 240612 476174 241487 476176
rect 240612 476172 240618 476174
rect 241421 476171 241487 476174
rect 241830 476172 241836 476236
rect 241900 476234 241906 476236
rect 242801 476234 242867 476237
rect 241900 476232 242867 476234
rect 241900 476176 242806 476232
rect 242862 476176 242867 476232
rect 241900 476174 242867 476176
rect 241900 476172 241906 476174
rect 242801 476171 242867 476174
rect 245653 476234 245719 476237
rect 246430 476234 246436 476236
rect 245653 476232 246436 476234
rect 245653 476176 245658 476232
rect 245714 476176 246436 476232
rect 245653 476174 246436 476176
rect 245653 476171 245719 476174
rect 246430 476172 246436 476174
rect 246500 476172 246506 476236
rect 247217 476234 247283 476237
rect 247534 476234 247540 476236
rect 247217 476232 247540 476234
rect 247217 476176 247222 476232
rect 247278 476176 247540 476232
rect 247217 476174 247540 476176
rect 247217 476171 247283 476174
rect 247534 476172 247540 476174
rect 247604 476172 247610 476236
rect 248638 476172 248644 476236
rect 248708 476234 248714 476236
rect 249793 476234 249859 476237
rect 248708 476232 249859 476234
rect 248708 476176 249798 476232
rect 249854 476176 249859 476232
rect 248708 476174 249859 476176
rect 248708 476172 248714 476174
rect 249793 476171 249859 476174
rect 250110 476172 250116 476236
rect 250180 476234 250186 476236
rect 251081 476234 251147 476237
rect 250180 476232 251147 476234
rect 250180 476176 251086 476232
rect 251142 476176 251147 476232
rect 250180 476174 251147 476176
rect 250180 476172 250186 476174
rect 251081 476171 251147 476174
rect 251398 476172 251404 476236
rect 251468 476234 251474 476236
rect 252461 476234 252527 476237
rect 251468 476232 252527 476234
rect 251468 476176 252466 476232
rect 252522 476176 252527 476232
rect 251468 476174 252527 476176
rect 251468 476172 251474 476174
rect 252461 476171 252527 476174
rect 253422 476172 253428 476236
rect 253492 476234 253498 476236
rect 253841 476234 253907 476237
rect 253492 476232 253907 476234
rect 253492 476176 253846 476232
rect 253902 476176 253907 476232
rect 253492 476174 253907 476176
rect 253492 476172 253498 476174
rect 253841 476171 253907 476174
rect 254526 476172 254532 476236
rect 254596 476234 254602 476236
rect 255221 476234 255287 476237
rect 254596 476232 255287 476234
rect 254596 476176 255226 476232
rect 255282 476176 255287 476232
rect 254596 476174 255287 476176
rect 254596 476172 254602 476174
rect 255221 476171 255287 476174
rect 255814 476172 255820 476236
rect 255884 476234 255890 476236
rect 256601 476234 256667 476237
rect 255884 476232 256667 476234
rect 255884 476176 256606 476232
rect 256662 476176 256667 476232
rect 255884 476174 256667 476176
rect 255884 476172 255890 476174
rect 256601 476171 256667 476174
rect 257102 476172 257108 476236
rect 257172 476234 257178 476236
rect 257981 476234 258047 476237
rect 257172 476232 258047 476234
rect 257172 476176 257986 476232
rect 258042 476176 258047 476232
rect 257172 476174 258047 476176
rect 257172 476172 257178 476174
rect 257981 476171 258047 476174
rect 259494 476172 259500 476236
rect 259564 476234 259570 476236
rect 260741 476234 260807 476237
rect 259564 476232 260807 476234
rect 259564 476176 260746 476232
rect 260802 476176 260807 476232
rect 259564 476174 260807 476176
rect 259564 476172 259570 476174
rect 260741 476171 260807 476174
rect 261702 476172 261708 476236
rect 261772 476234 261778 476236
rect 262857 476234 262923 476237
rect 261772 476232 262923 476234
rect 261772 476176 262862 476232
rect 262918 476176 262923 476232
rect 261772 476174 262923 476176
rect 261772 476172 261778 476174
rect 262857 476171 262923 476174
rect 263910 476172 263916 476236
rect 263980 476234 263986 476236
rect 264881 476234 264947 476237
rect 263980 476232 264947 476234
rect 263980 476176 264886 476232
rect 264942 476176 264947 476232
rect 263980 476174 264947 476176
rect 263980 476172 263986 476174
rect 264881 476171 264947 476174
rect 265382 476172 265388 476236
rect 265452 476234 265458 476236
rect 266261 476234 266327 476237
rect 267641 476236 267707 476237
rect 267590 476234 267596 476236
rect 265452 476232 266327 476234
rect 265452 476176 266266 476232
rect 266322 476176 266327 476232
rect 265452 476174 266327 476176
rect 267550 476174 267596 476234
rect 267660 476232 267707 476236
rect 267702 476176 267707 476232
rect 265452 476172 265458 476174
rect 266261 476171 266327 476174
rect 267590 476172 267596 476174
rect 267660 476172 267707 476176
rect 268694 476172 268700 476236
rect 268764 476234 268770 476236
rect 269021 476234 269087 476237
rect 268764 476232 269087 476234
rect 268764 476176 269026 476232
rect 269082 476176 269087 476232
rect 268764 476174 269087 476176
rect 268764 476172 268770 476174
rect 267641 476171 267707 476172
rect 269021 476171 269087 476174
rect 269798 476172 269804 476236
rect 269868 476234 269874 476236
rect 270401 476234 270467 476237
rect 269868 476232 270467 476234
rect 269868 476176 270406 476232
rect 270462 476176 270467 476232
rect 269868 476174 270467 476176
rect 269868 476172 269874 476174
rect 270401 476171 270467 476174
rect 271270 476172 271276 476236
rect 271340 476234 271346 476236
rect 271781 476234 271847 476237
rect 271340 476232 271847 476234
rect 271340 476176 271786 476232
rect 271842 476176 271847 476232
rect 271340 476174 271847 476176
rect 271340 476172 271346 476174
rect 271781 476171 271847 476174
rect 272190 476172 272196 476236
rect 272260 476234 272266 476236
rect 273161 476234 273227 476237
rect 272260 476232 273227 476234
rect 272260 476176 273166 476232
rect 273222 476176 273227 476232
rect 272260 476174 273227 476176
rect 272260 476172 272266 476174
rect 273161 476171 273227 476174
rect 274398 476172 274404 476236
rect 274468 476234 274474 476236
rect 275277 476234 275343 476237
rect 274468 476232 275343 476234
rect 274468 476176 275282 476232
rect 275338 476176 275343 476232
rect 274468 476174 275343 476176
rect 274468 476172 274474 476174
rect 275277 476171 275343 476174
rect 275870 476172 275876 476236
rect 275940 476234 275946 476236
rect 276657 476234 276723 476237
rect 275940 476232 276723 476234
rect 275940 476176 276662 476232
rect 276718 476176 276723 476232
rect 275940 476174 276723 476176
rect 275940 476172 275946 476174
rect 276657 476171 276723 476174
rect 278078 476172 278084 476236
rect 278148 476234 278154 476236
rect 278681 476234 278747 476237
rect 278148 476232 278747 476234
rect 278148 476176 278686 476232
rect 278742 476176 278747 476232
rect 278148 476174 278747 476176
rect 278148 476172 278154 476174
rect 278681 476171 278747 476174
rect 279182 476172 279188 476236
rect 279252 476234 279258 476236
rect 280061 476234 280127 476237
rect 279252 476232 280127 476234
rect 279252 476176 280066 476232
rect 280122 476176 280127 476232
rect 279252 476174 280127 476176
rect 279252 476172 279258 476174
rect 280061 476171 280127 476174
rect 282913 476234 282979 476237
rect 283414 476234 283420 476236
rect 282913 476232 283420 476234
rect 282913 476176 282918 476232
rect 282974 476176 283420 476232
rect 282913 476174 283420 476176
rect 282913 476171 282979 476174
rect 283414 476172 283420 476174
rect 283484 476172 283490 476236
rect 285765 476234 285831 476237
rect 285990 476234 285996 476236
rect 285765 476232 285996 476234
rect 285765 476176 285770 476232
rect 285826 476176 285996 476232
rect 285765 476174 285996 476176
rect 285765 476171 285831 476174
rect 285990 476172 285996 476174
rect 286060 476172 286066 476236
rect 287145 476234 287211 476237
rect 288198 476234 288204 476236
rect 287145 476232 288204 476234
rect 287145 476176 287150 476232
rect 287206 476176 288204 476232
rect 287145 476174 288204 476176
rect 287145 476171 287211 476174
rect 288198 476172 288204 476174
rect 288268 476172 288274 476236
rect 289905 476234 289971 476237
rect 290958 476234 290964 476236
rect 289905 476232 290964 476234
rect 289905 476176 289910 476232
rect 289966 476176 290964 476232
rect 289905 476174 290964 476176
rect 289905 476171 289971 476174
rect 290958 476172 290964 476174
rect 291028 476172 291034 476236
rect 292665 476234 292731 476237
rect 293350 476234 293356 476236
rect 292665 476232 293356 476234
rect 292665 476176 292670 476232
rect 292726 476176 293356 476232
rect 292665 476174 293356 476176
rect 292665 476171 292731 476174
rect 293350 476172 293356 476174
rect 293420 476172 293426 476236
rect 295333 476234 295399 476237
rect 295926 476234 295932 476236
rect 295333 476232 295932 476234
rect 295333 476176 295338 476232
rect 295394 476176 295932 476232
rect 295333 476174 295932 476176
rect 295333 476171 295399 476174
rect 295926 476172 295932 476174
rect 295996 476172 296002 476236
rect 298093 476234 298159 476237
rect 300853 476236 300919 476237
rect 298502 476234 298508 476236
rect 298093 476232 298508 476234
rect 298093 476176 298098 476232
rect 298154 476176 298508 476232
rect 298093 476174 298508 476176
rect 298093 476171 298159 476174
rect 298502 476172 298508 476174
rect 298572 476172 298578 476236
rect 300853 476234 300900 476236
rect 300808 476232 300900 476234
rect 300808 476176 300858 476232
rect 300808 476174 300900 476176
rect 300853 476172 300900 476174
rect 300964 476172 300970 476236
rect 325785 476234 325851 476237
rect 325918 476234 325924 476236
rect 325785 476232 325924 476234
rect 325785 476176 325790 476232
rect 325846 476176 325924 476232
rect 325785 476174 325924 476176
rect 300853 476171 300919 476172
rect 325785 476171 325851 476174
rect 325918 476172 325924 476174
rect 325988 476172 325994 476236
rect -960 475690 480 475780
rect 3325 475690 3391 475693
rect -960 475688 3391 475690
rect -960 475632 3330 475688
rect 3386 475632 3391 475688
rect -960 475630 3391 475632
rect -960 475540 480 475630
rect 3325 475627 3391 475630
rect 583520 471324 584960 471564
rect -960 462634 480 462724
rect 3417 462634 3483 462637
rect -960 462632 3483 462634
rect -960 462576 3422 462632
rect 3478 462576 3483 462632
rect -960 462574 3483 462576
rect -960 462484 480 462574
rect 3417 462571 3483 462574
rect 583520 457996 584960 458236
rect -960 449578 480 449668
rect 2865 449578 2931 449581
rect -960 449576 2931 449578
rect -960 449520 2870 449576
rect 2926 449520 2931 449576
rect -960 449518 2931 449520
rect -960 449428 480 449518
rect 2865 449515 2931 449518
rect 296529 446178 296595 446181
rect 558177 446178 558243 446181
rect 296529 446176 558243 446178
rect 296529 446120 296534 446176
rect 296590 446120 558182 446176
rect 558238 446120 558243 446176
rect 296529 446118 558243 446120
rect 296529 446115 296595 446118
rect 558177 446115 558243 446118
rect 294965 446042 295031 446045
rect 369158 446042 369164 446044
rect 294965 446040 369164 446042
rect 294965 445984 294970 446040
rect 295026 445984 369164 446040
rect 294965 445982 369164 445984
rect 294965 445979 295031 445982
rect 369158 445980 369164 445982
rect 369228 445980 369234 446044
rect 295701 445906 295767 445909
rect 554037 445906 554103 445909
rect 295701 445904 554103 445906
rect 295701 445848 295706 445904
rect 295762 445848 554042 445904
rect 554098 445848 554103 445904
rect 295701 445846 554103 445848
rect 295701 445843 295767 445846
rect 554037 445843 554103 445846
rect 364926 444682 364932 444684
rect 354630 444622 364932 444682
rect 300393 444546 300459 444549
rect 354630 444546 354690 444622
rect 364926 444620 364932 444622
rect 364996 444620 365002 444684
rect 583520 444668 584960 444908
rect 300393 444544 354690 444546
rect 300393 444488 300398 444544
rect 300454 444488 354690 444544
rect 300393 444486 354690 444488
rect 300393 444483 300459 444486
rect 214414 444348 214420 444412
rect 214484 444410 214490 444412
rect 350993 444410 351059 444413
rect 214484 444408 351059 444410
rect 214484 444352 350998 444408
rect 351054 444352 351059 444408
rect 214484 444350 351059 444352
rect 214484 444348 214490 444350
rect 350993 444347 351059 444350
rect 362217 443458 362283 443461
rect 362769 443460 362835 443461
rect 362534 443458 362540 443460
rect 362217 443456 362540 443458
rect 362217 443400 362222 443456
rect 362278 443400 362540 443456
rect 362217 443398 362540 443400
rect 362217 443395 362283 443398
rect 362534 443396 362540 443398
rect 362604 443396 362610 443460
rect 362718 443458 362724 443460
rect 362678 443398 362724 443458
rect 362788 443456 362835 443460
rect 362830 443400 362835 443456
rect 362718 443396 362724 443398
rect 362788 443396 362835 443400
rect 362902 443396 362908 443460
rect 362972 443458 362978 443460
rect 363045 443458 363111 443461
rect 362972 443456 363111 443458
rect 362972 443400 363050 443456
rect 363106 443400 363111 443456
rect 362972 443398 363111 443400
rect 362972 443396 362978 443398
rect 362769 443395 362835 443396
rect 363045 443395 363111 443398
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3325 423602 3391 423605
rect -960 423600 3391 423602
rect -960 423544 3330 423600
rect 3386 423544 3391 423600
rect -960 423542 3391 423544
rect -960 423452 480 423542
rect 3325 423539 3391 423542
rect 583520 418148 584960 418388
rect -960 410546 480 410636
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 583520 404820 584960 405060
rect -960 397490 480 397580
rect 3969 397490 4035 397493
rect -960 397488 4035 397490
rect -960 397432 3974 397488
rect 4030 397432 4035 397488
rect -960 397430 4035 397432
rect -960 397340 480 397430
rect 3969 397427 4035 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 579613 378450 579679 378453
rect 583520 378450 584960 378540
rect 579613 378448 584960 378450
rect 579613 378392 579618 378448
rect 579674 378392 584960 378448
rect 579613 378390 584960 378392
rect 579613 378387 579679 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 583520 364972 584960 365212
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 583520 351780 584960 352020
rect -960 345402 480 345492
rect 3877 345402 3943 345405
rect -960 345400 3943 345402
rect -960 345344 3882 345400
rect 3938 345344 3943 345400
rect -960 345342 3943 345344
rect -960 345252 480 345342
rect 3877 345339 3943 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 579981 325274 580047 325277
rect 583520 325274 584960 325364
rect 579981 325272 584960 325274
rect 579981 325216 579986 325272
rect 580042 325216 584960 325272
rect 579981 325214 584960 325216
rect 579981 325211 580047 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 583520 311932 584960 312172
rect 346117 309090 346183 309093
rect 365161 309090 365227 309093
rect 346117 309088 365227 309090
rect 346117 309032 346122 309088
rect 346178 309032 365166 309088
rect 365222 309032 365227 309088
rect 346117 309030 365227 309032
rect 346117 309027 346183 309030
rect 365161 309027 365227 309030
rect 216990 308892 216996 308956
rect 217060 308954 217066 308956
rect 275553 308954 275619 308957
rect 217060 308952 275619 308954
rect 217060 308896 275558 308952
rect 275614 308896 275619 308952
rect 217060 308894 275619 308896
rect 217060 308892 217066 308894
rect 275553 308891 275619 308894
rect 346393 308954 346459 308957
rect 367829 308954 367895 308957
rect 346393 308952 367895 308954
rect 346393 308896 346398 308952
rect 346454 308896 367834 308952
rect 367890 308896 367895 308952
rect 346393 308894 367895 308896
rect 346393 308891 346459 308894
rect 367829 308891 367895 308894
rect 217174 308756 217180 308820
rect 217244 308818 217250 308820
rect 276933 308818 276999 308821
rect 217244 308816 276999 308818
rect 217244 308760 276938 308816
rect 276994 308760 276999 308816
rect 217244 308758 276999 308760
rect 217244 308756 217250 308758
rect 276933 308755 276999 308758
rect 347037 308818 347103 308821
rect 367461 308818 367527 308821
rect 347037 308816 367527 308818
rect 347037 308760 347042 308816
rect 347098 308760 367466 308816
rect 367522 308760 367527 308816
rect 347037 308758 367527 308760
rect 347037 308755 347103 308758
rect 367461 308755 367527 308758
rect 217358 308620 217364 308684
rect 217428 308682 217434 308684
rect 278313 308682 278379 308685
rect 217428 308680 278379 308682
rect 217428 308624 278318 308680
rect 278374 308624 278379 308680
rect 217428 308622 278379 308624
rect 217428 308620 217434 308622
rect 278313 308619 278379 308622
rect 347313 308682 347379 308685
rect 370037 308682 370103 308685
rect 347313 308680 370103 308682
rect 347313 308624 347318 308680
rect 347374 308624 370042 308680
rect 370098 308624 370103 308680
rect 347313 308622 370103 308624
rect 347313 308619 347379 308622
rect 370037 308619 370103 308622
rect 75177 308546 75243 308549
rect 233417 308546 233483 308549
rect 75177 308544 233483 308546
rect 75177 308488 75182 308544
rect 75238 308488 233422 308544
rect 233478 308488 233483 308544
rect 75177 308486 233483 308488
rect 75177 308483 75243 308486
rect 233417 308483 233483 308486
rect 298461 308546 298527 308549
rect 358854 308546 358860 308548
rect 298461 308544 358860 308546
rect 298461 308488 298466 308544
rect 298522 308488 358860 308544
rect 298461 308486 358860 308488
rect 298461 308483 298527 308486
rect 358854 308484 358860 308486
rect 358924 308484 358930 308548
rect 35157 308410 35223 308413
rect 234521 308410 234587 308413
rect 35157 308408 234587 308410
rect 35157 308352 35162 308408
rect 35218 308352 234526 308408
rect 234582 308352 234587 308408
rect 35157 308350 234587 308352
rect 35157 308347 35223 308350
rect 234521 308347 234587 308350
rect 299105 308410 299171 308413
rect 360326 308410 360332 308412
rect 299105 308408 360332 308410
rect 299105 308352 299110 308408
rect 299166 308352 360332 308408
rect 299105 308350 360332 308352
rect 299105 308347 299171 308350
rect 360326 308348 360332 308350
rect 360396 308348 360402 308412
rect 353753 308274 353819 308277
rect 368013 308274 368079 308277
rect 353753 308272 368079 308274
rect 353753 308216 353758 308272
rect 353814 308216 368018 308272
rect 368074 308216 368079 308272
rect 353753 308214 368079 308216
rect 353753 308211 353819 308214
rect 368013 308211 368079 308214
rect 358997 308002 359063 308005
rect 467833 308002 467899 308005
rect 358997 308000 467899 308002
rect 358997 307944 359002 308000
rect 359058 307944 467838 308000
rect 467894 307944 467899 308000
rect 358997 307942 467899 307944
rect 358997 307939 359063 307942
rect 467833 307939 467899 307942
rect 361481 307866 361547 307869
rect 471973 307866 472039 307869
rect 361481 307864 472039 307866
rect 361481 307808 361486 307864
rect 361542 307808 471978 307864
rect 472034 307808 472039 307864
rect 361481 307806 472039 307808
rect 361481 307803 361547 307806
rect 471973 307803 472039 307806
rect 218646 306988 218652 307052
rect 218716 307050 218722 307052
rect 274633 307050 274699 307053
rect 218716 307048 274699 307050
rect 218716 306992 274638 307048
rect 274694 306992 274699 307048
rect 218716 306990 274699 306992
rect 218716 306988 218722 306990
rect 274633 306987 274699 306990
rect 312721 307050 312787 307053
rect 368974 307050 368980 307052
rect 312721 307048 368980 307050
rect 312721 306992 312726 307048
rect 312782 306992 368980 307048
rect 312721 306990 368980 306992
rect 312721 306987 312787 306990
rect 368974 306988 368980 306990
rect 369044 306988 369050 307052
rect -960 306234 480 306324
rect 3785 306234 3851 306237
rect -960 306232 3851 306234
rect -960 306176 3790 306232
rect 3846 306176 3851 306232
rect -960 306174 3851 306176
rect -960 306084 480 306174
rect 3785 306171 3851 306174
rect 219198 306172 219204 306236
rect 219268 306234 219274 306236
rect 274909 306234 274975 306237
rect 219268 306232 274975 306234
rect 219268 306176 274914 306232
rect 274970 306176 274975 306232
rect 219268 306174 274975 306176
rect 219268 306172 219274 306174
rect 274909 306171 274975 306174
rect 349153 306234 349219 306237
rect 370221 306234 370287 306237
rect 349153 306232 370287 306234
rect 349153 306176 349158 306232
rect 349214 306176 370226 306232
rect 370282 306176 370287 306232
rect 349153 306174 370287 306176
rect 349153 306171 349219 306174
rect 370221 306171 370287 306174
rect 216070 306036 216076 306100
rect 216140 306098 216146 306100
rect 275369 306098 275435 306101
rect 216140 306096 275435 306098
rect 216140 306040 275374 306096
rect 275430 306040 275435 306096
rect 216140 306038 275435 306040
rect 216140 306036 216146 306038
rect 275369 306035 275435 306038
rect 311157 306098 311223 306101
rect 400213 306098 400279 306101
rect 311157 306096 400279 306098
rect 311157 306040 311162 306096
rect 311218 306040 400218 306096
rect 400274 306040 400279 306096
rect 311157 306038 400279 306040
rect 311157 306035 311223 306038
rect 400213 306035 400279 306038
rect 215150 305900 215156 305964
rect 215220 305962 215226 305964
rect 275829 305962 275895 305965
rect 215220 305960 275895 305962
rect 215220 305904 275834 305960
rect 275890 305904 275895 305960
rect 215220 305902 275895 305904
rect 215220 305900 215226 305902
rect 275829 305899 275895 305902
rect 311341 305962 311407 305965
rect 404353 305962 404419 305965
rect 311341 305960 404419 305962
rect 311341 305904 311346 305960
rect 311402 305904 404358 305960
rect 404414 305904 404419 305960
rect 311341 305902 404419 305904
rect 311341 305899 311407 305902
rect 404353 305899 404419 305902
rect 214782 305764 214788 305828
rect 214852 305826 214858 305828
rect 276013 305826 276079 305829
rect 214852 305824 276079 305826
rect 214852 305768 276018 305824
rect 276074 305768 276079 305824
rect 214852 305766 276079 305768
rect 214852 305764 214858 305766
rect 276013 305763 276079 305766
rect 312537 305826 312603 305829
rect 407113 305826 407179 305829
rect 312537 305824 407179 305826
rect 312537 305768 312542 305824
rect 312598 305768 407118 305824
rect 407174 305768 407179 305824
rect 312537 305766 407179 305768
rect 312537 305763 312603 305766
rect 407113 305763 407179 305766
rect 217542 305628 217548 305692
rect 217612 305690 217618 305692
rect 281349 305690 281415 305693
rect 217612 305688 281415 305690
rect 217612 305632 281354 305688
rect 281410 305632 281415 305688
rect 217612 305630 281415 305632
rect 217612 305628 217618 305630
rect 281349 305627 281415 305630
rect 316309 305690 316375 305693
rect 429193 305690 429259 305693
rect 316309 305688 429259 305690
rect 316309 305632 316314 305688
rect 316370 305632 429198 305688
rect 429254 305632 429259 305688
rect 316309 305630 429259 305632
rect 316309 305627 316375 305630
rect 429193 305627 429259 305630
rect 309777 304330 309843 304333
rect 365110 304330 365116 304332
rect 309777 304328 365116 304330
rect 309777 304272 309782 304328
rect 309838 304272 365116 304328
rect 309777 304270 365116 304272
rect 309777 304267 309843 304270
rect 365110 304268 365116 304270
rect 365180 304268 365186 304332
rect 309961 304194 310027 304197
rect 367686 304194 367692 304196
rect 309961 304192 367692 304194
rect 309961 304136 309966 304192
rect 310022 304136 367692 304192
rect 309961 304134 367692 304136
rect 309961 304131 310027 304134
rect 367686 304132 367692 304134
rect 367756 304132 367762 304196
rect 216438 303316 216444 303380
rect 216508 303378 216514 303380
rect 276749 303378 276815 303381
rect 216508 303376 276815 303378
rect 216508 303320 276754 303376
rect 276810 303320 276815 303376
rect 216508 303318 276815 303320
rect 216508 303316 216514 303318
rect 276749 303315 276815 303318
rect 212942 303180 212948 303244
rect 213012 303242 213018 303244
rect 278129 303242 278195 303245
rect 213012 303240 278195 303242
rect 213012 303184 278134 303240
rect 278190 303184 278195 303240
rect 213012 303182 278195 303184
rect 213012 303180 213018 303182
rect 278129 303179 278195 303182
rect 212073 303106 212139 303109
rect 277393 303106 277459 303109
rect 212073 303104 277459 303106
rect 212073 303048 212078 303104
rect 212134 303048 277398 303104
rect 277454 303048 277459 303104
rect 212073 303046 277459 303048
rect 212073 303043 212139 303046
rect 277393 303043 277459 303046
rect 213269 302970 213335 302973
rect 279509 302970 279575 302973
rect 213269 302968 279575 302970
rect 213269 302912 213274 302968
rect 213330 302912 279514 302968
rect 279570 302912 279575 302968
rect 213269 302910 279575 302912
rect 213269 302907 213335 302910
rect 279509 302907 279575 302910
rect 211981 302834 212047 302837
rect 278773 302834 278839 302837
rect 211981 302832 278839 302834
rect 211981 302776 211986 302832
rect 212042 302776 278778 302832
rect 278834 302776 278839 302832
rect 211981 302774 278839 302776
rect 211981 302771 212047 302774
rect 278773 302771 278839 302774
rect 315481 302834 315547 302837
rect 392577 302834 392643 302837
rect 315481 302832 392643 302834
rect 315481 302776 315486 302832
rect 315542 302776 392582 302832
rect 392638 302776 392643 302832
rect 315481 302774 392643 302776
rect 315481 302771 315547 302774
rect 392577 302771 392643 302774
rect 214925 300114 214991 300117
rect 283189 300114 283255 300117
rect 214925 300112 283255 300114
rect 214925 300056 214930 300112
rect 214986 300056 283194 300112
rect 283250 300056 283255 300112
rect 214925 300054 283255 300056
rect 214925 300051 214991 300054
rect 283189 300051 283255 300054
rect 304073 298754 304139 298757
rect 365662 298754 365668 298756
rect 304073 298752 365668 298754
rect 304073 298696 304078 298752
rect 304134 298696 365668 298752
rect 304073 298694 365668 298696
rect 304073 298691 304139 298694
rect 365662 298692 365668 298694
rect 365732 298692 365738 298756
rect 583520 298604 584960 298844
rect -960 293178 480 293268
rect 3693 293178 3759 293181
rect -960 293176 3759 293178
rect -960 293120 3698 293176
rect 3754 293120 3759 293176
rect -960 293118 3759 293120
rect -960 293028 480 293118
rect 3693 293115 3759 293118
rect 303889 286378 303955 286381
rect 367134 286378 367140 286380
rect 303889 286376 367140 286378
rect 303889 286320 303894 286376
rect 303950 286320 367140 286376
rect 303889 286318 367140 286320
rect 303889 286315 303955 286318
rect 367134 286316 367140 286318
rect 367204 286316 367210 286380
rect 583520 285276 584960 285516
rect 302693 284882 302759 284885
rect 360326 284882 360332 284884
rect 302693 284880 360332 284882
rect 302693 284824 302698 284880
rect 302754 284824 360332 284880
rect 302693 284822 360332 284824
rect 302693 284819 302759 284822
rect 360326 284820 360332 284822
rect 360396 284820 360402 284884
rect -960 279972 480 280212
rect 216254 275164 216260 275228
rect 216324 275226 216330 275228
rect 273713 275226 273779 275229
rect 216324 275224 273779 275226
rect 216324 275168 273718 275224
rect 273774 275168 273779 275224
rect 216324 275166 273779 275168
rect 216324 275164 216330 275166
rect 273713 275163 273779 275166
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect 303797 269786 303863 269789
rect 369894 269786 369900 269788
rect 303797 269784 369900 269786
rect 303797 269728 303802 269784
rect 303858 269728 369900 269784
rect 303797 269726 369900 269728
rect 303797 269723 303863 269726
rect 369894 269724 369900 269726
rect 369964 269724 369970 269788
rect -960 267202 480 267292
rect 3233 267202 3299 267205
rect -960 267200 3299 267202
rect -960 267144 3238 267200
rect 3294 267144 3299 267200
rect -960 267142 3299 267144
rect -960 267052 480 267142
rect 3233 267139 3299 267142
rect 302601 267066 302667 267069
rect 363086 267066 363092 267068
rect 302601 267064 363092 267066
rect 302601 267008 302606 267064
rect 302662 267008 363092 267064
rect 302601 267006 363092 267008
rect 302601 267003 302667 267006
rect 363086 267004 363092 267006
rect 363156 267004 363162 267068
rect 214966 265508 214972 265572
rect 215036 265570 215042 265572
rect 273529 265570 273595 265573
rect 215036 265568 273595 265570
rect 215036 265512 273534 265568
rect 273590 265512 273595 265568
rect 215036 265510 273595 265512
rect 215036 265508 215042 265510
rect 273529 265507 273595 265510
rect 215886 262788 215892 262852
rect 215956 262850 215962 262852
rect 270493 262850 270559 262853
rect 215956 262848 270559 262850
rect 215956 262792 270498 262848
rect 270554 262792 270559 262848
rect 215956 262790 270559 262792
rect 215956 262788 215962 262790
rect 270493 262787 270559 262790
rect 329925 262850 329991 262853
rect 363454 262850 363460 262852
rect 329925 262848 363460 262850
rect 329925 262792 329930 262848
rect 329986 262792 363460 262848
rect 329925 262790 363460 262792
rect 329925 262787 329991 262790
rect 363454 262788 363460 262790
rect 363524 262788 363530 262852
rect 302509 260130 302575 260133
rect 359038 260130 359044 260132
rect 302509 260128 359044 260130
rect 302509 260072 302514 260128
rect 302570 260072 359044 260128
rect 302509 260070 359044 260072
rect 302509 260067 302575 260070
rect 359038 260068 359044 260070
rect 359108 260068 359114 260132
rect 583520 258756 584960 258996
rect 303613 254554 303679 254557
rect 368422 254554 368428 254556
rect 303613 254552 368428 254554
rect 303613 254496 303618 254552
rect 303674 254496 368428 254552
rect 303613 254494 368428 254496
rect 303613 254491 303679 254494
rect 368422 254492 368428 254494
rect 368492 254492 368498 254556
rect -960 254146 480 254236
rect 2773 254146 2839 254149
rect -960 254144 2839 254146
rect -960 254088 2778 254144
rect 2834 254088 2839 254144
rect -960 254086 2839 254088
rect -960 253996 480 254086
rect 2773 254083 2839 254086
rect 301129 250746 301195 250749
rect 360694 250746 360700 250748
rect 301129 250744 360700 250746
rect 301129 250688 301134 250744
rect 301190 250688 360700 250744
rect 301129 250686 360700 250688
rect 301129 250683 301195 250686
rect 360694 250684 360700 250686
rect 360764 250684 360770 250748
rect 317597 250610 317663 250613
rect 438853 250610 438919 250613
rect 317597 250608 438919 250610
rect 317597 250552 317602 250608
rect 317658 250552 438858 250608
rect 438914 250552 438919 250608
rect 317597 250550 438919 250552
rect 317597 250547 317663 250550
rect 438853 250547 438919 250550
rect 338205 250474 338271 250477
rect 546493 250474 546559 250477
rect 338205 250472 546559 250474
rect 338205 250416 338210 250472
rect 338266 250416 546498 250472
rect 546554 250416 546559 250472
rect 338205 250414 546559 250416
rect 338205 250411 338271 250414
rect 546493 250411 546559 250414
rect 213126 249052 213132 249116
rect 213196 249114 213202 249116
rect 273345 249114 273411 249117
rect 213196 249112 273411 249114
rect 213196 249056 273350 249112
rect 273406 249056 273411 249112
rect 213196 249054 273411 249056
rect 213196 249052 213202 249054
rect 273345 249051 273411 249054
rect 302325 249114 302391 249117
rect 364374 249114 364380 249116
rect 302325 249112 364380 249114
rect 302325 249056 302330 249112
rect 302386 249056 364380 249112
rect 302325 249054 364380 249056
rect 302325 249051 302391 249054
rect 364374 249052 364380 249054
rect 364444 249052 364450 249116
rect 295517 248162 295583 248165
rect 358118 248162 358124 248164
rect 295517 248160 358124 248162
rect 295517 248104 295522 248160
rect 295578 248104 358124 248160
rect 295517 248102 358124 248104
rect 295517 248099 295583 248102
rect 358118 248100 358124 248102
rect 358188 248100 358194 248164
rect 322933 248026 322999 248029
rect 465165 248026 465231 248029
rect 322933 248024 465231 248026
rect 322933 247968 322938 248024
rect 322994 247968 465170 248024
rect 465226 247968 465231 248024
rect 322933 247966 465231 247968
rect 322933 247963 322999 247966
rect 465165 247963 465231 247966
rect 323117 247890 323183 247893
rect 469213 247890 469279 247893
rect 323117 247888 469279 247890
rect 323117 247832 323122 247888
rect 323178 247832 469218 247888
rect 469274 247832 469279 247888
rect 323117 247830 469279 247832
rect 323117 247827 323183 247830
rect 469213 247827 469279 247830
rect 324497 247754 324563 247757
rect 473445 247754 473511 247757
rect 324497 247752 473511 247754
rect 324497 247696 324502 247752
rect 324558 247696 473450 247752
rect 473506 247696 473511 247752
rect 324497 247694 473511 247696
rect 324497 247691 324563 247694
rect 473445 247691 473511 247694
rect 324313 247618 324379 247621
rect 476113 247618 476179 247621
rect 324313 247616 476179 247618
rect 324313 247560 324318 247616
rect 324374 247560 476118 247616
rect 476174 247560 476179 247616
rect 324313 247558 476179 247560
rect 324313 247555 324379 247558
rect 476113 247555 476179 247558
rect 219014 246196 219020 246260
rect 219084 246258 219090 246260
rect 274633 246258 274699 246261
rect 219084 246256 274699 246258
rect 219084 246200 274638 246256
rect 274694 246200 274699 246256
rect 219084 246198 274699 246200
rect 219084 246196 219090 246198
rect 274633 246195 274699 246198
rect 302233 245578 302299 245581
rect 358302 245578 358308 245580
rect 302233 245576 358308 245578
rect 302233 245520 302238 245576
rect 302294 245520 358308 245576
rect 302233 245518 358308 245520
rect 302233 245515 302299 245518
rect 358302 245516 358308 245518
rect 358372 245516 358378 245580
rect 299473 245442 299539 245445
rect 359222 245442 359228 245444
rect 299473 245440 359228 245442
rect 299473 245384 299478 245440
rect 299534 245384 359228 245440
rect 299473 245382 359228 245384
rect 299473 245379 299539 245382
rect 359222 245380 359228 245382
rect 359292 245380 359298 245444
rect 583520 245428 584960 245668
rect 300853 245306 300919 245309
rect 356605 245306 356671 245309
rect 359406 245306 359412 245308
rect 300853 245304 356671 245306
rect 300853 245248 300858 245304
rect 300914 245248 356610 245304
rect 356666 245248 356671 245304
rect 300853 245246 356671 245248
rect 300853 245243 300919 245246
rect 356605 245243 356671 245246
rect 357022 245246 359412 245306
rect 296713 245170 296779 245173
rect 357022 245170 357082 245246
rect 359406 245244 359412 245246
rect 359476 245244 359482 245308
rect 296713 245168 357082 245170
rect 296713 245112 296718 245168
rect 296774 245112 357082 245168
rect 296713 245110 357082 245112
rect 357433 245170 357499 245173
rect 357934 245170 357940 245172
rect 357433 245168 357940 245170
rect 357433 245112 357438 245168
rect 357494 245112 357940 245168
rect 357433 245110 357940 245112
rect 296713 245107 296779 245110
rect 357433 245107 357499 245110
rect 357934 245108 357940 245110
rect 358004 245108 358010 245172
rect 295425 245034 295491 245037
rect 358486 245034 358492 245036
rect 295425 245032 358492 245034
rect 295425 244976 295430 245032
rect 295486 244976 358492 245032
rect 295425 244974 358492 244976
rect 295425 244971 295491 244974
rect 358486 244972 358492 244974
rect 358556 244972 358562 245036
rect 296897 244898 296963 244901
rect 360510 244898 360516 244900
rect 296897 244896 360516 244898
rect 296897 244840 296902 244896
rect 296958 244840 360516 244896
rect 296897 244838 360516 244840
rect 296897 244835 296963 244838
rect 360510 244836 360516 244838
rect 360580 244836 360586 244900
rect 356881 244762 356947 244765
rect 367318 244762 367324 244764
rect 356881 244760 367324 244762
rect 356881 244704 356886 244760
rect 356942 244704 367324 244760
rect 356881 244702 367324 244704
rect 356881 244699 356947 244702
rect 367318 244700 367324 244702
rect 367388 244700 367394 244764
rect 356605 244626 356671 244629
rect 363270 244626 363276 244628
rect 356605 244624 363276 244626
rect 356605 244568 356610 244624
rect 356666 244568 363276 244624
rect 356605 244566 363276 244568
rect 356605 244563 356671 244566
rect 363270 244564 363276 244566
rect 363340 244564 363346 244628
rect 218094 243340 218100 243404
rect 218164 243402 218170 243404
rect 218421 243402 218487 243405
rect 218164 243400 218487 243402
rect 218164 243344 218426 243400
rect 218482 243344 218487 243400
rect 218164 243342 218487 243344
rect 218164 243340 218170 243342
rect 218421 243339 218487 243342
rect -960 241090 480 241180
rect 3601 241090 3667 241093
rect -960 241088 3667 241090
rect -960 241032 3606 241088
rect 3662 241032 3667 241088
rect -960 241030 3667 241032
rect -960 240940 480 241030
rect 3601 241027 3667 241030
rect 580625 232386 580691 232389
rect 583520 232386 584960 232476
rect 580625 232384 584960 232386
rect 580625 232328 580630 232384
rect 580686 232328 584960 232384
rect 580625 232326 584960 232328
rect 580625 232323 580691 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 583520 205580 584960 205820
rect -960 201922 480 202012
rect 3693 201922 3759 201925
rect -960 201920 3759 201922
rect -960 201864 3698 201920
rect 3754 201864 3759 201920
rect -960 201862 3759 201864
rect -960 201772 480 201862
rect 3693 201859 3759 201862
rect 217409 196890 217475 196893
rect 219390 196890 220064 196924
rect 217409 196888 220064 196890
rect 217409 196832 217414 196888
rect 217470 196864 220064 196888
rect 217470 196832 219450 196864
rect 217409 196830 219450 196832
rect 217409 196827 217475 196830
rect 217501 195938 217567 195941
rect 219390 195938 220064 195972
rect 217501 195936 220064 195938
rect 217501 195880 217506 195936
rect 217562 195912 220064 195936
rect 217562 195880 219450 195912
rect 217501 195878 219450 195880
rect 217501 195875 217567 195878
rect 217041 193762 217107 193765
rect 219390 193762 220064 193796
rect 217041 193760 220064 193762
rect 217041 193704 217046 193760
rect 217102 193736 220064 193760
rect 217102 193704 219450 193736
rect 217041 193702 219450 193704
rect 217041 193699 217107 193702
rect 216673 192810 216739 192813
rect 219390 192810 220064 192844
rect 216673 192808 220064 192810
rect 216673 192752 216678 192808
rect 216734 192784 220064 192808
rect 216734 192752 219450 192784
rect 216673 192750 219450 192752
rect 216673 192747 216739 192750
rect 580533 192538 580599 192541
rect 583520 192538 584960 192628
rect 580533 192536 584960 192538
rect 580533 192480 580538 192536
rect 580594 192480 584960 192536
rect 580533 192478 584960 192480
rect 580533 192475 580599 192478
rect 583520 192388 584960 192478
rect 218605 191042 218671 191045
rect 219390 191042 220064 191076
rect 218605 191040 220064 191042
rect 218605 190984 218610 191040
rect 218666 191016 220064 191040
rect 218666 190984 219450 191016
rect 218605 190982 219450 190984
rect 218605 190979 218671 190982
rect 218513 189954 218579 189957
rect 219390 189954 220064 189988
rect 218513 189952 220064 189954
rect 218513 189896 218518 189952
rect 218574 189928 220064 189952
rect 218574 189896 219450 189928
rect 218513 189894 219450 189896
rect 218513 189891 218579 189894
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 216673 188186 216739 188189
rect 219390 188186 220064 188220
rect 216673 188184 220064 188186
rect 216673 188128 216678 188184
rect 216734 188160 220064 188184
rect 216734 188128 219450 188160
rect 216673 188126 219450 188128
rect 216673 188123 216739 188126
rect 583520 179060 584960 179300
rect 369158 177244 369164 177308
rect 369228 177306 369234 177308
rect 581085 177306 581151 177309
rect 369228 177304 581151 177306
rect 369228 177248 581090 177304
rect 581146 177248 581151 177304
rect 369228 177246 581151 177248
rect 369228 177244 369234 177246
rect 581085 177243 581151 177246
rect -960 175796 480 176036
rect 217133 169962 217199 169965
rect 219390 169962 220064 169996
rect 217133 169960 220064 169962
rect 217133 169904 217138 169960
rect 217194 169936 220064 169960
rect 217194 169904 219450 169936
rect 217133 169902 219450 169904
rect 217133 169899 217199 169902
rect 217593 168330 217659 168333
rect 219390 168330 220064 168364
rect 217593 168328 220064 168330
rect 217593 168272 217598 168328
rect 217654 168304 220064 168328
rect 217654 168272 219450 168304
rect 217593 168270 219450 168272
rect 217593 168267 217659 168270
rect 217685 168058 217751 168061
rect 219390 168058 220064 168092
rect 217685 168056 220064 168058
rect 217685 168000 217690 168056
rect 217746 168032 220064 168056
rect 217746 168000 219450 168032
rect 217685 167998 219450 168000
rect 217685 167995 217751 167998
rect 583520 165732 584960 165972
rect -960 162890 480 162980
rect 218094 162890 218100 162892
rect -960 162830 218100 162890
rect -960 162740 480 162830
rect 218094 162828 218100 162830
rect 218164 162828 218170 162892
rect 273345 159900 273411 159901
rect 278129 159900 278195 159901
rect 273312 159898 273318 159900
rect 273254 159838 273318 159898
rect 273382 159896 273411 159900
rect 278072 159898 278078 159900
rect 273406 159840 273411 159896
rect 273312 159836 273318 159838
rect 273382 159836 273411 159840
rect 278038 159838 278078 159898
rect 278142 159896 278195 159900
rect 278190 159840 278195 159896
rect 278072 159836 278078 159838
rect 278142 159836 278195 159840
rect 273345 159835 273411 159836
rect 278129 159835 278195 159836
rect 261109 159764 261175 159765
rect 261072 159762 261078 159764
rect 261018 159702 261078 159762
rect 261142 159760 261175 159764
rect 261170 159704 261175 159760
rect 261072 159700 261078 159702
rect 261142 159700 261175 159704
rect 261109 159699 261175 159700
rect 355317 159762 355383 159765
rect 357709 159762 357775 159765
rect 355317 159760 357775 159762
rect 355317 159704 355322 159760
rect 355378 159704 357714 159760
rect 357770 159704 357775 159760
rect 355317 159702 357775 159704
rect 355317 159699 355383 159702
rect 357709 159699 357775 159702
rect 275829 159628 275895 159629
rect 277025 159628 277091 159629
rect 279233 159628 279299 159629
rect 260664 159564 260670 159628
rect 260734 159626 260740 159628
rect 275760 159626 275766 159628
rect 260734 159566 267750 159626
rect 275738 159566 275766 159626
rect 260734 159564 260740 159566
rect 267690 159354 267750 159566
rect 275760 159564 275766 159566
rect 275830 159624 275895 159628
rect 276984 159626 276990 159628
rect 275830 159568 275834 159624
rect 275890 159568 275895 159624
rect 275830 159564 275895 159568
rect 276934 159566 276990 159626
rect 277054 159624 277091 159628
rect 279160 159626 279166 159628
rect 277086 159568 277091 159624
rect 276984 159564 276990 159566
rect 277054 159564 277091 159568
rect 279142 159566 279166 159626
rect 279160 159564 279166 159566
rect 279230 159624 279299 159628
rect 279230 159568 279238 159624
rect 279294 159568 279299 159624
rect 279230 159564 279299 159568
rect 275829 159563 275895 159564
rect 277025 159563 277091 159564
rect 279233 159563 279299 159564
rect 366449 159490 366515 159493
rect 354630 159488 366515 159490
rect 354630 159432 366454 159488
rect 366510 159432 366515 159488
rect 354630 159430 366515 159432
rect 354630 159354 354690 159430
rect 366449 159427 366515 159430
rect 267690 159294 354690 159354
rect 357433 159354 357499 159357
rect 357934 159354 357940 159356
rect 357433 159352 357940 159354
rect 357433 159296 357438 159352
rect 357494 159296 357940 159352
rect 357433 159294 357940 159296
rect 357433 159291 357499 159294
rect 357934 159292 357940 159294
rect 358004 159292 358010 159356
rect 360694 159292 360700 159356
rect 360764 159354 360770 159356
rect 361113 159354 361179 159357
rect 360764 159352 361179 159354
rect 360764 159296 361118 159352
rect 361174 159296 361179 159352
rect 360764 159294 361179 159296
rect 360764 159292 360770 159294
rect 361113 159291 361179 159294
rect 363270 159292 363276 159356
rect 363340 159354 363346 159356
rect 363873 159354 363939 159357
rect 363340 159352 363939 159354
rect 363340 159296 363878 159352
rect 363934 159296 363939 159352
rect 363340 159294 363939 159296
rect 363340 159292 363346 159294
rect 363873 159291 363939 159294
rect 259494 159156 259500 159220
rect 259564 159218 259570 159220
rect 367921 159218 367987 159221
rect 259564 159216 367987 159218
rect 259564 159160 367926 159216
rect 367982 159160 367987 159216
rect 259564 159158 367987 159160
rect 259564 159156 259570 159158
rect 367921 159155 367987 159158
rect 254526 159020 254532 159084
rect 254596 159082 254602 159084
rect 368013 159082 368079 159085
rect 254596 159080 368079 159082
rect 254596 159024 368018 159080
rect 368074 159024 368079 159080
rect 254596 159022 368079 159024
rect 254596 159020 254602 159022
rect 368013 159019 368079 159022
rect 253606 158884 253612 158948
rect 253676 158946 253682 158948
rect 370681 158946 370747 158949
rect 253676 158944 370747 158946
rect 253676 158888 370686 158944
rect 370742 158888 370747 158944
rect 253676 158886 370747 158888
rect 253676 158884 253682 158886
rect 370681 158883 370747 158886
rect 243118 158748 243124 158812
rect 243188 158810 243194 158812
rect 367829 158810 367895 158813
rect 243188 158808 367895 158810
rect 243188 158752 367834 158808
rect 367890 158752 367895 158808
rect 243188 158750 367895 158752
rect 243188 158748 243194 158750
rect 367829 158747 367895 158750
rect 216990 158612 216996 158676
rect 217060 158674 217066 158676
rect 220813 158674 220879 158677
rect 217060 158672 220879 158674
rect 217060 158616 220818 158672
rect 220874 158616 220879 158672
rect 217060 158614 220879 158616
rect 217060 158612 217066 158614
rect 220813 158611 220879 158614
rect 238109 158676 238175 158677
rect 239581 158676 239647 158677
rect 238109 158672 238156 158676
rect 238220 158674 238226 158676
rect 238109 158616 238114 158672
rect 238109 158612 238156 158616
rect 238220 158614 238266 158674
rect 239581 158672 239628 158676
rect 239692 158674 239698 158676
rect 239581 158616 239586 158672
rect 238220 158612 238226 158614
rect 239581 158612 239628 158616
rect 239692 158614 239738 158674
rect 239692 158612 239698 158614
rect 241830 158612 241836 158676
rect 241900 158674 241906 158676
rect 242433 158674 242499 158677
rect 241900 158672 242499 158674
rect 241900 158616 242438 158672
rect 242494 158616 242499 158672
rect 241900 158614 242499 158616
rect 241900 158612 241906 158614
rect 238109 158611 238175 158612
rect 239581 158611 239647 158612
rect 242433 158611 242499 158614
rect 244222 158612 244228 158676
rect 244292 158674 244298 158676
rect 244641 158674 244707 158677
rect 245561 158676 245627 158677
rect 248321 158676 248387 158677
rect 252369 158676 252435 158677
rect 255865 158676 255931 158677
rect 245510 158674 245516 158676
rect 244292 158672 244707 158674
rect 244292 158616 244646 158672
rect 244702 158616 244707 158672
rect 244292 158614 244707 158616
rect 245470 158614 245516 158674
rect 245580 158672 245627 158676
rect 248270 158674 248276 158676
rect 245622 158616 245627 158672
rect 244292 158612 244298 158614
rect 244641 158611 244707 158614
rect 245510 158612 245516 158614
rect 245580 158612 245627 158616
rect 248230 158614 248276 158674
rect 248340 158672 248387 158676
rect 252318 158674 252324 158676
rect 248382 158616 248387 158672
rect 248270 158612 248276 158614
rect 248340 158612 248387 158616
rect 252278 158614 252324 158674
rect 252388 158672 252435 158676
rect 255814 158674 255820 158676
rect 252430 158616 252435 158672
rect 252318 158612 252324 158614
rect 252388 158612 252435 158616
rect 255774 158614 255820 158674
rect 255884 158672 255931 158676
rect 255926 158616 255931 158672
rect 255814 158612 255820 158614
rect 255884 158612 255931 158616
rect 257102 158612 257108 158676
rect 257172 158674 257178 158676
rect 257245 158674 257311 158677
rect 261753 158676 261819 158677
rect 265433 158676 265499 158677
rect 265985 158676 266051 158677
rect 266537 158676 266603 158677
rect 268745 158676 268811 158677
rect 261702 158674 261708 158676
rect 257172 158672 257311 158674
rect 257172 158616 257250 158672
rect 257306 158616 257311 158672
rect 257172 158614 257311 158616
rect 261662 158614 261708 158674
rect 261772 158672 261819 158676
rect 265382 158674 265388 158676
rect 261814 158616 261819 158672
rect 257172 158612 257178 158614
rect 245561 158611 245627 158612
rect 248321 158611 248387 158612
rect 252369 158611 252435 158612
rect 255865 158611 255931 158612
rect 257245 158611 257311 158614
rect 261702 158612 261708 158614
rect 261772 158612 261819 158616
rect 265342 158614 265388 158674
rect 265452 158672 265499 158676
rect 265934 158674 265940 158676
rect 265494 158616 265499 158672
rect 265382 158612 265388 158614
rect 265452 158612 265499 158616
rect 265894 158614 265940 158674
rect 266004 158672 266051 158676
rect 266486 158674 266492 158676
rect 266046 158616 266051 158672
rect 265934 158612 265940 158614
rect 266004 158612 266051 158616
rect 266446 158614 266492 158674
rect 266556 158672 266603 158676
rect 268694 158674 268700 158676
rect 266598 158616 266603 158672
rect 266486 158612 266492 158614
rect 266556 158612 266603 158616
rect 268654 158614 268700 158674
rect 268764 158672 268811 158676
rect 268806 158616 268811 158672
rect 268694 158612 268700 158614
rect 268764 158612 268811 158616
rect 269798 158612 269804 158676
rect 269868 158674 269874 158676
rect 269941 158674 270007 158677
rect 270953 158676 271019 158677
rect 272241 158676 272307 158677
rect 274449 158676 274515 158677
rect 276105 158676 276171 158677
rect 281073 158676 281139 158677
rect 288249 158676 288315 158677
rect 291009 158676 291075 158677
rect 293585 158676 293651 158677
rect 295977 158676 296043 158677
rect 298553 158676 298619 158677
rect 300945 158676 301011 158677
rect 303521 158676 303587 158677
rect 306097 158676 306163 158677
rect 308673 158676 308739 158677
rect 311065 158676 311131 158677
rect 313457 158676 313523 158677
rect 315849 158676 315915 158677
rect 318609 158676 318675 158677
rect 321001 158676 321067 158677
rect 323393 158676 323459 158677
rect 325969 158676 326035 158677
rect 270902 158674 270908 158676
rect 269868 158672 270007 158674
rect 269868 158616 269946 158672
rect 270002 158616 270007 158672
rect 269868 158614 270007 158616
rect 270862 158614 270908 158674
rect 270972 158672 271019 158676
rect 272190 158674 272196 158676
rect 271014 158616 271019 158672
rect 269868 158612 269874 158614
rect 261753 158611 261819 158612
rect 265433 158611 265499 158612
rect 265985 158611 266051 158612
rect 266537 158611 266603 158612
rect 268745 158611 268811 158612
rect 269941 158611 270007 158614
rect 270902 158612 270908 158614
rect 270972 158612 271019 158616
rect 272150 158614 272196 158674
rect 272260 158672 272307 158676
rect 274398 158674 274404 158676
rect 272302 158616 272307 158672
rect 272190 158612 272196 158614
rect 272260 158612 272307 158616
rect 274358 158614 274404 158674
rect 274468 158672 274515 158676
rect 276054 158674 276060 158676
rect 274510 158616 274515 158672
rect 274398 158612 274404 158614
rect 274468 158612 274515 158616
rect 276014 158614 276060 158674
rect 276124 158672 276171 158676
rect 281022 158674 281028 158676
rect 276166 158616 276171 158672
rect 276054 158612 276060 158614
rect 276124 158612 276171 158616
rect 280982 158614 281028 158674
rect 281092 158672 281139 158676
rect 288198 158674 288204 158676
rect 281134 158616 281139 158672
rect 281022 158612 281028 158614
rect 281092 158612 281139 158616
rect 288158 158614 288204 158674
rect 288268 158672 288315 158676
rect 290958 158674 290964 158676
rect 288310 158616 288315 158672
rect 288198 158612 288204 158614
rect 288268 158612 288315 158616
rect 290918 158614 290964 158674
rect 291028 158672 291075 158676
rect 293534 158674 293540 158676
rect 291070 158616 291075 158672
rect 290958 158612 290964 158614
rect 291028 158612 291075 158616
rect 293494 158614 293540 158674
rect 293604 158672 293651 158676
rect 295926 158674 295932 158676
rect 293646 158616 293651 158672
rect 293534 158612 293540 158614
rect 293604 158612 293651 158616
rect 295886 158614 295932 158674
rect 295996 158672 296043 158676
rect 298502 158674 298508 158676
rect 296038 158616 296043 158672
rect 295926 158612 295932 158614
rect 295996 158612 296043 158616
rect 298462 158614 298508 158674
rect 298572 158672 298619 158676
rect 300894 158674 300900 158676
rect 298614 158616 298619 158672
rect 298502 158612 298508 158614
rect 298572 158612 298619 158616
rect 300854 158614 300900 158674
rect 300964 158672 301011 158676
rect 303470 158674 303476 158676
rect 301006 158616 301011 158672
rect 300894 158612 300900 158614
rect 300964 158612 301011 158616
rect 303430 158614 303476 158674
rect 303540 158672 303587 158676
rect 306046 158674 306052 158676
rect 303582 158616 303587 158672
rect 303470 158612 303476 158614
rect 303540 158612 303587 158616
rect 306006 158614 306052 158674
rect 306116 158672 306163 158676
rect 308622 158674 308628 158676
rect 306158 158616 306163 158672
rect 306046 158612 306052 158614
rect 306116 158612 306163 158616
rect 308582 158614 308628 158674
rect 308692 158672 308739 158676
rect 311014 158674 311020 158676
rect 308734 158616 308739 158672
rect 308622 158612 308628 158614
rect 308692 158612 308739 158616
rect 310974 158614 311020 158674
rect 311084 158672 311131 158676
rect 313406 158674 313412 158676
rect 311126 158616 311131 158672
rect 311014 158612 311020 158614
rect 311084 158612 311131 158616
rect 313366 158614 313412 158674
rect 313476 158672 313523 158676
rect 315798 158674 315804 158676
rect 313518 158616 313523 158672
rect 313406 158612 313412 158614
rect 313476 158612 313523 158616
rect 315758 158614 315804 158674
rect 315868 158672 315915 158676
rect 318558 158674 318564 158676
rect 315910 158616 315915 158672
rect 315798 158612 315804 158614
rect 315868 158612 315915 158616
rect 318518 158614 318564 158674
rect 318628 158672 318675 158676
rect 320950 158674 320956 158676
rect 318670 158616 318675 158672
rect 318558 158612 318564 158614
rect 318628 158612 318675 158616
rect 320910 158614 320956 158674
rect 321020 158672 321067 158676
rect 323342 158674 323348 158676
rect 321062 158616 321067 158672
rect 320950 158612 320956 158614
rect 321020 158612 321067 158616
rect 323302 158614 323348 158674
rect 323412 158672 323459 158676
rect 325918 158674 325924 158676
rect 323454 158616 323459 158672
rect 323342 158612 323348 158614
rect 323412 158612 323459 158616
rect 325878 158614 325924 158674
rect 325988 158672 326035 158676
rect 326030 158616 326035 158672
rect 325918 158612 325924 158614
rect 325988 158612 326035 158616
rect 270953 158611 271019 158612
rect 272241 158611 272307 158612
rect 274449 158611 274515 158612
rect 276105 158611 276171 158612
rect 281073 158611 281139 158612
rect 288249 158611 288315 158612
rect 291009 158611 291075 158612
rect 293585 158611 293651 158612
rect 295977 158611 296043 158612
rect 298553 158611 298619 158612
rect 300945 158611 301011 158612
rect 303521 158611 303587 158612
rect 306097 158611 306163 158612
rect 308673 158611 308739 158612
rect 311065 158611 311131 158612
rect 313457 158611 313523 158612
rect 315849 158611 315915 158612
rect 318609 158611 318675 158612
rect 321001 158611 321067 158612
rect 323393 158611 323459 158612
rect 325969 158611 326035 158612
rect 218881 158538 218947 158541
rect 224953 158538 225019 158541
rect 218881 158536 225019 158538
rect 218881 158480 218886 158536
rect 218942 158480 224958 158536
rect 225014 158480 225019 158536
rect 218881 158478 225019 158480
rect 218881 158475 218947 158478
rect 224953 158475 225019 158478
rect 236126 158476 236132 158540
rect 236196 158538 236202 158540
rect 365161 158538 365227 158541
rect 236196 158536 365227 158538
rect 236196 158480 365166 158536
rect 365222 158480 365227 158536
rect 236196 158478 365227 158480
rect 236196 158476 236202 158478
rect 365161 158475 365227 158478
rect 216070 158340 216076 158404
rect 216140 158402 216146 158404
rect 219433 158402 219499 158405
rect 216140 158400 219499 158402
rect 216140 158344 219438 158400
rect 219494 158344 219499 158400
rect 216140 158342 219499 158344
rect 216140 158340 216146 158342
rect 219433 158339 219499 158342
rect 258206 158340 258212 158404
rect 258276 158402 258282 158404
rect 367553 158402 367619 158405
rect 258276 158400 367619 158402
rect 258276 158344 367558 158400
rect 367614 158344 367619 158400
rect 258276 158342 367619 158344
rect 258276 158340 258282 158342
rect 367553 158339 367619 158342
rect 217174 158204 217180 158268
rect 217244 158266 217250 158268
rect 227713 158266 227779 158269
rect 217244 158264 227779 158266
rect 217244 158208 227718 158264
rect 227774 158208 227779 158264
rect 217244 158206 227779 158208
rect 217244 158204 217250 158206
rect 227713 158203 227779 158206
rect 240542 158204 240548 158268
rect 240612 158266 240618 158268
rect 241421 158266 241487 158269
rect 240612 158264 241487 158266
rect 240612 158208 241426 158264
rect 241482 158208 241487 158264
rect 240612 158206 241487 158208
rect 240612 158204 240618 158206
rect 241421 158203 241487 158206
rect 258574 158204 258580 158268
rect 258644 158266 258650 158268
rect 366541 158266 366607 158269
rect 258644 158264 366607 158266
rect 258644 158208 366546 158264
rect 366602 158208 366607 158264
rect 258644 158206 366607 158208
rect 258644 158204 258650 158206
rect 366541 158203 366607 158206
rect 217358 158068 217364 158132
rect 217428 158130 217434 158132
rect 234613 158130 234679 158133
rect 217428 158128 234679 158130
rect 217428 158072 234618 158128
rect 234674 158072 234679 158128
rect 217428 158070 234679 158072
rect 217428 158068 217434 158070
rect 234613 158067 234679 158070
rect 262622 158068 262628 158132
rect 262692 158130 262698 158132
rect 369117 158130 369183 158133
rect 262692 158128 369183 158130
rect 262692 158072 369122 158128
rect 369178 158072 369183 158128
rect 262692 158070 369183 158072
rect 262692 158068 262698 158070
rect 369117 158067 369183 158070
rect 214782 157932 214788 157996
rect 214852 157994 214858 157996
rect 223573 157994 223639 157997
rect 234705 157994 234771 157997
rect 246665 157996 246731 157997
rect 246614 157994 246620 157996
rect 214852 157992 223639 157994
rect 214852 157936 223578 157992
rect 223634 157936 223639 157992
rect 214852 157934 223639 157936
rect 214852 157932 214858 157934
rect 223573 157931 223639 157934
rect 229050 157992 234771 157994
rect 229050 157936 234710 157992
rect 234766 157936 234771 157992
rect 229050 157934 234771 157936
rect 246574 157934 246620 157994
rect 246684 157992 246731 157996
rect 246726 157936 246731 157992
rect 212942 157796 212948 157860
rect 213012 157858 213018 157860
rect 229050 157858 229110 157934
rect 234705 157931 234771 157934
rect 246614 157932 246620 157934
rect 246684 157932 246731 157936
rect 247718 157932 247724 157996
rect 247788 157994 247794 157996
rect 247953 157994 248019 157997
rect 247788 157992 248019 157994
rect 247788 157936 247958 157992
rect 248014 157936 248019 157992
rect 247788 157934 248019 157936
rect 247788 157932 247794 157934
rect 246665 157931 246731 157932
rect 247953 157931 248019 157934
rect 250846 157932 250852 157996
rect 250916 157994 250922 157996
rect 251081 157994 251147 157997
rect 250916 157992 251147 157994
rect 250916 157936 251086 157992
rect 251142 157936 251147 157992
rect 250916 157934 251147 157936
rect 250916 157932 250922 157934
rect 251081 157931 251147 157934
rect 267038 157932 267044 157996
rect 267108 157994 267114 157996
rect 370497 157994 370563 157997
rect 267108 157992 370563 157994
rect 267108 157936 370502 157992
rect 370558 157936 370563 157992
rect 267108 157934 370563 157936
rect 267108 157932 267114 157934
rect 370497 157931 370563 157934
rect 248689 157860 248755 157861
rect 248638 157858 248644 157860
rect 213012 157798 229110 157858
rect 248598 157798 248644 157858
rect 248708 157856 248755 157860
rect 248750 157800 248755 157856
rect 213012 157796 213018 157798
rect 248638 157796 248644 157798
rect 248708 157796 248755 157800
rect 250110 157796 250116 157860
rect 250180 157858 250186 157860
rect 250437 157858 250503 157861
rect 250180 157856 250503 157858
rect 250180 157800 250442 157856
rect 250498 157800 250503 157856
rect 250180 157798 250503 157800
rect 250180 157796 250186 157798
rect 248689 157795 248755 157796
rect 250437 157795 250503 157798
rect 251398 157796 251404 157860
rect 251468 157858 251474 157860
rect 252461 157858 252527 157861
rect 253473 157860 253539 157861
rect 253422 157858 253428 157860
rect 251468 157856 252527 157858
rect 251468 157800 252466 157856
rect 252522 157800 252527 157856
rect 251468 157798 252527 157800
rect 253382 157798 253428 157858
rect 253492 157856 253539 157860
rect 253534 157800 253539 157856
rect 251468 157796 251474 157798
rect 252461 157795 252527 157798
rect 253422 157796 253428 157798
rect 253492 157796 253539 157800
rect 263910 157796 263916 157860
rect 263980 157858 263986 157860
rect 355317 157858 355383 157861
rect 263980 157856 355383 157858
rect 263980 157800 355322 157856
rect 355378 157800 355383 157856
rect 263980 157798 355383 157800
rect 263980 157796 263986 157798
rect 253473 157795 253539 157796
rect 355317 157795 355383 157798
rect 268377 157724 268443 157725
rect 271321 157724 271387 157725
rect 273713 157724 273779 157725
rect 278497 157724 278563 157725
rect 268326 157722 268332 157724
rect 268286 157662 268332 157722
rect 268396 157720 268443 157724
rect 271270 157722 271276 157724
rect 268438 157664 268443 157720
rect 268326 157660 268332 157662
rect 268396 157660 268443 157664
rect 271230 157662 271276 157722
rect 271340 157720 271387 157724
rect 273662 157722 273668 157724
rect 271382 157664 271387 157720
rect 271270 157660 271276 157662
rect 271340 157660 271387 157664
rect 273622 157662 273668 157722
rect 273732 157720 273779 157724
rect 278446 157722 278452 157724
rect 273774 157664 273779 157720
rect 273662 157660 273668 157662
rect 273732 157660 273779 157664
rect 278406 157662 278452 157722
rect 278516 157720 278563 157724
rect 278558 157664 278563 157720
rect 278446 157660 278452 157662
rect 278516 157660 278563 157664
rect 268377 157659 268443 157660
rect 271321 157659 271387 157660
rect 273713 157659 273779 157660
rect 278497 157659 278563 157660
rect 256233 157588 256299 157589
rect 256182 157586 256188 157588
rect 256142 157526 256188 157586
rect 256252 157584 256299 157588
rect 256294 157528 256299 157584
rect 256182 157524 256188 157526
rect 256252 157524 256299 157528
rect 263542 157524 263548 157588
rect 263612 157586 263618 157588
rect 263685 157586 263751 157589
rect 283649 157588 283715 157589
rect 286041 157588 286107 157589
rect 283598 157586 283604 157588
rect 263612 157584 263751 157586
rect 263612 157528 263690 157584
rect 263746 157528 263751 157584
rect 263612 157526 263751 157528
rect 283558 157526 283604 157586
rect 283668 157584 283715 157588
rect 285990 157586 285996 157588
rect 283710 157528 283715 157584
rect 263612 157524 263618 157526
rect 256233 157523 256299 157524
rect 263685 157523 263751 157526
rect 283598 157524 283604 157526
rect 283668 157524 283715 157528
rect 285950 157526 285996 157586
rect 286060 157584 286107 157588
rect 286102 157528 286107 157584
rect 285990 157524 285996 157526
rect 286060 157524 286107 157528
rect 283649 157523 283715 157524
rect 286041 157523 286107 157524
rect 237230 157388 237236 157452
rect 237300 157450 237306 157452
rect 367461 157450 367527 157453
rect 237300 157448 367527 157450
rect 237300 157392 367466 157448
rect 367522 157392 367527 157448
rect 237300 157390 367527 157392
rect 237300 157388 237306 157390
rect 367461 157387 367527 157390
rect 213545 155954 213611 155957
rect 253933 155954 253999 155957
rect 213545 155952 253999 155954
rect 213545 155896 213550 155952
rect 213606 155896 253938 155952
rect 253994 155896 253999 155952
rect 213545 155894 253999 155896
rect 213545 155891 213611 155894
rect 253933 155891 253999 155894
rect 211061 155818 211127 155821
rect 255313 155818 255379 155821
rect 211061 155816 255379 155818
rect 211061 155760 211066 155816
rect 211122 155760 255318 155816
rect 255374 155760 255379 155816
rect 211061 155758 255379 155760
rect 211061 155755 211127 155758
rect 255313 155755 255379 155758
rect 212349 155682 212415 155685
rect 259545 155682 259611 155685
rect 212349 155680 259611 155682
rect 212349 155624 212354 155680
rect 212410 155624 259550 155680
rect 259606 155624 259611 155680
rect 212349 155622 259611 155624
rect 212349 155619 212415 155622
rect 259545 155619 259611 155622
rect 210877 155546 210943 155549
rect 267825 155546 267891 155549
rect 210877 155544 267891 155546
rect 210877 155488 210882 155544
rect 210938 155488 267830 155544
rect 267886 155488 267891 155544
rect 210877 155486 267891 155488
rect 210877 155483 210943 155486
rect 267825 155483 267891 155486
rect 210969 155410 211035 155413
rect 269113 155410 269179 155413
rect 210969 155408 269179 155410
rect 210969 155352 210974 155408
rect 211030 155352 269118 155408
rect 269174 155352 269179 155408
rect 210969 155350 269179 155352
rect 210969 155347 211035 155350
rect 269113 155347 269179 155350
rect 213177 155274 213243 155277
rect 274633 155274 274699 155277
rect 213177 155272 274699 155274
rect 213177 155216 213182 155272
rect 213238 155216 274638 155272
rect 274694 155216 274699 155272
rect 213177 155214 274699 155216
rect 213177 155211 213243 155214
rect 274633 155211 274699 155214
rect 580441 152690 580507 152693
rect 583520 152690 584960 152780
rect 580441 152688 584960 152690
rect 580441 152632 580446 152688
rect 580502 152632 584960 152688
rect 580441 152630 584960 152632
rect 580441 152627 580507 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3509 149834 3575 149837
rect -960 149832 3575 149834
rect -960 149776 3514 149832
rect 3570 149776 3575 149832
rect -960 149774 3575 149776
rect -960 149684 480 149774
rect 3509 149771 3575 149774
rect 583520 139212 584960 139452
rect -960 136778 480 136868
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 580349 112842 580415 112845
rect 583520 112842 584960 112932
rect 580349 112840 584960 112842
rect 580349 112784 580354 112840
rect 580410 112784 584960 112840
rect 580349 112782 584960 112784
rect 580349 112779 580415 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect -960 110606 6930 110666
rect -960 110516 480 110606
rect 6870 110530 6930 110606
rect 214414 110530 214420 110532
rect 6870 110470 214420 110530
rect 214414 110468 214420 110470
rect 214484 110468 214490 110532
rect 583520 99364 584960 99604
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 583520 86036 584960 86276
rect -960 84690 480 84780
rect -960 84630 6930 84690
rect -960 84540 480 84630
rect 6870 84282 6930 84630
rect 362534 84282 362540 84284
rect 6870 84222 362540 84282
rect 362534 84220 362540 84222
rect 362604 84220 362610 84284
rect 583520 72994 584960 73084
rect 583342 72934 584960 72994
rect 583342 72858 583402 72934
rect 583520 72858 584960 72934
rect 583342 72844 584960 72858
rect 583342 72798 583586 72844
rect 364926 71844 364932 71908
rect 364996 71906 365002 71908
rect 583526 71906 583586 72798
rect 364996 71846 583586 71906
rect 364996 71844 365002 71846
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45522 480 45612
rect -960 45462 674 45522
rect -960 45386 480 45462
rect 614 45386 674 45462
rect -960 45372 674 45386
rect 246 45326 674 45372
rect 246 44842 306 45326
rect 246 44782 6930 44842
rect 6870 44298 6930 44782
rect 362718 44298 362724 44300
rect 6870 44238 362724 44298
rect 362718 44236 362724 44238
rect 362788 44236 362794 44300
rect 580257 33146 580323 33149
rect 583520 33146 584960 33236
rect 580257 33144 584960 33146
rect 580257 33088 580262 33144
rect 580318 33088 584960 33144
rect 580257 33086 584960 33088
rect 580257 33083 580323 33086
rect 583520 32996 584960 33086
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect 322105 8938 322171 8941
rect 368657 8938 368723 8941
rect 322105 8936 368723 8938
rect 322105 8880 322110 8936
rect 322166 8880 368662 8936
rect 368718 8880 368723 8936
rect 322105 8878 368723 8880
rect 322105 8875 322171 8878
rect 368657 8875 368723 8878
rect 351637 6762 351703 6765
rect 361665 6762 361731 6765
rect 351637 6760 361731 6762
rect 351637 6704 351642 6760
rect 351698 6704 361670 6760
rect 361726 6704 361731 6760
rect 351637 6702 361731 6704
rect 351637 6699 351703 6702
rect 361665 6699 361731 6702
rect 348049 6626 348115 6629
rect 364701 6626 364767 6629
rect 348049 6624 364767 6626
rect -960 6490 480 6580
rect 348049 6568 348054 6624
rect 348110 6568 364706 6624
rect 364762 6568 364767 6624
rect 348049 6566 364767 6568
rect 348049 6563 348115 6566
rect 364701 6563 364767 6566
rect 346945 6490 347011 6493
rect 364793 6490 364859 6493
rect -960 6430 674 6490
rect -960 6354 480 6430
rect 614 6354 674 6430
rect 346945 6488 364859 6490
rect 346945 6432 346950 6488
rect 347006 6432 364798 6488
rect 364854 6432 364859 6488
rect 583520 6476 584960 6716
rect 346945 6430 364859 6432
rect 346945 6427 347011 6430
rect 364793 6427 364859 6430
rect -960 6340 674 6354
rect 246 6294 674 6340
rect 344553 6354 344619 6357
rect 366173 6354 366239 6357
rect 344553 6352 366239 6354
rect 344553 6296 344558 6352
rect 344614 6296 366178 6352
rect 366234 6296 366239 6352
rect 344553 6294 366239 6296
rect 246 5810 306 6294
rect 344553 6291 344619 6294
rect 366173 6291 366239 6294
rect 320909 6218 320975 6221
rect 367318 6218 367324 6220
rect 320909 6216 367324 6218
rect 320909 6160 320914 6216
rect 320970 6160 367324 6216
rect 320909 6158 367324 6160
rect 320909 6155 320975 6158
rect 367318 6156 367324 6158
rect 367388 6156 367394 6220
rect 246 5750 6930 5810
rect 6870 5674 6930 5750
rect 362902 5674 362908 5676
rect 6870 5614 362908 5674
rect 362902 5612 362908 5614
rect 362972 5612 362978 5676
rect 342161 4042 342227 4045
rect 360142 4042 360148 4044
rect 342161 4040 360148 4042
rect 342161 3984 342166 4040
rect 342222 3984 360148 4040
rect 342161 3982 360148 3984
rect 342161 3979 342227 3982
rect 360142 3980 360148 3982
rect 360212 3980 360218 4044
rect 215150 3844 215156 3908
rect 215220 3906 215226 3908
rect 222745 3906 222811 3909
rect 215220 3904 222811 3906
rect 215220 3848 222750 3904
rect 222806 3848 222811 3904
rect 215220 3846 222811 3848
rect 215220 3844 215226 3846
rect 222745 3843 222811 3846
rect 338665 3906 338731 3909
rect 358854 3906 358860 3908
rect 338665 3904 358860 3906
rect 338665 3848 338670 3904
rect 338726 3848 358860 3904
rect 338665 3846 358860 3848
rect 338665 3843 338731 3846
rect 358854 3844 358860 3846
rect 358924 3844 358930 3908
rect 365110 3844 365116 3908
rect 365180 3906 365186 3908
rect 365180 3846 374010 3906
rect 365180 3844 365186 3846
rect 216438 3708 216444 3772
rect 216508 3770 216514 3772
rect 227529 3770 227595 3773
rect 216508 3768 227595 3770
rect 216508 3712 227534 3768
rect 227590 3712 227595 3768
rect 216508 3710 227595 3712
rect 216508 3708 216514 3710
rect 227529 3707 227595 3710
rect 335077 3770 335143 3773
rect 360510 3770 360516 3772
rect 335077 3768 360516 3770
rect 335077 3712 335082 3768
rect 335138 3712 360516 3768
rect 335077 3710 360516 3712
rect 335077 3707 335143 3710
rect 360510 3708 360516 3710
rect 360580 3708 360586 3772
rect 367686 3708 367692 3772
rect 367756 3770 367762 3772
rect 373950 3770 374010 3846
rect 394233 3770 394299 3773
rect 367756 3710 371066 3770
rect 373950 3768 394299 3770
rect 373950 3712 394238 3768
rect 394294 3712 394299 3768
rect 373950 3710 394299 3712
rect 367756 3708 367762 3710
rect 218053 3634 218119 3637
rect 219198 3634 219204 3636
rect 218053 3632 219204 3634
rect 218053 3576 218058 3632
rect 218114 3576 219204 3632
rect 218053 3574 219204 3576
rect 218053 3571 218119 3574
rect 219198 3572 219204 3574
rect 219268 3572 219274 3636
rect 219341 3634 219407 3637
rect 331581 3634 331647 3637
rect 359406 3634 359412 3636
rect 219341 3632 219450 3634
rect 219341 3576 219346 3632
rect 219402 3576 219450 3632
rect 219341 3571 219450 3576
rect 331581 3632 359412 3634
rect 331581 3576 331586 3632
rect 331642 3576 359412 3632
rect 331581 3574 359412 3576
rect 331581 3571 331647 3574
rect 359406 3572 359412 3574
rect 359476 3572 359482 3636
rect 368974 3572 368980 3636
rect 369044 3634 369050 3636
rect 371006 3634 371066 3710
rect 394233 3707 394299 3710
rect 397729 3634 397795 3637
rect 369044 3574 370882 3634
rect 371006 3632 397795 3634
rect 371006 3576 397734 3632
rect 397790 3576 397795 3632
rect 371006 3574 397795 3576
rect 369044 3572 369050 3574
rect 213126 3436 213132 3500
rect 213196 3498 213202 3500
rect 213361 3498 213427 3501
rect 213196 3496 213427 3498
rect 213196 3440 213366 3496
rect 213422 3440 213427 3496
rect 213196 3438 213427 3440
rect 213196 3436 213202 3438
rect 213361 3435 213427 3438
rect 214465 3498 214531 3501
rect 214966 3498 214972 3500
rect 214465 3496 214972 3498
rect 214465 3440 214470 3496
rect 214526 3440 214972 3496
rect 214465 3438 214972 3440
rect 214465 3435 214531 3438
rect 214966 3436 214972 3438
rect 215036 3436 215042 3500
rect 215661 3498 215727 3501
rect 216254 3498 216260 3500
rect 215661 3496 216260 3498
rect 215661 3440 215666 3496
rect 215722 3440 216260 3496
rect 215661 3438 216260 3440
rect 215661 3435 215727 3438
rect 216254 3436 216260 3438
rect 216324 3436 216330 3500
rect 216857 3498 216923 3501
rect 218646 3498 218652 3500
rect 216857 3496 218652 3498
rect 216857 3440 216862 3496
rect 216918 3440 218652 3496
rect 216857 3438 218652 3440
rect 216857 3435 216923 3438
rect 218646 3436 218652 3438
rect 218716 3436 218722 3500
rect 219014 3436 219020 3500
rect 219084 3498 219090 3500
rect 219249 3498 219315 3501
rect 219084 3496 219315 3498
rect 219084 3440 219254 3496
rect 219310 3440 219315 3496
rect 219084 3438 219315 3440
rect 219390 3498 219450 3571
rect 237005 3498 237071 3501
rect 219390 3496 237071 3498
rect 219390 3440 237010 3496
rect 237066 3440 237071 3496
rect 219390 3438 237071 3440
rect 219084 3436 219090 3438
rect 219249 3435 219315 3438
rect 237005 3435 237071 3438
rect 325601 3498 325667 3501
rect 358118 3498 358124 3500
rect 325601 3496 358124 3498
rect 325601 3440 325606 3496
rect 325662 3440 358124 3496
rect 325601 3438 358124 3440
rect 325601 3435 325667 3438
rect 358118 3436 358124 3438
rect 358188 3436 358194 3500
rect 358302 3436 358308 3500
rect 358372 3498 358378 3500
rect 358721 3498 358787 3501
rect 358372 3496 358787 3498
rect 358372 3440 358726 3496
rect 358782 3440 358787 3496
rect 358372 3438 358787 3440
rect 358372 3436 358378 3438
rect 358721 3435 358787 3438
rect 359038 3436 359044 3500
rect 359108 3498 359114 3500
rect 359917 3498 359983 3501
rect 359108 3496 359983 3498
rect 359108 3440 359922 3496
rect 359978 3440 359983 3496
rect 359108 3438 359983 3440
rect 359108 3436 359114 3438
rect 359917 3435 359983 3438
rect 360326 3436 360332 3500
rect 360396 3498 360402 3500
rect 361113 3498 361179 3501
rect 360396 3496 361179 3498
rect 360396 3440 361118 3496
rect 361174 3440 361179 3496
rect 360396 3438 361179 3440
rect 360396 3436 360402 3438
rect 361113 3435 361179 3438
rect 363086 3436 363092 3500
rect 363156 3498 363162 3500
rect 363505 3498 363571 3501
rect 363156 3496 363571 3498
rect 363156 3440 363510 3496
rect 363566 3440 363571 3496
rect 363156 3438 363571 3440
rect 363156 3436 363162 3438
rect 363505 3435 363571 3438
rect 364374 3436 364380 3500
rect 364444 3498 364450 3500
rect 364609 3498 364675 3501
rect 364444 3496 364675 3498
rect 364444 3440 364614 3496
rect 364670 3440 364675 3496
rect 364444 3438 364675 3440
rect 364444 3436 364450 3438
rect 364609 3435 364675 3438
rect 365662 3436 365668 3500
rect 365732 3498 365738 3500
rect 365805 3498 365871 3501
rect 365732 3496 365871 3498
rect 365732 3440 365810 3496
rect 365866 3440 365871 3496
rect 365732 3438 365871 3440
rect 365732 3436 365738 3438
rect 365805 3435 365871 3438
rect 367134 3436 367140 3500
rect 367204 3498 367210 3500
rect 368197 3498 368263 3501
rect 367204 3496 368263 3498
rect 367204 3440 368202 3496
rect 368258 3440 368263 3496
rect 367204 3438 368263 3440
rect 367204 3436 367210 3438
rect 368197 3435 368263 3438
rect 368422 3436 368428 3500
rect 368492 3498 368498 3500
rect 369393 3498 369459 3501
rect 368492 3496 369459 3498
rect 368492 3440 369398 3496
rect 369454 3440 369459 3496
rect 368492 3438 369459 3440
rect 368492 3436 368498 3438
rect 369393 3435 369459 3438
rect 369894 3436 369900 3500
rect 369964 3498 369970 3500
rect 370589 3498 370655 3501
rect 369964 3496 370655 3498
rect 369964 3440 370594 3496
rect 370650 3440 370655 3496
rect 369964 3438 370655 3440
rect 370822 3498 370882 3574
rect 397729 3571 397795 3574
rect 411897 3498 411963 3501
rect 370822 3496 411963 3498
rect 370822 3440 411902 3496
rect 411958 3440 411963 3496
rect 370822 3438 411963 3440
rect 369964 3436 369970 3438
rect 370589 3435 370655 3438
rect 411897 3435 411963 3438
rect 200297 3362 200363 3365
rect 215886 3362 215892 3364
rect 200297 3360 215892 3362
rect 200297 3304 200302 3360
rect 200358 3304 215892 3360
rect 200297 3302 215892 3304
rect 200297 3299 200363 3302
rect 215886 3300 215892 3302
rect 215956 3300 215962 3364
rect 217542 3300 217548 3364
rect 217612 3362 217618 3364
rect 324405 3362 324471 3365
rect 358486 3362 358492 3364
rect 217612 3302 238770 3362
rect 217612 3300 217618 3302
rect 215109 3226 215175 3229
rect 226333 3226 226399 3229
rect 215109 3224 226399 3226
rect 215109 3168 215114 3224
rect 215170 3168 226338 3224
rect 226394 3168 226399 3224
rect 215109 3166 226399 3168
rect 238710 3226 238770 3302
rect 324405 3360 358492 3362
rect 324405 3304 324410 3360
rect 324466 3304 358492 3360
rect 324405 3302 358492 3304
rect 324405 3299 324471 3302
rect 358486 3300 358492 3302
rect 358556 3300 358562 3364
rect 363454 3300 363460 3364
rect 363524 3362 363530 3364
rect 501781 3362 501847 3365
rect 363524 3360 501847 3362
rect 363524 3304 501786 3360
rect 501842 3304 501847 3360
rect 363524 3302 501847 3304
rect 363524 3300 363530 3302
rect 501781 3299 501847 3302
rect 251173 3226 251239 3229
rect 238710 3224 251239 3226
rect 238710 3168 251178 3224
rect 251234 3168 251239 3224
rect 238710 3166 251239 3168
rect 215109 3163 215175 3166
rect 226333 3163 226399 3166
rect 251173 3163 251239 3166
rect 345749 3226 345815 3229
rect 359222 3226 359228 3228
rect 345749 3224 359228 3226
rect 345749 3168 345754 3224
rect 345810 3168 359228 3224
rect 345749 3166 359228 3168
rect 345749 3163 345815 3166
rect 359222 3164 359228 3166
rect 359292 3164 359298 3228
rect 216581 3090 216647 3093
rect 219341 3090 219407 3093
rect 216581 3088 219407 3090
rect 216581 3032 216586 3088
rect 216642 3032 219346 3088
rect 219402 3032 219407 3088
rect 216581 3030 219407 3032
rect 216581 3027 216647 3030
rect 219341 3027 219407 3030
<< via3 >>
rect 265940 477260 266004 477324
rect 268332 477260 268396 477324
rect 256188 477124 256252 477188
rect 280844 476988 280908 477052
rect 305868 476988 305932 477052
rect 308444 476988 308508 477052
rect 258028 476852 258092 476916
rect 278452 476852 278516 476916
rect 311020 476852 311084 476916
rect 253612 476716 253676 476780
rect 270908 476716 270972 476780
rect 276980 476716 277044 476780
rect 303476 476716 303540 476780
rect 323348 476716 323412 476780
rect 244228 476640 244292 476644
rect 244228 476584 244278 476640
rect 244278 476584 244292 476640
rect 244228 476580 244292 476584
rect 248276 476580 248340 476644
rect 250668 476580 250732 476644
rect 258396 476580 258460 476644
rect 263548 476640 263612 476644
rect 263548 476584 263598 476640
rect 263598 476584 263612 476640
rect 263548 476580 263612 476584
rect 260972 476444 261036 476508
rect 273484 476444 273548 476508
rect 313412 476444 313476 476508
rect 315804 476444 315868 476508
rect 238156 476308 238220 476372
rect 243124 476308 243188 476372
rect 245332 476308 245396 476372
rect 252324 476368 252388 476372
rect 252324 476312 252374 476368
rect 252374 476312 252388 476368
rect 252324 476308 252388 476312
rect 260788 476308 260852 476372
rect 262812 476308 262876 476372
rect 266492 476308 266556 476372
rect 273300 476308 273364 476372
rect 276060 476368 276124 476372
rect 276060 476312 276074 476368
rect 276074 476312 276124 476368
rect 276060 476308 276124 476312
rect 318380 476308 318444 476372
rect 320956 476308 321020 476372
rect 235948 476232 236012 476236
rect 235948 476176 235962 476232
rect 235962 476176 236012 476232
rect 235948 476172 236012 476176
rect 237236 476172 237300 476236
rect 239628 476172 239692 476236
rect 240548 476172 240612 476236
rect 241836 476172 241900 476236
rect 246436 476172 246500 476236
rect 247540 476172 247604 476236
rect 248644 476172 248708 476236
rect 250116 476172 250180 476236
rect 251404 476172 251468 476236
rect 253428 476172 253492 476236
rect 254532 476172 254596 476236
rect 255820 476172 255884 476236
rect 257108 476172 257172 476236
rect 259500 476172 259564 476236
rect 261708 476172 261772 476236
rect 263916 476172 263980 476236
rect 265388 476172 265452 476236
rect 267596 476232 267660 476236
rect 267596 476176 267646 476232
rect 267646 476176 267660 476232
rect 267596 476172 267660 476176
rect 268700 476172 268764 476236
rect 269804 476172 269868 476236
rect 271276 476172 271340 476236
rect 272196 476172 272260 476236
rect 274404 476172 274468 476236
rect 275876 476172 275940 476236
rect 278084 476172 278148 476236
rect 279188 476172 279252 476236
rect 283420 476172 283484 476236
rect 285996 476172 286060 476236
rect 288204 476172 288268 476236
rect 290964 476172 291028 476236
rect 293356 476172 293420 476236
rect 295932 476172 295996 476236
rect 298508 476172 298572 476236
rect 300900 476232 300964 476236
rect 300900 476176 300914 476232
rect 300914 476176 300964 476232
rect 300900 476172 300964 476176
rect 325924 476172 325988 476236
rect 369164 445980 369228 446044
rect 364932 444620 364996 444684
rect 214420 444348 214484 444412
rect 362540 443396 362604 443460
rect 362724 443456 362788 443460
rect 362724 443400 362774 443456
rect 362774 443400 362788 443456
rect 362724 443396 362788 443400
rect 362908 443396 362972 443460
rect 216996 308892 217060 308956
rect 217180 308756 217244 308820
rect 217364 308620 217428 308684
rect 358860 308484 358924 308548
rect 360332 308348 360396 308412
rect 218652 306988 218716 307052
rect 368980 306988 369044 307052
rect 219204 306172 219268 306236
rect 216076 306036 216140 306100
rect 215156 305900 215220 305964
rect 214788 305764 214852 305828
rect 217548 305628 217612 305692
rect 365116 304268 365180 304332
rect 367692 304132 367756 304196
rect 216444 303316 216508 303380
rect 212948 303180 213012 303244
rect 365668 298692 365732 298756
rect 367140 286316 367204 286380
rect 360332 284820 360396 284884
rect 216260 275164 216324 275228
rect 369900 269724 369964 269788
rect 363092 267004 363156 267068
rect 214972 265508 215036 265572
rect 215892 262788 215956 262852
rect 363460 262788 363524 262852
rect 359044 260068 359108 260132
rect 368428 254492 368492 254556
rect 360700 250684 360764 250748
rect 213132 249052 213196 249116
rect 364380 249052 364444 249116
rect 358124 248100 358188 248164
rect 219020 246196 219084 246260
rect 358308 245516 358372 245580
rect 359228 245380 359292 245444
rect 359412 245244 359476 245308
rect 357940 245108 358004 245172
rect 358492 244972 358556 245036
rect 360516 244836 360580 244900
rect 367324 244700 367388 244764
rect 363276 244564 363340 244628
rect 218100 243340 218164 243404
rect 369164 177244 369228 177308
rect 218100 162828 218164 162892
rect 273318 159896 273382 159900
rect 273318 159840 273350 159896
rect 273350 159840 273382 159896
rect 273318 159836 273382 159840
rect 278078 159896 278142 159900
rect 278078 159840 278134 159896
rect 278134 159840 278142 159896
rect 278078 159836 278142 159840
rect 261078 159760 261142 159764
rect 261078 159704 261114 159760
rect 261114 159704 261142 159760
rect 261078 159700 261142 159704
rect 260670 159564 260734 159628
rect 275766 159564 275830 159628
rect 276990 159624 277054 159628
rect 276990 159568 277030 159624
rect 277030 159568 277054 159624
rect 276990 159564 277054 159568
rect 279166 159564 279230 159628
rect 357940 159292 358004 159356
rect 360700 159292 360764 159356
rect 363276 159292 363340 159356
rect 259500 159156 259564 159220
rect 254532 159020 254596 159084
rect 253612 158884 253676 158948
rect 243124 158748 243188 158812
rect 216996 158612 217060 158676
rect 238156 158672 238220 158676
rect 238156 158616 238170 158672
rect 238170 158616 238220 158672
rect 238156 158612 238220 158616
rect 239628 158672 239692 158676
rect 239628 158616 239642 158672
rect 239642 158616 239692 158672
rect 239628 158612 239692 158616
rect 241836 158612 241900 158676
rect 244228 158612 244292 158676
rect 245516 158672 245580 158676
rect 245516 158616 245566 158672
rect 245566 158616 245580 158672
rect 245516 158612 245580 158616
rect 248276 158672 248340 158676
rect 248276 158616 248326 158672
rect 248326 158616 248340 158672
rect 248276 158612 248340 158616
rect 252324 158672 252388 158676
rect 252324 158616 252374 158672
rect 252374 158616 252388 158672
rect 252324 158612 252388 158616
rect 255820 158672 255884 158676
rect 255820 158616 255870 158672
rect 255870 158616 255884 158672
rect 255820 158612 255884 158616
rect 257108 158612 257172 158676
rect 261708 158672 261772 158676
rect 261708 158616 261758 158672
rect 261758 158616 261772 158672
rect 261708 158612 261772 158616
rect 265388 158672 265452 158676
rect 265388 158616 265438 158672
rect 265438 158616 265452 158672
rect 265388 158612 265452 158616
rect 265940 158672 266004 158676
rect 265940 158616 265990 158672
rect 265990 158616 266004 158672
rect 265940 158612 266004 158616
rect 266492 158672 266556 158676
rect 266492 158616 266542 158672
rect 266542 158616 266556 158672
rect 266492 158612 266556 158616
rect 268700 158672 268764 158676
rect 268700 158616 268750 158672
rect 268750 158616 268764 158672
rect 268700 158612 268764 158616
rect 269804 158612 269868 158676
rect 270908 158672 270972 158676
rect 270908 158616 270958 158672
rect 270958 158616 270972 158672
rect 270908 158612 270972 158616
rect 272196 158672 272260 158676
rect 272196 158616 272246 158672
rect 272246 158616 272260 158672
rect 272196 158612 272260 158616
rect 274404 158672 274468 158676
rect 274404 158616 274454 158672
rect 274454 158616 274468 158672
rect 274404 158612 274468 158616
rect 276060 158672 276124 158676
rect 276060 158616 276110 158672
rect 276110 158616 276124 158672
rect 276060 158612 276124 158616
rect 281028 158672 281092 158676
rect 281028 158616 281078 158672
rect 281078 158616 281092 158672
rect 281028 158612 281092 158616
rect 288204 158672 288268 158676
rect 288204 158616 288254 158672
rect 288254 158616 288268 158672
rect 288204 158612 288268 158616
rect 290964 158672 291028 158676
rect 290964 158616 291014 158672
rect 291014 158616 291028 158672
rect 290964 158612 291028 158616
rect 293540 158672 293604 158676
rect 293540 158616 293590 158672
rect 293590 158616 293604 158672
rect 293540 158612 293604 158616
rect 295932 158672 295996 158676
rect 295932 158616 295982 158672
rect 295982 158616 295996 158672
rect 295932 158612 295996 158616
rect 298508 158672 298572 158676
rect 298508 158616 298558 158672
rect 298558 158616 298572 158672
rect 298508 158612 298572 158616
rect 300900 158672 300964 158676
rect 300900 158616 300950 158672
rect 300950 158616 300964 158672
rect 300900 158612 300964 158616
rect 303476 158672 303540 158676
rect 303476 158616 303526 158672
rect 303526 158616 303540 158672
rect 303476 158612 303540 158616
rect 306052 158672 306116 158676
rect 306052 158616 306102 158672
rect 306102 158616 306116 158672
rect 306052 158612 306116 158616
rect 308628 158672 308692 158676
rect 308628 158616 308678 158672
rect 308678 158616 308692 158672
rect 308628 158612 308692 158616
rect 311020 158672 311084 158676
rect 311020 158616 311070 158672
rect 311070 158616 311084 158672
rect 311020 158612 311084 158616
rect 313412 158672 313476 158676
rect 313412 158616 313462 158672
rect 313462 158616 313476 158672
rect 313412 158612 313476 158616
rect 315804 158672 315868 158676
rect 315804 158616 315854 158672
rect 315854 158616 315868 158672
rect 315804 158612 315868 158616
rect 318564 158672 318628 158676
rect 318564 158616 318614 158672
rect 318614 158616 318628 158672
rect 318564 158612 318628 158616
rect 320956 158672 321020 158676
rect 320956 158616 321006 158672
rect 321006 158616 321020 158672
rect 320956 158612 321020 158616
rect 323348 158672 323412 158676
rect 323348 158616 323398 158672
rect 323398 158616 323412 158672
rect 323348 158612 323412 158616
rect 325924 158672 325988 158676
rect 325924 158616 325974 158672
rect 325974 158616 325988 158672
rect 325924 158612 325988 158616
rect 236132 158476 236196 158540
rect 216076 158340 216140 158404
rect 258212 158340 258276 158404
rect 217180 158204 217244 158268
rect 240548 158204 240612 158268
rect 258580 158204 258644 158268
rect 217364 158068 217428 158132
rect 262628 158068 262692 158132
rect 214788 157932 214852 157996
rect 246620 157992 246684 157996
rect 246620 157936 246670 157992
rect 246670 157936 246684 157992
rect 212948 157796 213012 157860
rect 246620 157932 246684 157936
rect 247724 157932 247788 157996
rect 250852 157932 250916 157996
rect 267044 157932 267108 157996
rect 248644 157856 248708 157860
rect 248644 157800 248694 157856
rect 248694 157800 248708 157856
rect 248644 157796 248708 157800
rect 250116 157796 250180 157860
rect 251404 157796 251468 157860
rect 253428 157856 253492 157860
rect 253428 157800 253478 157856
rect 253478 157800 253492 157856
rect 253428 157796 253492 157800
rect 263916 157796 263980 157860
rect 268332 157720 268396 157724
rect 268332 157664 268382 157720
rect 268382 157664 268396 157720
rect 268332 157660 268396 157664
rect 271276 157720 271340 157724
rect 271276 157664 271326 157720
rect 271326 157664 271340 157720
rect 271276 157660 271340 157664
rect 273668 157720 273732 157724
rect 273668 157664 273718 157720
rect 273718 157664 273732 157720
rect 273668 157660 273732 157664
rect 278452 157720 278516 157724
rect 278452 157664 278502 157720
rect 278502 157664 278516 157720
rect 278452 157660 278516 157664
rect 256188 157584 256252 157588
rect 256188 157528 256238 157584
rect 256238 157528 256252 157584
rect 256188 157524 256252 157528
rect 263548 157524 263612 157588
rect 283604 157584 283668 157588
rect 283604 157528 283654 157584
rect 283654 157528 283668 157584
rect 283604 157524 283668 157528
rect 285996 157584 286060 157588
rect 285996 157528 286046 157584
rect 286046 157528 286060 157584
rect 285996 157524 286060 157528
rect 237236 157388 237300 157452
rect 214420 110468 214484 110532
rect 362540 84220 362604 84284
rect 364932 71844 364996 71908
rect 362724 44236 362788 44300
rect 367324 6156 367388 6220
rect 362908 5612 362972 5676
rect 360148 3980 360212 4044
rect 215156 3844 215220 3908
rect 358860 3844 358924 3908
rect 365116 3844 365180 3908
rect 216444 3708 216508 3772
rect 360516 3708 360580 3772
rect 367692 3708 367756 3772
rect 219204 3572 219268 3636
rect 359412 3572 359476 3636
rect 368980 3572 369044 3636
rect 213132 3436 213196 3500
rect 214972 3436 215036 3500
rect 216260 3436 216324 3500
rect 218652 3436 218716 3500
rect 219020 3436 219084 3500
rect 358124 3436 358188 3500
rect 358308 3436 358372 3500
rect 359044 3436 359108 3500
rect 360332 3436 360396 3500
rect 363092 3436 363156 3500
rect 364380 3436 364444 3500
rect 365668 3436 365732 3500
rect 367140 3436 367204 3500
rect 368428 3436 368492 3500
rect 369900 3436 369964 3500
rect 215892 3300 215956 3364
rect 217548 3300 217612 3364
rect 358492 3300 358556 3364
rect 363460 3300 363524 3364
rect 359228 3164 359292 3228
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 60294 205954 60914 241398
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 214954 69914 250398
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 223954 78914 259398
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 228454 83414 263898
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 232954 87914 268398
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 241954 96914 277398
rect 96294 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 96914 241954
rect 96294 241634 96914 241718
rect 96294 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 96914 241634
rect 96294 205954 96914 241398
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 246454 101414 281898
rect 100794 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 101414 246454
rect 100794 246134 101414 246218
rect 100794 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 101414 246134
rect 100794 210454 101414 245898
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 100794 174454 101414 209898
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 138454 101414 173898
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 214954 105914 250398
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 105294 142954 105914 178398
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 259954 114914 295398
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 223954 114914 259398
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 151954 114914 187398
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114294 115954 114914 151398
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118794 228454 119414 263898
rect 118794 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 119414 228454
rect 118794 228134 119414 228218
rect 118794 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 119414 228134
rect 118794 192454 119414 227898
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 120454 119414 155898
rect 118794 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 119414 120454
rect 118794 120134 119414 120218
rect 118794 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 119414 120134
rect 118794 84454 119414 119898
rect 118794 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 119414 84454
rect 118794 84134 119414 84218
rect 118794 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 119414 84134
rect 118794 48454 119414 83898
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 232954 123914 268398
rect 123294 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 123914 232954
rect 123294 232634 123914 232718
rect 123294 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 123914 232634
rect 123294 196954 123914 232398
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 123294 124954 123914 160398
rect 123294 124718 123326 124954
rect 123562 124718 123646 124954
rect 123882 124718 123914 124954
rect 123294 124634 123914 124718
rect 123294 124398 123326 124634
rect 123562 124398 123646 124634
rect 123882 124398 123914 124634
rect 123294 88954 123914 124398
rect 123294 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 123914 88954
rect 123294 88634 123914 88718
rect 123294 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 123914 88634
rect 123294 52954 123914 88398
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 241954 132914 277398
rect 132294 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 132914 241954
rect 132294 241634 132914 241718
rect 132294 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 132914 241634
rect 132294 205954 132914 241398
rect 132294 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 132914 205954
rect 132294 205634 132914 205718
rect 132294 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 132914 205634
rect 132294 169954 132914 205398
rect 132294 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 132914 169954
rect 132294 169634 132914 169718
rect 132294 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 132914 169634
rect 132294 133954 132914 169398
rect 132294 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 132914 133954
rect 132294 133634 132914 133718
rect 132294 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 132914 133634
rect 132294 97954 132914 133398
rect 132294 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 132914 97954
rect 132294 97634 132914 97718
rect 132294 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 132914 97634
rect 132294 61954 132914 97398
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 246454 137414 281898
rect 136794 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 137414 246454
rect 136794 246134 137414 246218
rect 136794 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 137414 246134
rect 136794 210454 137414 245898
rect 136794 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 137414 210454
rect 136794 210134 137414 210218
rect 136794 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 137414 210134
rect 136794 174454 137414 209898
rect 136794 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 137414 174454
rect 136794 174134 137414 174218
rect 136794 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 137414 174134
rect 136794 138454 137414 173898
rect 136794 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 137414 138454
rect 136794 138134 137414 138218
rect 136794 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 137414 138134
rect 136794 102454 137414 137898
rect 136794 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 137414 102454
rect 136794 102134 137414 102218
rect 136794 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 137414 102134
rect 136794 66454 137414 101898
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6106 137414 29898
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 214954 141914 250398
rect 141294 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 141914 214954
rect 141294 214634 141914 214718
rect 141294 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 141914 214634
rect 141294 178954 141914 214398
rect 141294 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 141914 178954
rect 141294 178634 141914 178718
rect 141294 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 141914 178634
rect 141294 142954 141914 178398
rect 141294 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 141914 142954
rect 141294 142634 141914 142718
rect 141294 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 141914 142634
rect 141294 106954 141914 142398
rect 141294 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 141914 106954
rect 141294 106634 141914 106718
rect 141294 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 141914 106634
rect 141294 70954 141914 106398
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7066 141914 34398
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 223954 150914 259398
rect 150294 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 150914 223954
rect 150294 223634 150914 223718
rect 150294 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 150914 223634
rect 150294 187954 150914 223398
rect 150294 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 150914 187954
rect 150294 187634 150914 187718
rect 150294 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 150914 187634
rect 150294 151954 150914 187398
rect 150294 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 150914 151954
rect 150294 151634 150914 151718
rect 150294 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 150914 151634
rect 150294 115954 150914 151398
rect 150294 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 150914 115954
rect 150294 115634 150914 115718
rect 150294 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 150914 115634
rect 150294 79954 150914 115398
rect 150294 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 150914 79954
rect 150294 79634 150914 79718
rect 150294 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 150914 79634
rect 150294 43954 150914 79398
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 228454 155414 263898
rect 154794 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 155414 228454
rect 154794 228134 155414 228218
rect 154794 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 155414 228134
rect 154794 192454 155414 227898
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 154794 156454 155414 191898
rect 154794 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 155414 156454
rect 154794 156134 155414 156218
rect 154794 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 155414 156134
rect 154794 120454 155414 155898
rect 154794 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 155414 120454
rect 154794 120134 155414 120218
rect 154794 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 155414 120134
rect 154794 84454 155414 119898
rect 154794 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 155414 84454
rect 154794 84134 155414 84218
rect 154794 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 155414 84134
rect 154794 48454 155414 83898
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 232954 159914 268398
rect 159294 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 159914 232954
rect 159294 232634 159914 232718
rect 159294 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 159914 232634
rect 159294 196954 159914 232398
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 159294 160954 159914 196398
rect 159294 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 159914 160954
rect 159294 160634 159914 160718
rect 159294 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 159914 160634
rect 159294 124954 159914 160398
rect 159294 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 159914 124954
rect 159294 124634 159914 124718
rect 159294 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 159914 124634
rect 159294 88954 159914 124398
rect 159294 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 159914 88954
rect 159294 88634 159914 88718
rect 159294 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 159914 88634
rect 159294 52954 159914 88398
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 241954 168914 277398
rect 168294 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 168914 241954
rect 168294 241634 168914 241718
rect 168294 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 168914 241634
rect 168294 205954 168914 241398
rect 168294 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 168914 205954
rect 168294 205634 168914 205718
rect 168294 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 168914 205634
rect 168294 169954 168914 205398
rect 168294 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 168914 169954
rect 168294 169634 168914 169718
rect 168294 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 168914 169634
rect 168294 133954 168914 169398
rect 168294 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 168914 133954
rect 168294 133634 168914 133718
rect 168294 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 168914 133634
rect 168294 97954 168914 133398
rect 168294 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 168914 97954
rect 168294 97634 168914 97718
rect 168294 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 168914 97634
rect 168294 61954 168914 97398
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 246454 173414 281898
rect 172794 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 173414 246454
rect 172794 246134 173414 246218
rect 172794 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 173414 246134
rect 172794 210454 173414 245898
rect 172794 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 173414 210454
rect 172794 210134 173414 210218
rect 172794 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 173414 210134
rect 172794 174454 173414 209898
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 172794 138454 173414 173898
rect 172794 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 173414 138454
rect 172794 138134 173414 138218
rect 172794 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 173414 138134
rect 172794 102454 173414 137898
rect 172794 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 173414 102454
rect 172794 102134 173414 102218
rect 172794 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 173414 102134
rect 172794 66454 173414 101898
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 214954 177914 250398
rect 177294 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 177914 214954
rect 177294 214634 177914 214718
rect 177294 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 177914 214634
rect 177294 178954 177914 214398
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 106954 177914 142398
rect 177294 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 177914 106954
rect 177294 106634 177914 106718
rect 177294 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 177914 106634
rect 177294 70954 177914 106398
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 259954 186914 295398
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 223954 186914 259398
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 187954 186914 223398
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 115954 186914 151398
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 186294 79954 186914 115398
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 186294 79634 186914 79718
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 228454 191414 263898
rect 190794 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 191414 228454
rect 190794 228134 191414 228218
rect 190794 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 191414 228134
rect 190794 192454 191414 227898
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 120454 191414 155898
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 84454 191414 119898
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 195294 232954 195914 268398
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 196954 195914 232398
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 241954 204914 277398
rect 204294 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 204914 241954
rect 204294 241634 204914 241718
rect 204294 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 204914 241634
rect 204294 205954 204914 241398
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 565308 218414 578898
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 565308 222914 583398
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 565308 227414 587898
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 565308 231914 592398
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 565308 236414 596898
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 565308 240914 565398
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 565308 245414 569898
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 565308 249914 574398
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 565308 254414 578898
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 565308 258914 583398
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 565308 263414 587898
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 565308 267914 592398
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 565308 272414 596898
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 565308 276914 565398
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 565308 281414 569898
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 565308 285914 574398
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 565308 290414 578898
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 565308 294914 583398
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 565308 299414 587898
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 565308 303914 592398
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 565308 308414 596898
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 565308 312914 565398
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 565308 317414 569898
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 565308 321914 574398
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 565308 326414 578898
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 565308 330914 583398
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 565308 335414 587898
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 565308 339914 592398
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 565308 344414 596898
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 565308 348914 565398
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 565308 353414 569898
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 565308 357914 574398
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 220272 547954 220620 547986
rect 220272 547718 220328 547954
rect 220564 547718 220620 547954
rect 220272 547634 220620 547718
rect 220272 547398 220328 547634
rect 220564 547398 220620 547634
rect 220272 547366 220620 547398
rect 356000 547954 356348 547986
rect 356000 547718 356056 547954
rect 356292 547718 356348 547954
rect 356000 547634 356348 547718
rect 356000 547398 356056 547634
rect 356292 547398 356348 547634
rect 356000 547366 356348 547398
rect 220952 543454 221300 543486
rect 220952 543218 221008 543454
rect 221244 543218 221300 543454
rect 220952 543134 221300 543218
rect 220952 542898 221008 543134
rect 221244 542898 221300 543134
rect 220952 542866 221300 542898
rect 355320 543454 355668 543486
rect 355320 543218 355376 543454
rect 355612 543218 355668 543454
rect 355320 543134 355668 543218
rect 355320 542898 355376 543134
rect 355612 542898 355668 543134
rect 355320 542866 355668 542898
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 220272 511954 220620 511986
rect 220272 511718 220328 511954
rect 220564 511718 220620 511954
rect 220272 511634 220620 511718
rect 220272 511398 220328 511634
rect 220564 511398 220620 511634
rect 220272 511366 220620 511398
rect 356000 511954 356348 511986
rect 356000 511718 356056 511954
rect 356292 511718 356348 511954
rect 356000 511634 356348 511718
rect 356000 511398 356056 511634
rect 356292 511398 356348 511634
rect 356000 511366 356348 511398
rect 220952 507454 221300 507486
rect 220952 507218 221008 507454
rect 221244 507218 221300 507454
rect 220952 507134 221300 507218
rect 220952 506898 221008 507134
rect 221244 506898 221300 507134
rect 220952 506866 221300 506898
rect 355320 507454 355668 507486
rect 355320 507218 355376 507454
rect 355612 507218 355668 507454
rect 355320 507134 355668 507218
rect 355320 506898 355376 507134
rect 355612 506898 355668 507134
rect 355320 506866 355668 506898
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 236056 479770 236116 480080
rect 235950 479710 236116 479770
rect 237144 479770 237204 480080
rect 238232 479770 238292 480080
rect 237144 479710 237298 479770
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 217794 471454 218414 478000
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 214419 444412 214485 444413
rect 214419 444348 214420 444412
rect 214484 444348 214485 444412
rect 214419 444347 214485 444348
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 212947 303244 213013 303245
rect 212947 303180 212948 303244
rect 213012 303180 213013 303244
rect 212947 303179 213013 303180
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 246454 209414 281898
rect 208794 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 209414 246454
rect 208794 246134 209414 246218
rect 208794 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 209414 246134
rect 208794 210454 209414 245898
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 212950 157861 213010 303179
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213131 249116 213197 249117
rect 213131 249052 213132 249116
rect 213196 249052 213197 249116
rect 213131 249051 213197 249052
rect 212947 157860 213013 157861
rect 212947 157796 212948 157860
rect 213012 157796 213013 157860
rect 212947 157795 213013 157796
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 213134 3501 213194 249051
rect 213294 214954 213914 250398
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 214422 110533 214482 444347
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 216995 308956 217061 308957
rect 216995 308892 216996 308956
rect 217060 308892 217061 308956
rect 216995 308891 217061 308892
rect 216075 306100 216141 306101
rect 216075 306036 216076 306100
rect 216140 306036 216141 306100
rect 216075 306035 216141 306036
rect 215155 305964 215221 305965
rect 215155 305900 215156 305964
rect 215220 305900 215221 305964
rect 215155 305899 215221 305900
rect 214787 305828 214853 305829
rect 214787 305764 214788 305828
rect 214852 305764 214853 305828
rect 214787 305763 214853 305764
rect 214790 157997 214850 305763
rect 214971 265572 215037 265573
rect 214971 265508 214972 265572
rect 215036 265508 215037 265572
rect 214971 265507 215037 265508
rect 214787 157996 214853 157997
rect 214787 157932 214788 157996
rect 214852 157932 214853 157996
rect 214787 157931 214853 157932
rect 214419 110532 214485 110533
rect 214419 110468 214420 110532
rect 214484 110468 214485 110532
rect 214419 110467 214485 110468
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213131 3500 213197 3501
rect 213131 3436 213132 3500
rect 213196 3436 213197 3500
rect 213131 3435 213197 3436
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 -7066 213914 34398
rect 214974 3501 215034 265507
rect 215158 3909 215218 305899
rect 215891 262852 215957 262853
rect 215891 262788 215892 262852
rect 215956 262788 215957 262852
rect 215891 262787 215957 262788
rect 215155 3908 215221 3909
rect 215155 3844 215156 3908
rect 215220 3844 215221 3908
rect 215155 3843 215221 3844
rect 214971 3500 215037 3501
rect 214971 3436 214972 3500
rect 215036 3436 215037 3500
rect 214971 3435 215037 3436
rect 215894 3365 215954 262787
rect 216078 158405 216138 306035
rect 216443 303380 216509 303381
rect 216443 303316 216444 303380
rect 216508 303316 216509 303380
rect 216443 303315 216509 303316
rect 216259 275228 216325 275229
rect 216259 275164 216260 275228
rect 216324 275164 216325 275228
rect 216259 275163 216325 275164
rect 216075 158404 216141 158405
rect 216075 158340 216076 158404
rect 216140 158340 216141 158404
rect 216075 158339 216141 158340
rect 216262 3501 216322 275163
rect 216446 3773 216506 303315
rect 216998 158677 217058 308891
rect 217179 308820 217245 308821
rect 217179 308756 217180 308820
rect 217244 308756 217245 308820
rect 217179 308755 217245 308756
rect 216995 158676 217061 158677
rect 216995 158612 216996 158676
rect 217060 158612 217061 158676
rect 216995 158611 217061 158612
rect 217182 158269 217242 308755
rect 217363 308684 217429 308685
rect 217363 308620 217364 308684
rect 217428 308620 217429 308684
rect 217363 308619 217429 308620
rect 217179 158268 217245 158269
rect 217179 158204 217180 158268
rect 217244 158204 217245 158268
rect 217179 158203 217245 158204
rect 217366 158133 217426 308619
rect 217547 305692 217613 305693
rect 217547 305628 217548 305692
rect 217612 305628 217613 305692
rect 217547 305627 217613 305628
rect 217363 158132 217429 158133
rect 217363 158068 217364 158132
rect 217428 158068 217429 158132
rect 217363 158067 217429 158068
rect 216443 3772 216509 3773
rect 216443 3708 216444 3772
rect 216508 3708 216509 3772
rect 216443 3707 216509 3708
rect 216259 3500 216325 3501
rect 216259 3436 216260 3500
rect 216324 3436 216325 3500
rect 216259 3435 216325 3436
rect 217550 3365 217610 305627
rect 217794 291454 218414 326898
rect 222294 475954 222914 478000
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 218651 307052 218717 307053
rect 218651 306988 218652 307052
rect 218716 306988 218717 307052
rect 218651 306987 218717 306988
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 245308 218414 254898
rect 218099 243404 218165 243405
rect 218099 243340 218100 243404
rect 218164 243340 218165 243404
rect 218099 243339 218165 243340
rect 218102 162893 218162 243339
rect 218099 162892 218165 162893
rect 218099 162828 218100 162892
rect 218164 162828 218165 162892
rect 218099 162827 218165 162828
rect 217794 147454 218414 158000
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 218654 3501 218714 306987
rect 219203 306236 219269 306237
rect 219203 306172 219204 306236
rect 219268 306172 219269 306236
rect 219203 306171 219269 306172
rect 219019 246260 219085 246261
rect 219019 246196 219020 246260
rect 219084 246196 219085 246260
rect 219019 246195 219085 246196
rect 219022 3501 219082 246195
rect 219206 3637 219266 306171
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 245308 222914 259398
rect 226794 444454 227414 478000
rect 235950 476237 236010 479710
rect 237238 476237 237298 479710
rect 238158 479710 238292 479770
rect 239592 479770 239652 480080
rect 240544 479770 240604 480080
rect 241768 479770 241828 480080
rect 243128 479770 243188 480080
rect 239592 479710 239690 479770
rect 240544 479710 240610 479770
rect 241768 479710 241898 479770
rect 238158 476373 238218 479710
rect 238155 476372 238221 476373
rect 238155 476308 238156 476372
rect 238220 476308 238221 476372
rect 238155 476307 238221 476308
rect 239630 476237 239690 479710
rect 240550 476237 240610 479710
rect 241838 476237 241898 479710
rect 243126 479710 243188 479770
rect 244216 479770 244276 480080
rect 245440 479770 245500 480080
rect 246528 479770 246588 480080
rect 247616 479770 247676 480080
rect 248296 479770 248356 480080
rect 248704 479770 248764 480080
rect 244216 479710 244290 479770
rect 243126 476373 243186 479710
rect 244230 476645 244290 479710
rect 245334 479710 245500 479770
rect 246438 479710 246588 479770
rect 247542 479710 247676 479770
rect 248278 479710 248356 479770
rect 248646 479710 248764 479770
rect 250064 479770 250124 480080
rect 250744 479770 250804 480080
rect 250064 479710 250178 479770
rect 244227 476644 244293 476645
rect 244227 476580 244228 476644
rect 244292 476580 244293 476644
rect 244227 476579 244293 476580
rect 245334 476373 245394 479710
rect 243123 476372 243189 476373
rect 243123 476308 243124 476372
rect 243188 476308 243189 476372
rect 243123 476307 243189 476308
rect 245331 476372 245397 476373
rect 245331 476308 245332 476372
rect 245396 476308 245397 476372
rect 245331 476307 245397 476308
rect 246438 476237 246498 479710
rect 247542 476237 247602 479710
rect 248278 476645 248338 479710
rect 248275 476644 248341 476645
rect 248275 476580 248276 476644
rect 248340 476580 248341 476644
rect 248275 476579 248341 476580
rect 248646 476237 248706 479710
rect 250118 476237 250178 479710
rect 250670 479710 250804 479770
rect 251288 479770 251348 480080
rect 252376 479770 252436 480080
rect 253464 479770 253524 480080
rect 251288 479710 251466 479770
rect 250670 476645 250730 479710
rect 250667 476644 250733 476645
rect 250667 476580 250668 476644
rect 250732 476580 250733 476644
rect 250667 476579 250733 476580
rect 251406 476237 251466 479710
rect 252326 479710 252436 479770
rect 253430 479710 253524 479770
rect 253600 479770 253660 480080
rect 254552 479770 254612 480080
rect 255912 479770 255972 480080
rect 253600 479710 253674 479770
rect 252326 476373 252386 479710
rect 252323 476372 252389 476373
rect 252323 476308 252324 476372
rect 252388 476308 252389 476372
rect 252323 476307 252389 476308
rect 253430 476237 253490 479710
rect 253614 476781 253674 479710
rect 254534 479710 254612 479770
rect 255822 479710 255972 479770
rect 256048 479770 256108 480080
rect 257000 479770 257060 480080
rect 258088 479770 258148 480080
rect 258496 479770 258556 480080
rect 256048 479710 256250 479770
rect 257000 479710 257170 479770
rect 253611 476780 253677 476781
rect 253611 476716 253612 476780
rect 253676 476716 253677 476780
rect 253611 476715 253677 476716
rect 254534 476237 254594 479710
rect 255822 476237 255882 479710
rect 256190 477189 256250 479710
rect 256187 477188 256253 477189
rect 256187 477124 256188 477188
rect 256252 477124 256253 477188
rect 256187 477123 256253 477124
rect 257110 476237 257170 479710
rect 257846 479710 258148 479770
rect 258398 479710 258556 479770
rect 259448 479770 259508 480080
rect 260672 479770 260732 480080
rect 261080 479770 261140 480080
rect 261760 479770 261820 480080
rect 262848 479770 262908 480080
rect 259448 479710 259562 479770
rect 260672 479710 260850 479770
rect 257846 476914 257906 479710
rect 258027 476916 258093 476917
rect 258027 476914 258028 476916
rect 257846 476854 258028 476914
rect 258027 476852 258028 476854
rect 258092 476852 258093 476916
rect 258027 476851 258093 476852
rect 258398 476645 258458 479710
rect 258395 476644 258461 476645
rect 258395 476580 258396 476644
rect 258460 476580 258461 476644
rect 258395 476579 258461 476580
rect 259502 476237 259562 479710
rect 260790 476373 260850 479710
rect 260974 479710 261140 479770
rect 261710 479710 261820 479770
rect 262814 479710 262908 479770
rect 263528 479770 263588 480080
rect 263936 479770 263996 480080
rect 263528 479710 263610 479770
rect 260974 476509 261034 479710
rect 260971 476508 261037 476509
rect 260971 476444 260972 476508
rect 261036 476444 261037 476508
rect 260971 476443 261037 476444
rect 260787 476372 260853 476373
rect 260787 476308 260788 476372
rect 260852 476308 260853 476372
rect 260787 476307 260853 476308
rect 261710 476237 261770 479710
rect 262814 476373 262874 479710
rect 263550 476645 263610 479710
rect 263918 479710 263996 479770
rect 265296 479770 265356 480080
rect 265976 479770 266036 480080
rect 265296 479710 265450 479770
rect 263547 476644 263613 476645
rect 263547 476580 263548 476644
rect 263612 476580 263613 476644
rect 263547 476579 263613 476580
rect 262811 476372 262877 476373
rect 262811 476308 262812 476372
rect 262876 476308 262877 476372
rect 262811 476307 262877 476308
rect 263918 476237 263978 479710
rect 265390 476237 265450 479710
rect 265942 479710 266036 479770
rect 266384 479770 266444 480080
rect 267608 479770 267668 480080
rect 266384 479710 266554 479770
rect 265942 477325 266002 479710
rect 265939 477324 266005 477325
rect 265939 477260 265940 477324
rect 266004 477260 266005 477324
rect 265939 477259 266005 477260
rect 266494 476373 266554 479710
rect 267598 479710 267668 479770
rect 268288 479770 268348 480080
rect 268696 479770 268756 480080
rect 269784 479770 269844 480080
rect 271008 479770 271068 480080
rect 268288 479710 268394 479770
rect 268696 479710 268762 479770
rect 269784 479710 269866 479770
rect 266491 476372 266557 476373
rect 266491 476308 266492 476372
rect 266556 476308 266557 476372
rect 266491 476307 266557 476308
rect 267598 476237 267658 479710
rect 268334 477325 268394 479710
rect 268331 477324 268397 477325
rect 268331 477260 268332 477324
rect 268396 477260 268397 477324
rect 268331 477259 268397 477260
rect 268702 476237 268762 479710
rect 269806 476237 269866 479710
rect 270910 479710 271068 479770
rect 271144 479770 271204 480080
rect 272232 479770 272292 480080
rect 273320 479770 273380 480080
rect 273592 479770 273652 480080
rect 274408 479770 274468 480080
rect 271144 479710 271338 479770
rect 270910 476781 270970 479710
rect 270907 476780 270973 476781
rect 270907 476716 270908 476780
rect 270972 476716 270973 476780
rect 270907 476715 270973 476716
rect 271278 476237 271338 479710
rect 272198 479710 272292 479770
rect 273302 479710 273380 479770
rect 273486 479710 273652 479770
rect 274406 479710 274468 479770
rect 275768 479770 275828 480080
rect 276040 479770 276100 480080
rect 276992 479770 277052 480080
rect 275768 479710 275938 479770
rect 276040 479710 276122 479770
rect 272198 476237 272258 479710
rect 273302 476373 273362 479710
rect 273486 476509 273546 479710
rect 273483 476508 273549 476509
rect 273483 476444 273484 476508
rect 273548 476444 273549 476508
rect 273483 476443 273549 476444
rect 273299 476372 273365 476373
rect 273299 476308 273300 476372
rect 273364 476308 273365 476372
rect 273299 476307 273365 476308
rect 274406 476237 274466 479710
rect 275878 476237 275938 479710
rect 276062 476373 276122 479710
rect 276982 479710 277052 479770
rect 278080 479770 278140 480080
rect 278488 479770 278548 480080
rect 278080 479710 278146 479770
rect 276982 476781 277042 479710
rect 276979 476780 277045 476781
rect 276979 476716 276980 476780
rect 277044 476716 277045 476780
rect 276979 476715 277045 476716
rect 276059 476372 276125 476373
rect 276059 476308 276060 476372
rect 276124 476308 276125 476372
rect 276059 476307 276125 476308
rect 278086 476237 278146 479710
rect 278454 479710 278548 479770
rect 279168 479770 279228 480080
rect 280936 479770 280996 480080
rect 283520 479770 283580 480080
rect 279168 479710 279250 479770
rect 278454 476917 278514 479710
rect 278451 476916 278517 476917
rect 278451 476852 278452 476916
rect 278516 476852 278517 476916
rect 278451 476851 278517 476852
rect 279190 476237 279250 479710
rect 280846 479710 280996 479770
rect 283422 479710 283580 479770
rect 285968 479770 286028 480080
rect 288280 479770 288340 480080
rect 291000 479770 291060 480080
rect 293448 479770 293508 480080
rect 285968 479710 286058 479770
rect 280846 477053 280906 479710
rect 280843 477052 280909 477053
rect 280843 476988 280844 477052
rect 280908 476988 280909 477052
rect 280843 476987 280909 476988
rect 283422 476237 283482 479710
rect 285998 476237 286058 479710
rect 288206 479710 288340 479770
rect 290966 479710 291060 479770
rect 293358 479710 293508 479770
rect 295896 479770 295956 480080
rect 298480 479770 298540 480080
rect 300928 479770 300988 480080
rect 303512 479770 303572 480080
rect 305960 479770 306020 480080
rect 308544 479770 308604 480080
rect 295896 479710 295994 479770
rect 298480 479710 298570 479770
rect 288206 476237 288266 479710
rect 290966 476237 291026 479710
rect 293358 476237 293418 479710
rect 295934 476237 295994 479710
rect 298510 476237 298570 479710
rect 300902 479710 300988 479770
rect 303478 479710 303572 479770
rect 305870 479710 306020 479770
rect 308446 479710 308604 479770
rect 310992 479770 311052 480080
rect 313440 479770 313500 480080
rect 315888 479770 315948 480080
rect 318472 479770 318532 480080
rect 310992 479710 311082 479770
rect 300902 476237 300962 479710
rect 303478 476781 303538 479710
rect 305870 477053 305930 479710
rect 308446 477053 308506 479710
rect 305867 477052 305933 477053
rect 305867 476988 305868 477052
rect 305932 476988 305933 477052
rect 305867 476987 305933 476988
rect 308443 477052 308509 477053
rect 308443 476988 308444 477052
rect 308508 476988 308509 477052
rect 308443 476987 308509 476988
rect 311022 476917 311082 479710
rect 313414 479710 313500 479770
rect 315806 479710 315948 479770
rect 318382 479710 318532 479770
rect 320920 479770 320980 480080
rect 323368 479770 323428 480080
rect 325952 479770 326012 480080
rect 320920 479710 321018 479770
rect 311019 476916 311085 476917
rect 311019 476852 311020 476916
rect 311084 476852 311085 476916
rect 311019 476851 311085 476852
rect 303475 476780 303541 476781
rect 303475 476716 303476 476780
rect 303540 476716 303541 476780
rect 303475 476715 303541 476716
rect 313414 476509 313474 479710
rect 315806 476509 315866 479710
rect 313411 476508 313477 476509
rect 313411 476444 313412 476508
rect 313476 476444 313477 476508
rect 313411 476443 313477 476444
rect 315803 476508 315869 476509
rect 315803 476444 315804 476508
rect 315868 476444 315869 476508
rect 315803 476443 315869 476444
rect 318382 476373 318442 479710
rect 320958 476373 321018 479710
rect 323350 479710 323428 479770
rect 325926 479710 326012 479770
rect 323350 476781 323410 479710
rect 323347 476780 323413 476781
rect 323347 476716 323348 476780
rect 323412 476716 323413 476780
rect 323347 476715 323413 476716
rect 318379 476372 318445 476373
rect 318379 476308 318380 476372
rect 318444 476308 318445 476372
rect 318379 476307 318445 476308
rect 320955 476372 321021 476373
rect 320955 476308 320956 476372
rect 321020 476308 321021 476372
rect 320955 476307 321021 476308
rect 325926 476237 325986 479710
rect 235947 476236 236013 476237
rect 235947 476172 235948 476236
rect 236012 476172 236013 476236
rect 235947 476171 236013 476172
rect 237235 476236 237301 476237
rect 237235 476172 237236 476236
rect 237300 476172 237301 476236
rect 237235 476171 237301 476172
rect 239627 476236 239693 476237
rect 239627 476172 239628 476236
rect 239692 476172 239693 476236
rect 239627 476171 239693 476172
rect 240547 476236 240613 476237
rect 240547 476172 240548 476236
rect 240612 476172 240613 476236
rect 240547 476171 240613 476172
rect 241835 476236 241901 476237
rect 241835 476172 241836 476236
rect 241900 476172 241901 476236
rect 241835 476171 241901 476172
rect 246435 476236 246501 476237
rect 246435 476172 246436 476236
rect 246500 476172 246501 476236
rect 246435 476171 246501 476172
rect 247539 476236 247605 476237
rect 247539 476172 247540 476236
rect 247604 476172 247605 476236
rect 247539 476171 247605 476172
rect 248643 476236 248709 476237
rect 248643 476172 248644 476236
rect 248708 476172 248709 476236
rect 248643 476171 248709 476172
rect 250115 476236 250181 476237
rect 250115 476172 250116 476236
rect 250180 476172 250181 476236
rect 250115 476171 250181 476172
rect 251403 476236 251469 476237
rect 251403 476172 251404 476236
rect 251468 476172 251469 476236
rect 251403 476171 251469 476172
rect 253427 476236 253493 476237
rect 253427 476172 253428 476236
rect 253492 476172 253493 476236
rect 253427 476171 253493 476172
rect 254531 476236 254597 476237
rect 254531 476172 254532 476236
rect 254596 476172 254597 476236
rect 254531 476171 254597 476172
rect 255819 476236 255885 476237
rect 255819 476172 255820 476236
rect 255884 476172 255885 476236
rect 255819 476171 255885 476172
rect 257107 476236 257173 476237
rect 257107 476172 257108 476236
rect 257172 476172 257173 476236
rect 257107 476171 257173 476172
rect 259499 476236 259565 476237
rect 259499 476172 259500 476236
rect 259564 476172 259565 476236
rect 259499 476171 259565 476172
rect 261707 476236 261773 476237
rect 261707 476172 261708 476236
rect 261772 476172 261773 476236
rect 261707 476171 261773 476172
rect 263915 476236 263981 476237
rect 263915 476172 263916 476236
rect 263980 476172 263981 476236
rect 263915 476171 263981 476172
rect 265387 476236 265453 476237
rect 265387 476172 265388 476236
rect 265452 476172 265453 476236
rect 265387 476171 265453 476172
rect 267595 476236 267661 476237
rect 267595 476172 267596 476236
rect 267660 476172 267661 476236
rect 267595 476171 267661 476172
rect 268699 476236 268765 476237
rect 268699 476172 268700 476236
rect 268764 476172 268765 476236
rect 268699 476171 268765 476172
rect 269803 476236 269869 476237
rect 269803 476172 269804 476236
rect 269868 476172 269869 476236
rect 269803 476171 269869 476172
rect 271275 476236 271341 476237
rect 271275 476172 271276 476236
rect 271340 476172 271341 476236
rect 271275 476171 271341 476172
rect 272195 476236 272261 476237
rect 272195 476172 272196 476236
rect 272260 476172 272261 476236
rect 272195 476171 272261 476172
rect 274403 476236 274469 476237
rect 274403 476172 274404 476236
rect 274468 476172 274469 476236
rect 274403 476171 274469 476172
rect 275875 476236 275941 476237
rect 275875 476172 275876 476236
rect 275940 476172 275941 476236
rect 275875 476171 275941 476172
rect 278083 476236 278149 476237
rect 278083 476172 278084 476236
rect 278148 476172 278149 476236
rect 278083 476171 278149 476172
rect 279187 476236 279253 476237
rect 279187 476172 279188 476236
rect 279252 476172 279253 476236
rect 279187 476171 279253 476172
rect 283419 476236 283485 476237
rect 283419 476172 283420 476236
rect 283484 476172 283485 476236
rect 283419 476171 283485 476172
rect 285995 476236 286061 476237
rect 285995 476172 285996 476236
rect 286060 476172 286061 476236
rect 285995 476171 286061 476172
rect 288203 476236 288269 476237
rect 288203 476172 288204 476236
rect 288268 476172 288269 476236
rect 288203 476171 288269 476172
rect 290963 476236 291029 476237
rect 290963 476172 290964 476236
rect 291028 476172 291029 476236
rect 290963 476171 291029 476172
rect 293355 476236 293421 476237
rect 293355 476172 293356 476236
rect 293420 476172 293421 476236
rect 293355 476171 293421 476172
rect 295931 476236 295997 476237
rect 295931 476172 295932 476236
rect 295996 476172 295997 476236
rect 295931 476171 295997 476172
rect 298507 476236 298573 476237
rect 298507 476172 298508 476236
rect 298572 476172 298573 476236
rect 298507 476171 298573 476172
rect 300899 476236 300965 476237
rect 300899 476172 300900 476236
rect 300964 476172 300965 476236
rect 300899 476171 300965 476172
rect 325923 476236 325989 476237
rect 325923 476172 325924 476236
rect 325988 476172 325989 476236
rect 325923 476171 325989 476172
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 446026 362414 470898
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 364931 444684 364997 444685
rect 364931 444620 364932 444684
rect 364996 444620 364997 444684
rect 364931 444619 364997 444620
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 362539 443460 362605 443461
rect 362539 443396 362540 443460
rect 362604 443396 362605 443460
rect 362539 443395 362605 443396
rect 362723 443460 362789 443461
rect 362723 443396 362724 443460
rect 362788 443396 362789 443460
rect 362723 443395 362789 443396
rect 362907 443460 362973 443461
rect 362907 443396 362908 443460
rect 362972 443396 362973 443460
rect 362907 443395 362973 443396
rect 251968 439954 252288 439986
rect 251968 439718 252010 439954
rect 252246 439718 252288 439954
rect 251968 439634 252288 439718
rect 251968 439398 252010 439634
rect 252246 439398 252288 439634
rect 251968 439366 252288 439398
rect 282688 439954 283008 439986
rect 282688 439718 282730 439954
rect 282966 439718 283008 439954
rect 282688 439634 283008 439718
rect 282688 439398 282730 439634
rect 282966 439398 283008 439634
rect 282688 439366 283008 439398
rect 313408 439954 313728 439986
rect 313408 439718 313450 439954
rect 313686 439718 313728 439954
rect 313408 439634 313728 439718
rect 313408 439398 313450 439634
rect 313686 439398 313728 439634
rect 313408 439366 313728 439398
rect 344128 439954 344448 439986
rect 344128 439718 344170 439954
rect 344406 439718 344448 439954
rect 344128 439634 344448 439718
rect 344128 439398 344170 439634
rect 344406 439398 344448 439634
rect 344128 439366 344448 439398
rect 236608 435454 236928 435486
rect 236608 435218 236650 435454
rect 236886 435218 236928 435454
rect 236608 435134 236928 435218
rect 236608 434898 236650 435134
rect 236886 434898 236928 435134
rect 236608 434866 236928 434898
rect 267328 435454 267648 435486
rect 267328 435218 267370 435454
rect 267606 435218 267648 435454
rect 267328 435134 267648 435218
rect 267328 434898 267370 435134
rect 267606 434898 267648 435134
rect 267328 434866 267648 434898
rect 298048 435454 298368 435486
rect 298048 435218 298090 435454
rect 298326 435218 298368 435454
rect 298048 435134 298368 435218
rect 298048 434898 298090 435134
rect 298326 434898 298368 435134
rect 298048 434866 298368 434898
rect 328768 435454 329088 435486
rect 328768 435218 328810 435454
rect 329046 435218 329088 435454
rect 328768 435134 329088 435218
rect 328768 434898 328810 435134
rect 329046 434898 329088 435134
rect 328768 434866 329088 434898
rect 359488 435454 359808 435486
rect 359488 435218 359530 435454
rect 359766 435218 359808 435454
rect 359488 435134 359808 435218
rect 359488 434898 359530 435134
rect 359766 434898 359808 435134
rect 359488 434866 359808 434898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 251968 403954 252288 403986
rect 251968 403718 252010 403954
rect 252246 403718 252288 403954
rect 251968 403634 252288 403718
rect 251968 403398 252010 403634
rect 252246 403398 252288 403634
rect 251968 403366 252288 403398
rect 282688 403954 283008 403986
rect 282688 403718 282730 403954
rect 282966 403718 283008 403954
rect 282688 403634 283008 403718
rect 282688 403398 282730 403634
rect 282966 403398 283008 403634
rect 282688 403366 283008 403398
rect 313408 403954 313728 403986
rect 313408 403718 313450 403954
rect 313686 403718 313728 403954
rect 313408 403634 313728 403718
rect 313408 403398 313450 403634
rect 313686 403398 313728 403634
rect 313408 403366 313728 403398
rect 344128 403954 344448 403986
rect 344128 403718 344170 403954
rect 344406 403718 344448 403954
rect 344128 403634 344448 403718
rect 344128 403398 344170 403634
rect 344406 403398 344448 403634
rect 344128 403366 344448 403398
rect 236608 399454 236928 399486
rect 236608 399218 236650 399454
rect 236886 399218 236928 399454
rect 236608 399134 236928 399218
rect 236608 398898 236650 399134
rect 236886 398898 236928 399134
rect 236608 398866 236928 398898
rect 267328 399454 267648 399486
rect 267328 399218 267370 399454
rect 267606 399218 267648 399454
rect 267328 399134 267648 399218
rect 267328 398898 267370 399134
rect 267606 398898 267648 399134
rect 267328 398866 267648 398898
rect 298048 399454 298368 399486
rect 298048 399218 298090 399454
rect 298326 399218 298368 399454
rect 298048 399134 298368 399218
rect 298048 398898 298090 399134
rect 298326 398898 298368 399134
rect 298048 398866 298368 398898
rect 328768 399454 329088 399486
rect 328768 399218 328810 399454
rect 329046 399218 329088 399454
rect 328768 399134 329088 399218
rect 328768 398898 328810 399134
rect 329046 398898 329088 399134
rect 328768 398866 329088 398898
rect 359488 399454 359808 399486
rect 359488 399218 359530 399454
rect 359766 399218 359808 399454
rect 359488 399134 359808 399218
rect 359488 398898 359530 399134
rect 359766 398898 359808 399134
rect 359488 398866 359808 398898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 251968 367954 252288 367986
rect 251968 367718 252010 367954
rect 252246 367718 252288 367954
rect 251968 367634 252288 367718
rect 251968 367398 252010 367634
rect 252246 367398 252288 367634
rect 251968 367366 252288 367398
rect 282688 367954 283008 367986
rect 282688 367718 282730 367954
rect 282966 367718 283008 367954
rect 282688 367634 283008 367718
rect 282688 367398 282730 367634
rect 282966 367398 283008 367634
rect 282688 367366 283008 367398
rect 313408 367954 313728 367986
rect 313408 367718 313450 367954
rect 313686 367718 313728 367954
rect 313408 367634 313728 367718
rect 313408 367398 313450 367634
rect 313686 367398 313728 367634
rect 313408 367366 313728 367398
rect 344128 367954 344448 367986
rect 344128 367718 344170 367954
rect 344406 367718 344448 367954
rect 344128 367634 344448 367718
rect 344128 367398 344170 367634
rect 344406 367398 344448 367634
rect 344128 367366 344448 367398
rect 236608 363454 236928 363486
rect 236608 363218 236650 363454
rect 236886 363218 236928 363454
rect 236608 363134 236928 363218
rect 236608 362898 236650 363134
rect 236886 362898 236928 363134
rect 236608 362866 236928 362898
rect 267328 363454 267648 363486
rect 267328 363218 267370 363454
rect 267606 363218 267648 363454
rect 267328 363134 267648 363218
rect 267328 362898 267370 363134
rect 267606 362898 267648 363134
rect 267328 362866 267648 362898
rect 298048 363454 298368 363486
rect 298048 363218 298090 363454
rect 298326 363218 298368 363454
rect 298048 363134 298368 363218
rect 298048 362898 298090 363134
rect 298326 362898 298368 363134
rect 298048 362866 298368 362898
rect 328768 363454 329088 363486
rect 328768 363218 328810 363454
rect 329046 363218 329088 363454
rect 328768 363134 329088 363218
rect 328768 362898 328810 363134
rect 329046 362898 329088 363134
rect 328768 362866 329088 362898
rect 359488 363454 359808 363486
rect 359488 363218 359530 363454
rect 359766 363218 359808 363454
rect 359488 363134 359808 363218
rect 359488 362898 359530 363134
rect 359766 362898 359808 363134
rect 359488 362866 359808 362898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 251968 331954 252288 331986
rect 251968 331718 252010 331954
rect 252246 331718 252288 331954
rect 251968 331634 252288 331718
rect 251968 331398 252010 331634
rect 252246 331398 252288 331634
rect 251968 331366 252288 331398
rect 282688 331954 283008 331986
rect 282688 331718 282730 331954
rect 282966 331718 283008 331954
rect 282688 331634 283008 331718
rect 282688 331398 282730 331634
rect 282966 331398 283008 331634
rect 282688 331366 283008 331398
rect 313408 331954 313728 331986
rect 313408 331718 313450 331954
rect 313686 331718 313728 331954
rect 313408 331634 313728 331718
rect 313408 331398 313450 331634
rect 313686 331398 313728 331634
rect 313408 331366 313728 331398
rect 344128 331954 344448 331986
rect 344128 331718 344170 331954
rect 344406 331718 344448 331954
rect 344128 331634 344448 331718
rect 344128 331398 344170 331634
rect 344406 331398 344448 331634
rect 344128 331366 344448 331398
rect 236608 327454 236928 327486
rect 236608 327218 236650 327454
rect 236886 327218 236928 327454
rect 236608 327134 236928 327218
rect 236608 326898 236650 327134
rect 236886 326898 236928 327134
rect 236608 326866 236928 326898
rect 267328 327454 267648 327486
rect 267328 327218 267370 327454
rect 267606 327218 267648 327454
rect 267328 327134 267648 327218
rect 267328 326898 267370 327134
rect 267606 326898 267648 327134
rect 267328 326866 267648 326898
rect 298048 327454 298368 327486
rect 298048 327218 298090 327454
rect 298326 327218 298368 327454
rect 298048 327134 298368 327218
rect 298048 326898 298090 327134
rect 298326 326898 298368 327134
rect 298048 326866 298368 326898
rect 328768 327454 329088 327486
rect 328768 327218 328810 327454
rect 329046 327218 329088 327454
rect 328768 327134 329088 327218
rect 328768 326898 328810 327134
rect 329046 326898 329088 327134
rect 328768 326866 329088 326898
rect 359488 327454 359808 327486
rect 359488 327218 359530 327454
rect 359766 327218 359808 327454
rect 359488 327134 359808 327218
rect 359488 326898 359530 327134
rect 359766 326898 359808 327134
rect 359488 326866 359808 326898
rect 358859 308548 358925 308549
rect 358859 308484 358860 308548
rect 358924 308484 358925 308548
rect 358859 308483 358925 308484
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 245308 227414 263898
rect 231294 304954 231914 308400
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 245308 231914 268398
rect 244794 282454 245414 308400
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 246454 245414 281898
rect 244794 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 245414 246454
rect 244794 246134 245414 246218
rect 244794 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 245414 246134
rect 244794 245308 245414 245898
rect 249294 286954 249914 308400
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 245308 249914 250398
rect 253794 291454 254414 308400
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 245308 254414 254898
rect 258294 295954 258914 308400
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 245308 258914 259398
rect 262794 300454 263414 308400
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 245308 263414 263898
rect 267294 304954 267914 308400
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 245308 267914 268398
rect 280794 282454 281414 308400
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 246454 281414 281898
rect 280794 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 281414 246454
rect 280794 246134 281414 246218
rect 280794 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 281414 246134
rect 280794 245308 281414 245898
rect 285294 286954 285914 308400
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 245308 285914 250398
rect 289794 291454 290414 308400
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 245308 290414 254898
rect 294294 295954 294914 308400
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 245308 294914 259398
rect 298794 300454 299414 308400
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 245308 299414 263898
rect 303294 304954 303914 308400
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 245308 303914 268398
rect 316794 282454 317414 308400
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 246454 317414 281898
rect 316794 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 317414 246454
rect 316794 246134 317414 246218
rect 316794 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 317414 246134
rect 316794 245308 317414 245898
rect 321294 286954 321914 308400
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 245308 321914 250398
rect 325794 291454 326414 308400
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 245308 326414 254898
rect 330294 295954 330914 308400
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 245308 330914 259398
rect 334794 300454 335414 308400
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 245308 335414 263898
rect 339294 304954 339914 308400
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 245308 339914 268398
rect 352794 282454 353414 308400
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 245308 353414 245898
rect 357294 286954 357914 308400
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 245308 357914 250398
rect 358123 248164 358189 248165
rect 358123 248100 358124 248164
rect 358188 248100 358189 248164
rect 358123 248099 358189 248100
rect 357939 245172 358005 245173
rect 357939 245108 357940 245172
rect 358004 245108 358005 245172
rect 357939 245107 358005 245108
rect 220272 223954 220620 223986
rect 220272 223718 220328 223954
rect 220564 223718 220620 223954
rect 220272 223634 220620 223718
rect 220272 223398 220328 223634
rect 220564 223398 220620 223634
rect 220272 223366 220620 223398
rect 356000 223954 356348 223986
rect 356000 223718 356056 223954
rect 356292 223718 356348 223954
rect 356000 223634 356348 223718
rect 356000 223398 356056 223634
rect 356292 223398 356348 223634
rect 356000 223366 356348 223398
rect 220952 219454 221300 219486
rect 220952 219218 221008 219454
rect 221244 219218 221300 219454
rect 220952 219134 221300 219218
rect 220952 218898 221008 219134
rect 221244 218898 221300 219134
rect 220952 218866 221300 218898
rect 355320 219454 355668 219486
rect 355320 219218 355376 219454
rect 355612 219218 355668 219454
rect 355320 219134 355668 219218
rect 355320 218898 355376 219134
rect 355612 218898 355668 219134
rect 355320 218866 355668 218898
rect 220272 187954 220620 187986
rect 220272 187718 220328 187954
rect 220564 187718 220620 187954
rect 220272 187634 220620 187718
rect 220272 187398 220328 187634
rect 220564 187398 220620 187634
rect 220272 187366 220620 187398
rect 356000 187954 356348 187986
rect 356000 187718 356056 187954
rect 356292 187718 356348 187954
rect 356000 187634 356348 187718
rect 356000 187398 356056 187634
rect 356292 187398 356348 187634
rect 356000 187366 356348 187398
rect 220952 183454 221300 183486
rect 220952 183218 221008 183454
rect 221244 183218 221300 183454
rect 220952 183134 221300 183218
rect 220952 182898 221008 183134
rect 221244 182898 221300 183134
rect 220952 182866 221300 182898
rect 355320 183454 355668 183486
rect 355320 183218 355376 183454
rect 355612 183218 355668 183454
rect 355320 183134 355668 183218
rect 355320 182898 355376 183134
rect 355612 182898 355668 183134
rect 355320 182866 355668 182898
rect 236056 159490 236116 160106
rect 237144 159490 237204 160106
rect 238232 159490 238292 160106
rect 236056 159430 236194 159490
rect 237144 159430 237298 159490
rect 236134 158541 236194 159430
rect 236131 158540 236197 158541
rect 236131 158476 236132 158540
rect 236196 158476 236197 158540
rect 236131 158475 236197 158476
rect 222294 151954 222914 158000
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 219203 3636 219269 3637
rect 219203 3572 219204 3636
rect 219268 3572 219269 3636
rect 219203 3571 219269 3572
rect 215891 3364 215957 3365
rect 215891 3300 215892 3364
rect 215956 3300 215957 3364
rect 215891 3299 215957 3300
rect 217547 3364 217613 3365
rect 217547 3300 217548 3364
rect 217612 3300 217613 3364
rect 217547 3299 217613 3300
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 218651 3500 218717 3501
rect 218651 3436 218652 3500
rect 218716 3436 218717 3500
rect 218651 3435 218717 3436
rect 219019 3500 219085 3501
rect 219019 3436 219020 3500
rect 219084 3436 219085 3500
rect 219019 3435 219085 3436
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 156454 227414 158000
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 124954 231914 158000
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 129454 236414 158000
rect 237238 157453 237298 159430
rect 238158 159430 238292 159490
rect 239592 159490 239652 160106
rect 240544 159490 240604 160106
rect 241768 159490 241828 160106
rect 243128 159490 243188 160106
rect 239592 159430 239690 159490
rect 240544 159430 240610 159490
rect 241768 159430 241898 159490
rect 238158 158677 238218 159430
rect 239630 158677 239690 159430
rect 238155 158676 238221 158677
rect 238155 158612 238156 158676
rect 238220 158612 238221 158676
rect 238155 158611 238221 158612
rect 239627 158676 239693 158677
rect 239627 158612 239628 158676
rect 239692 158612 239693 158676
rect 239627 158611 239693 158612
rect 240550 158269 240610 159430
rect 241838 158677 241898 159430
rect 243126 159430 243188 159490
rect 244216 159490 244276 160106
rect 245440 159490 245500 160106
rect 246528 159490 246588 160106
rect 247616 159490 247676 160106
rect 248296 159490 248356 160106
rect 248704 159490 248764 160106
rect 244216 159430 244290 159490
rect 245440 159430 245578 159490
rect 246528 159430 246682 159490
rect 247616 159430 247786 159490
rect 243126 158813 243186 159430
rect 243123 158812 243189 158813
rect 243123 158748 243124 158812
rect 243188 158748 243189 158812
rect 243123 158747 243189 158748
rect 244230 158677 244290 159430
rect 245518 158677 245578 159430
rect 241835 158676 241901 158677
rect 241835 158612 241836 158676
rect 241900 158612 241901 158676
rect 241835 158611 241901 158612
rect 244227 158676 244293 158677
rect 244227 158612 244228 158676
rect 244292 158612 244293 158676
rect 244227 158611 244293 158612
rect 245515 158676 245581 158677
rect 245515 158612 245516 158676
rect 245580 158612 245581 158676
rect 245515 158611 245581 158612
rect 240547 158268 240613 158269
rect 240547 158204 240548 158268
rect 240612 158204 240613 158268
rect 240547 158203 240613 158204
rect 237235 157452 237301 157453
rect 237235 157388 237236 157452
rect 237300 157388 237301 157452
rect 237235 157387 237301 157388
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 133954 240914 158000
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 138454 245414 158000
rect 246622 157997 246682 159430
rect 247726 157997 247786 159430
rect 248278 159430 248356 159490
rect 248646 159430 248764 159490
rect 250064 159490 250124 160106
rect 250744 159490 250804 160106
rect 251288 159490 251348 160106
rect 252376 159490 252436 160106
rect 253464 159490 253524 160106
rect 250064 159430 250178 159490
rect 250744 159430 250914 159490
rect 251288 159430 251466 159490
rect 248278 158677 248338 159430
rect 248275 158676 248341 158677
rect 248275 158612 248276 158676
rect 248340 158612 248341 158676
rect 248275 158611 248341 158612
rect 246619 157996 246685 157997
rect 246619 157932 246620 157996
rect 246684 157932 246685 157996
rect 246619 157931 246685 157932
rect 247723 157996 247789 157997
rect 247723 157932 247724 157996
rect 247788 157932 247789 157996
rect 247723 157931 247789 157932
rect 248646 157861 248706 159430
rect 248643 157860 248709 157861
rect 248643 157796 248644 157860
rect 248708 157796 248709 157860
rect 248643 157795 248709 157796
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 142954 249914 158000
rect 250118 157861 250178 159430
rect 250854 157997 250914 159430
rect 250851 157996 250917 157997
rect 250851 157932 250852 157996
rect 250916 157932 250917 157996
rect 250851 157931 250917 157932
rect 251406 157861 251466 159430
rect 252326 159430 252436 159490
rect 253430 159430 253524 159490
rect 253600 159490 253660 160106
rect 254552 159490 254612 160106
rect 255912 159490 255972 160106
rect 253600 159430 253674 159490
rect 252326 158677 252386 159430
rect 252323 158676 252389 158677
rect 252323 158612 252324 158676
rect 252388 158612 252389 158676
rect 252323 158611 252389 158612
rect 253430 157861 253490 159430
rect 253614 158949 253674 159430
rect 254534 159430 254612 159490
rect 255822 159430 255972 159490
rect 256048 159490 256108 160106
rect 257000 159490 257060 160106
rect 258088 159490 258148 160106
rect 258496 159490 258556 160106
rect 259448 159490 259508 160106
rect 260672 159629 260732 160106
rect 261080 159765 261140 160106
rect 261077 159764 261143 159765
rect 261077 159700 261078 159764
rect 261142 159700 261143 159764
rect 261077 159699 261143 159700
rect 260669 159628 260735 159629
rect 260669 159564 260670 159628
rect 260734 159564 260735 159628
rect 260669 159563 260735 159564
rect 261760 159490 261820 160106
rect 262848 159490 262908 160106
rect 256048 159430 256250 159490
rect 257000 159430 257170 159490
rect 258088 159430 258274 159490
rect 258496 159430 258642 159490
rect 259448 159430 259562 159490
rect 254534 159085 254594 159430
rect 254531 159084 254597 159085
rect 254531 159020 254532 159084
rect 254596 159020 254597 159084
rect 254531 159019 254597 159020
rect 253611 158948 253677 158949
rect 253611 158884 253612 158948
rect 253676 158884 253677 158948
rect 253611 158883 253677 158884
rect 255822 158677 255882 159430
rect 255819 158676 255885 158677
rect 255819 158612 255820 158676
rect 255884 158612 255885 158676
rect 255819 158611 255885 158612
rect 250115 157860 250181 157861
rect 250115 157796 250116 157860
rect 250180 157796 250181 157860
rect 250115 157795 250181 157796
rect 251403 157860 251469 157861
rect 251403 157796 251404 157860
rect 251468 157796 251469 157860
rect 251403 157795 251469 157796
rect 253427 157860 253493 157861
rect 253427 157796 253428 157860
rect 253492 157796 253493 157860
rect 253427 157795 253493 157796
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 147454 254414 158000
rect 256190 157589 256250 159430
rect 257110 158677 257170 159430
rect 257107 158676 257173 158677
rect 257107 158612 257108 158676
rect 257172 158612 257173 158676
rect 257107 158611 257173 158612
rect 258214 158405 258274 159430
rect 258211 158404 258277 158405
rect 258211 158340 258212 158404
rect 258276 158340 258277 158404
rect 258211 158339 258277 158340
rect 258582 158269 258642 159430
rect 259502 159221 259562 159430
rect 261710 159430 261820 159490
rect 262630 159430 262908 159490
rect 263528 159490 263588 160106
rect 263936 159490 263996 160106
rect 263528 159430 263610 159490
rect 259499 159220 259565 159221
rect 259499 159156 259500 159220
rect 259564 159156 259565 159220
rect 259499 159155 259565 159156
rect 261710 158677 261770 159430
rect 261707 158676 261773 158677
rect 261707 158612 261708 158676
rect 261772 158612 261773 158676
rect 261707 158611 261773 158612
rect 258579 158268 258645 158269
rect 258579 158204 258580 158268
rect 258644 158204 258645 158268
rect 258579 158203 258645 158204
rect 262630 158133 262690 159430
rect 262627 158132 262693 158133
rect 262627 158068 262628 158132
rect 262692 158068 262693 158132
rect 262627 158067 262693 158068
rect 256187 157588 256253 157589
rect 256187 157524 256188 157588
rect 256252 157524 256253 157588
rect 256187 157523 256253 157524
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 151954 258914 158000
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 156454 263414 158000
rect 263550 157589 263610 159430
rect 263918 159430 263996 159490
rect 265296 159490 265356 160106
rect 265976 159490 266036 160106
rect 265296 159430 265450 159490
rect 263918 157861 263978 159430
rect 265390 158677 265450 159430
rect 265942 159430 266036 159490
rect 266384 159490 266444 160106
rect 267608 159490 267668 160106
rect 266384 159430 266554 159490
rect 265942 158677 266002 159430
rect 266494 158677 266554 159430
rect 267046 159430 267668 159490
rect 268288 159490 268348 160106
rect 268696 159490 268756 160106
rect 269784 159490 269844 160106
rect 271008 159490 271068 160106
rect 268288 159430 268394 159490
rect 268696 159430 268762 159490
rect 269784 159430 269866 159490
rect 265387 158676 265453 158677
rect 265387 158612 265388 158676
rect 265452 158612 265453 158676
rect 265387 158611 265453 158612
rect 265939 158676 266005 158677
rect 265939 158612 265940 158676
rect 266004 158612 266005 158676
rect 265939 158611 266005 158612
rect 266491 158676 266557 158677
rect 266491 158612 266492 158676
rect 266556 158612 266557 158676
rect 266491 158611 266557 158612
rect 267046 157997 267106 159430
rect 267043 157996 267109 157997
rect 267043 157932 267044 157996
rect 267108 157932 267109 157996
rect 267043 157931 267109 157932
rect 263915 157860 263981 157861
rect 263915 157796 263916 157860
rect 263980 157796 263981 157860
rect 263915 157795 263981 157796
rect 263547 157588 263613 157589
rect 263547 157524 263548 157588
rect 263612 157524 263613 157588
rect 263547 157523 263613 157524
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 124954 267914 158000
rect 268334 157725 268394 159430
rect 268702 158677 268762 159430
rect 269806 158677 269866 159430
rect 270910 159430 271068 159490
rect 271144 159490 271204 160106
rect 272232 159490 272292 160106
rect 273320 159901 273380 160106
rect 273317 159900 273383 159901
rect 273317 159836 273318 159900
rect 273382 159836 273383 159900
rect 273317 159835 273383 159836
rect 271144 159430 271338 159490
rect 270910 158677 270970 159430
rect 268699 158676 268765 158677
rect 268699 158612 268700 158676
rect 268764 158612 268765 158676
rect 268699 158611 268765 158612
rect 269803 158676 269869 158677
rect 269803 158612 269804 158676
rect 269868 158612 269869 158676
rect 269803 158611 269869 158612
rect 270907 158676 270973 158677
rect 270907 158612 270908 158676
rect 270972 158612 270973 158676
rect 270907 158611 270973 158612
rect 271278 157725 271338 159430
rect 272198 159430 272292 159490
rect 273592 159490 273652 160106
rect 274408 159490 274468 160106
rect 275768 159629 275828 160106
rect 275765 159628 275831 159629
rect 275765 159564 275766 159628
rect 275830 159564 275831 159628
rect 275765 159563 275831 159564
rect 273592 159430 273730 159490
rect 272198 158677 272258 159430
rect 272195 158676 272261 158677
rect 272195 158612 272196 158676
rect 272260 158612 272261 158676
rect 272195 158611 272261 158612
rect 268331 157724 268397 157725
rect 268331 157660 268332 157724
rect 268396 157660 268397 157724
rect 268331 157659 268397 157660
rect 271275 157724 271341 157725
rect 271275 157660 271276 157724
rect 271340 157660 271341 157724
rect 271275 157659 271341 157660
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 129454 272414 158000
rect 273670 157725 273730 159430
rect 274406 159430 274468 159490
rect 276040 159490 276100 160106
rect 276992 159629 277052 160106
rect 278080 159901 278140 160106
rect 278077 159900 278143 159901
rect 278077 159836 278078 159900
rect 278142 159836 278143 159900
rect 278077 159835 278143 159836
rect 276989 159628 277055 159629
rect 276989 159564 276990 159628
rect 277054 159564 277055 159628
rect 276989 159563 277055 159564
rect 278488 159490 278548 160106
rect 279168 159629 279228 160106
rect 279165 159628 279231 159629
rect 279165 159564 279166 159628
rect 279230 159564 279231 159628
rect 280936 159626 280996 160106
rect 283520 159626 283580 160106
rect 280936 159566 281090 159626
rect 283520 159566 283666 159626
rect 279165 159563 279231 159564
rect 276040 159430 276122 159490
rect 274406 158677 274466 159430
rect 276062 158677 276122 159430
rect 278454 159430 278548 159490
rect 274403 158676 274469 158677
rect 274403 158612 274404 158676
rect 274468 158612 274469 158676
rect 274403 158611 274469 158612
rect 276059 158676 276125 158677
rect 276059 158612 276060 158676
rect 276124 158612 276125 158676
rect 276059 158611 276125 158612
rect 273667 157724 273733 157725
rect 273667 157660 273668 157724
rect 273732 157660 273733 157724
rect 273667 157659 273733 157660
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 133954 276914 158000
rect 278454 157725 278514 159430
rect 281030 158677 281090 159566
rect 281027 158676 281093 158677
rect 281027 158612 281028 158676
rect 281092 158612 281093 158676
rect 281027 158611 281093 158612
rect 278451 157724 278517 157725
rect 278451 157660 278452 157724
rect 278516 157660 278517 157724
rect 278451 157659 278517 157660
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 138454 281414 158000
rect 283606 157589 283666 159566
rect 285968 159490 286028 160106
rect 288280 159490 288340 160106
rect 291000 159490 291060 160106
rect 285968 159430 286058 159490
rect 283603 157588 283669 157589
rect 283603 157524 283604 157588
rect 283668 157524 283669 157588
rect 283603 157523 283669 157524
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 142954 285914 158000
rect 285998 157589 286058 159430
rect 288206 159430 288340 159490
rect 290966 159430 291060 159490
rect 293448 159490 293508 160106
rect 295896 159490 295956 160106
rect 298480 159490 298540 160106
rect 300928 159490 300988 160106
rect 303512 159490 303572 160106
rect 293448 159430 293602 159490
rect 295896 159430 295994 159490
rect 298480 159430 298570 159490
rect 288206 158677 288266 159430
rect 290966 158677 291026 159430
rect 293542 158677 293602 159430
rect 295934 158677 295994 159430
rect 298510 158677 298570 159430
rect 300902 159430 300988 159490
rect 303478 159430 303572 159490
rect 305960 159490 306020 160106
rect 308544 159490 308604 160106
rect 310992 159490 311052 160106
rect 313440 159490 313500 160106
rect 315888 159490 315948 160106
rect 305960 159430 306114 159490
rect 308544 159430 308690 159490
rect 310992 159430 311082 159490
rect 300902 158677 300962 159430
rect 303478 158677 303538 159430
rect 306054 158677 306114 159430
rect 308630 158677 308690 159430
rect 311022 158677 311082 159430
rect 313414 159430 313500 159490
rect 315806 159430 315948 159490
rect 318472 159490 318532 160106
rect 320920 159490 320980 160106
rect 323368 159490 323428 160106
rect 325952 159490 326012 160106
rect 318472 159430 318626 159490
rect 320920 159430 321018 159490
rect 313414 158677 313474 159430
rect 315806 158677 315866 159430
rect 318566 158677 318626 159430
rect 320958 158677 321018 159430
rect 323350 159430 323428 159490
rect 325926 159430 326012 159490
rect 323350 158677 323410 159430
rect 325926 158677 325986 159430
rect 357942 159357 358002 245107
rect 357939 159356 358005 159357
rect 357939 159292 357940 159356
rect 358004 159292 358005 159356
rect 357939 159291 358005 159292
rect 288203 158676 288269 158677
rect 288203 158612 288204 158676
rect 288268 158612 288269 158676
rect 288203 158611 288269 158612
rect 290963 158676 291029 158677
rect 290963 158612 290964 158676
rect 291028 158612 291029 158676
rect 290963 158611 291029 158612
rect 293539 158676 293605 158677
rect 293539 158612 293540 158676
rect 293604 158612 293605 158676
rect 293539 158611 293605 158612
rect 295931 158676 295997 158677
rect 295931 158612 295932 158676
rect 295996 158612 295997 158676
rect 295931 158611 295997 158612
rect 298507 158676 298573 158677
rect 298507 158612 298508 158676
rect 298572 158612 298573 158676
rect 298507 158611 298573 158612
rect 300899 158676 300965 158677
rect 300899 158612 300900 158676
rect 300964 158612 300965 158676
rect 300899 158611 300965 158612
rect 303475 158676 303541 158677
rect 303475 158612 303476 158676
rect 303540 158612 303541 158676
rect 303475 158611 303541 158612
rect 306051 158676 306117 158677
rect 306051 158612 306052 158676
rect 306116 158612 306117 158676
rect 306051 158611 306117 158612
rect 308627 158676 308693 158677
rect 308627 158612 308628 158676
rect 308692 158612 308693 158676
rect 308627 158611 308693 158612
rect 311019 158676 311085 158677
rect 311019 158612 311020 158676
rect 311084 158612 311085 158676
rect 311019 158611 311085 158612
rect 313411 158676 313477 158677
rect 313411 158612 313412 158676
rect 313476 158612 313477 158676
rect 313411 158611 313477 158612
rect 315803 158676 315869 158677
rect 315803 158612 315804 158676
rect 315868 158612 315869 158676
rect 315803 158611 315869 158612
rect 318563 158676 318629 158677
rect 318563 158612 318564 158676
rect 318628 158612 318629 158676
rect 318563 158611 318629 158612
rect 320955 158676 321021 158677
rect 320955 158612 320956 158676
rect 321020 158612 321021 158676
rect 320955 158611 321021 158612
rect 323347 158676 323413 158677
rect 323347 158612 323348 158676
rect 323412 158612 323413 158676
rect 323347 158611 323413 158612
rect 325923 158676 325989 158677
rect 325923 158612 325924 158676
rect 325988 158612 325989 158676
rect 325923 158611 325989 158612
rect 285995 157588 286061 157589
rect 285995 157524 285996 157588
rect 286060 157524 286061 157588
rect 285995 157523 286061 157524
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 147454 290414 158000
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 151954 294914 158000
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 156454 299414 158000
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 124954 303914 158000
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 129454 308414 158000
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 133954 312914 158000
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 138454 317414 158000
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 142954 321914 158000
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 147454 326414 158000
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 151954 330914 158000
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 156454 335414 158000
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 124954 339914 158000
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 129454 344414 158000
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 133954 348914 158000
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 138454 353414 158000
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 142954 357914 158000
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 358126 3501 358186 248099
rect 358307 245580 358373 245581
rect 358307 245516 358308 245580
rect 358372 245516 358373 245580
rect 358307 245515 358373 245516
rect 358310 3501 358370 245515
rect 358491 245036 358557 245037
rect 358491 244972 358492 245036
rect 358556 244972 358557 245036
rect 358491 244971 358557 244972
rect 358123 3500 358189 3501
rect 358123 3436 358124 3500
rect 358188 3436 358189 3500
rect 358123 3435 358189 3436
rect 358307 3500 358373 3501
rect 358307 3436 358308 3500
rect 358372 3436 358373 3500
rect 358307 3435 358373 3436
rect 358494 3365 358554 244971
rect 358862 3909 358922 308483
rect 360331 308412 360397 308413
rect 360331 308348 360332 308412
rect 360396 308348 360397 308412
rect 360331 308347 360397 308348
rect 360334 302250 360394 308347
rect 360150 302190 360394 302250
rect 359043 260132 359109 260133
rect 359043 260068 359044 260132
rect 359108 260068 359109 260132
rect 359043 260067 359109 260068
rect 358859 3908 358925 3909
rect 358859 3844 358860 3908
rect 358924 3844 358925 3908
rect 358859 3843 358925 3844
rect 359046 3501 359106 260067
rect 359227 245444 359293 245445
rect 359227 245380 359228 245444
rect 359292 245380 359293 245444
rect 359227 245379 359293 245380
rect 359043 3500 359109 3501
rect 359043 3436 359044 3500
rect 359108 3436 359109 3500
rect 359043 3435 359109 3436
rect 358491 3364 358557 3365
rect 358491 3300 358492 3364
rect 358556 3300 358557 3364
rect 358491 3299 358557 3300
rect 359230 3229 359290 245379
rect 359411 245308 359477 245309
rect 359411 245244 359412 245308
rect 359476 245244 359477 245308
rect 359411 245243 359477 245244
rect 359414 3637 359474 245243
rect 360150 4045 360210 302190
rect 361794 291454 362414 308400
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 360331 284884 360397 284885
rect 360331 284820 360332 284884
rect 360396 284820 360397 284884
rect 360331 284819 360397 284820
rect 360147 4044 360213 4045
rect 360147 3980 360148 4044
rect 360212 3980 360213 4044
rect 360147 3979 360213 3980
rect 359411 3636 359477 3637
rect 359411 3572 359412 3636
rect 359476 3572 359477 3636
rect 359411 3571 359477 3572
rect 360334 3501 360394 284819
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 360699 250748 360765 250749
rect 360699 250684 360700 250748
rect 360764 250684 360765 250748
rect 360699 250683 360765 250684
rect 360515 244900 360581 244901
rect 360515 244836 360516 244900
rect 360580 244836 360581 244900
rect 360515 244835 360581 244836
rect 360518 3773 360578 244835
rect 360702 159357 360762 250683
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 360699 159356 360765 159357
rect 360699 159292 360700 159356
rect 360764 159292 360765 159356
rect 360699 159291 360765 159292
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 362542 84285 362602 443395
rect 362539 84284 362605 84285
rect 362539 84220 362540 84284
rect 362604 84220 362605 84284
rect 362539 84219 362605 84220
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 362726 44301 362786 443395
rect 362723 44300 362789 44301
rect 362723 44236 362724 44300
rect 362788 44236 362789 44300
rect 362723 44235 362789 44236
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 360515 3772 360581 3773
rect 360515 3708 360516 3772
rect 360580 3708 360581 3772
rect 360515 3707 360581 3708
rect 360331 3500 360397 3501
rect 360331 3436 360332 3500
rect 360396 3436 360397 3500
rect 360331 3435 360397 3436
rect 361794 3454 362414 38898
rect 362910 5677 362970 443395
rect 363091 267068 363157 267069
rect 363091 267004 363092 267068
rect 363156 267004 363157 267068
rect 363091 267003 363157 267004
rect 362907 5676 362973 5677
rect 362907 5612 362908 5676
rect 362972 5612 362973 5676
rect 362907 5611 362973 5612
rect 363094 3501 363154 267003
rect 363459 262852 363525 262853
rect 363459 262788 363460 262852
rect 363524 262788 363525 262852
rect 363459 262787 363525 262788
rect 363275 244628 363341 244629
rect 363275 244564 363276 244628
rect 363340 244564 363341 244628
rect 363275 244563 363341 244564
rect 363278 159357 363338 244563
rect 363275 159356 363341 159357
rect 363275 159292 363276 159356
rect 363340 159292 363341 159356
rect 363275 159291 363341 159292
rect 359227 3228 359293 3229
rect 359227 3164 359228 3228
rect 359292 3164 359293 3228
rect 359227 3163 359293 3164
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 363091 3500 363157 3501
rect 363091 3436 363092 3500
rect 363156 3436 363157 3500
rect 363091 3435 363157 3436
rect 363462 3365 363522 262787
rect 364379 249116 364445 249117
rect 364379 249052 364380 249116
rect 364444 249052 364445 249116
rect 364379 249051 364445 249052
rect 364382 3501 364442 249051
rect 364934 71909 364994 444619
rect 366294 439954 366914 475398
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 369163 446044 369229 446045
rect 369163 445980 369164 446044
rect 369228 445980 369229 446044
rect 369163 445979 369229 445980
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 365115 304332 365181 304333
rect 365115 304268 365116 304332
rect 365180 304268 365181 304332
rect 365115 304267 365181 304268
rect 364931 71908 364997 71909
rect 364931 71844 364932 71908
rect 364996 71844 364997 71908
rect 364931 71843 364997 71844
rect 365118 3909 365178 304267
rect 365667 298756 365733 298757
rect 365667 298692 365668 298756
rect 365732 298692 365733 298756
rect 365667 298691 365733 298692
rect 365115 3908 365181 3909
rect 365115 3844 365116 3908
rect 365180 3844 365181 3908
rect 365115 3843 365181 3844
rect 365670 3501 365730 298691
rect 366294 295954 366914 331398
rect 368979 307052 369045 307053
rect 368979 306988 368980 307052
rect 369044 306988 369045 307052
rect 368979 306987 369045 306988
rect 367691 304196 367757 304197
rect 367691 304132 367692 304196
rect 367756 304132 367757 304196
rect 367691 304131 367757 304132
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 367139 286380 367205 286381
rect 367139 286316 367140 286380
rect 367204 286316 367205 286380
rect 367139 286315 367205 286316
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 364379 3500 364445 3501
rect 364379 3436 364380 3500
rect 364444 3436 364445 3500
rect 364379 3435 364445 3436
rect 365667 3500 365733 3501
rect 365667 3436 365668 3500
rect 365732 3436 365733 3500
rect 365667 3435 365733 3436
rect 363459 3364 363525 3365
rect 363459 3300 363460 3364
rect 363524 3300 363525 3364
rect 363459 3299 363525 3300
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 -1306 366914 7398
rect 367142 3501 367202 286315
rect 367323 244764 367389 244765
rect 367323 244700 367324 244764
rect 367388 244700 367389 244764
rect 367323 244699 367389 244700
rect 367326 6221 367386 244699
rect 367323 6220 367389 6221
rect 367323 6156 367324 6220
rect 367388 6156 367389 6220
rect 367323 6155 367389 6156
rect 367694 3773 367754 304131
rect 368427 254556 368493 254557
rect 368427 254492 368428 254556
rect 368492 254492 368493 254556
rect 368427 254491 368493 254492
rect 367691 3772 367757 3773
rect 367691 3708 367692 3772
rect 367756 3708 367757 3772
rect 367691 3707 367757 3708
rect 368430 3501 368490 254491
rect 368982 3637 369042 306987
rect 369166 177309 369226 445979
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 369899 269788 369965 269789
rect 369899 269724 369900 269788
rect 369964 269724 369965 269788
rect 369899 269723 369965 269724
rect 369163 177308 369229 177309
rect 369163 177244 369164 177308
rect 369228 177244 369229 177308
rect 369163 177243 369229 177244
rect 368979 3636 369045 3637
rect 368979 3572 368980 3636
rect 369044 3572 369045 3636
rect 368979 3571 369045 3572
rect 369902 3501 369962 269723
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 367139 3500 367205 3501
rect 367139 3436 367140 3500
rect 367204 3436 367205 3500
rect 367139 3435 367205 3436
rect 368427 3500 368493 3501
rect 368427 3436 368428 3500
rect 368492 3436 368493 3500
rect 368427 3435 368493 3436
rect 369899 3500 369965 3501
rect 369899 3436 369900 3500
rect 369964 3436 369965 3500
rect 369899 3435 369965 3436
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 210454 389414 245898
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 214954 393914 250398
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 96326 241718 96562 241954
rect 96646 241718 96882 241954
rect 96326 241398 96562 241634
rect 96646 241398 96882 241634
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 100826 246218 101062 246454
rect 101146 246218 101382 246454
rect 100826 245898 101062 246134
rect 101146 245898 101382 246134
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 118826 228218 119062 228454
rect 119146 228218 119382 228454
rect 118826 227898 119062 228134
rect 119146 227898 119382 228134
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 118826 120218 119062 120454
rect 119146 120218 119382 120454
rect 118826 119898 119062 120134
rect 119146 119898 119382 120134
rect 118826 84218 119062 84454
rect 119146 84218 119382 84454
rect 118826 83898 119062 84134
rect 119146 83898 119382 84134
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 123326 232718 123562 232954
rect 123646 232718 123882 232954
rect 123326 232398 123562 232634
rect 123646 232398 123882 232634
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 123326 124718 123562 124954
rect 123646 124718 123882 124954
rect 123326 124398 123562 124634
rect 123646 124398 123882 124634
rect 123326 88718 123562 88954
rect 123646 88718 123882 88954
rect 123326 88398 123562 88634
rect 123646 88398 123882 88634
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 132326 241718 132562 241954
rect 132646 241718 132882 241954
rect 132326 241398 132562 241634
rect 132646 241398 132882 241634
rect 132326 205718 132562 205954
rect 132646 205718 132882 205954
rect 132326 205398 132562 205634
rect 132646 205398 132882 205634
rect 132326 169718 132562 169954
rect 132646 169718 132882 169954
rect 132326 169398 132562 169634
rect 132646 169398 132882 169634
rect 132326 133718 132562 133954
rect 132646 133718 132882 133954
rect 132326 133398 132562 133634
rect 132646 133398 132882 133634
rect 132326 97718 132562 97954
rect 132646 97718 132882 97954
rect 132326 97398 132562 97634
rect 132646 97398 132882 97634
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 136826 246218 137062 246454
rect 137146 246218 137382 246454
rect 136826 245898 137062 246134
rect 137146 245898 137382 246134
rect 136826 210218 137062 210454
rect 137146 210218 137382 210454
rect 136826 209898 137062 210134
rect 137146 209898 137382 210134
rect 136826 174218 137062 174454
rect 137146 174218 137382 174454
rect 136826 173898 137062 174134
rect 137146 173898 137382 174134
rect 136826 138218 137062 138454
rect 137146 138218 137382 138454
rect 136826 137898 137062 138134
rect 137146 137898 137382 138134
rect 136826 102218 137062 102454
rect 137146 102218 137382 102454
rect 136826 101898 137062 102134
rect 137146 101898 137382 102134
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 141326 214718 141562 214954
rect 141646 214718 141882 214954
rect 141326 214398 141562 214634
rect 141646 214398 141882 214634
rect 141326 178718 141562 178954
rect 141646 178718 141882 178954
rect 141326 178398 141562 178634
rect 141646 178398 141882 178634
rect 141326 142718 141562 142954
rect 141646 142718 141882 142954
rect 141326 142398 141562 142634
rect 141646 142398 141882 142634
rect 141326 106718 141562 106954
rect 141646 106718 141882 106954
rect 141326 106398 141562 106634
rect 141646 106398 141882 106634
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 150326 223718 150562 223954
rect 150646 223718 150882 223954
rect 150326 223398 150562 223634
rect 150646 223398 150882 223634
rect 150326 187718 150562 187954
rect 150646 187718 150882 187954
rect 150326 187398 150562 187634
rect 150646 187398 150882 187634
rect 150326 151718 150562 151954
rect 150646 151718 150882 151954
rect 150326 151398 150562 151634
rect 150646 151398 150882 151634
rect 150326 115718 150562 115954
rect 150646 115718 150882 115954
rect 150326 115398 150562 115634
rect 150646 115398 150882 115634
rect 150326 79718 150562 79954
rect 150646 79718 150882 79954
rect 150326 79398 150562 79634
rect 150646 79398 150882 79634
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 154826 228218 155062 228454
rect 155146 228218 155382 228454
rect 154826 227898 155062 228134
rect 155146 227898 155382 228134
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 154826 156218 155062 156454
rect 155146 156218 155382 156454
rect 154826 155898 155062 156134
rect 155146 155898 155382 156134
rect 154826 120218 155062 120454
rect 155146 120218 155382 120454
rect 154826 119898 155062 120134
rect 155146 119898 155382 120134
rect 154826 84218 155062 84454
rect 155146 84218 155382 84454
rect 154826 83898 155062 84134
rect 155146 83898 155382 84134
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 159326 232718 159562 232954
rect 159646 232718 159882 232954
rect 159326 232398 159562 232634
rect 159646 232398 159882 232634
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 159326 160718 159562 160954
rect 159646 160718 159882 160954
rect 159326 160398 159562 160634
rect 159646 160398 159882 160634
rect 159326 124718 159562 124954
rect 159646 124718 159882 124954
rect 159326 124398 159562 124634
rect 159646 124398 159882 124634
rect 159326 88718 159562 88954
rect 159646 88718 159882 88954
rect 159326 88398 159562 88634
rect 159646 88398 159882 88634
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 168326 241718 168562 241954
rect 168646 241718 168882 241954
rect 168326 241398 168562 241634
rect 168646 241398 168882 241634
rect 168326 205718 168562 205954
rect 168646 205718 168882 205954
rect 168326 205398 168562 205634
rect 168646 205398 168882 205634
rect 168326 169718 168562 169954
rect 168646 169718 168882 169954
rect 168326 169398 168562 169634
rect 168646 169398 168882 169634
rect 168326 133718 168562 133954
rect 168646 133718 168882 133954
rect 168326 133398 168562 133634
rect 168646 133398 168882 133634
rect 168326 97718 168562 97954
rect 168646 97718 168882 97954
rect 168326 97398 168562 97634
rect 168646 97398 168882 97634
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 172826 246218 173062 246454
rect 173146 246218 173382 246454
rect 172826 245898 173062 246134
rect 173146 245898 173382 246134
rect 172826 210218 173062 210454
rect 173146 210218 173382 210454
rect 172826 209898 173062 210134
rect 173146 209898 173382 210134
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 172826 138218 173062 138454
rect 173146 138218 173382 138454
rect 172826 137898 173062 138134
rect 173146 137898 173382 138134
rect 172826 102218 173062 102454
rect 173146 102218 173382 102454
rect 172826 101898 173062 102134
rect 173146 101898 173382 102134
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 177326 214718 177562 214954
rect 177646 214718 177882 214954
rect 177326 214398 177562 214634
rect 177646 214398 177882 214634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 177326 106718 177562 106954
rect 177646 106718 177882 106954
rect 177326 106398 177562 106634
rect 177646 106398 177882 106634
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 190826 228218 191062 228454
rect 191146 228218 191382 228454
rect 190826 227898 191062 228134
rect 191146 227898 191382 228134
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 204326 241718 204562 241954
rect 204646 241718 204882 241954
rect 204326 241398 204562 241634
rect 204646 241398 204882 241634
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 220328 547718 220564 547954
rect 220328 547398 220564 547634
rect 356056 547718 356292 547954
rect 356056 547398 356292 547634
rect 221008 543218 221244 543454
rect 221008 542898 221244 543134
rect 355376 543218 355612 543454
rect 355376 542898 355612 543134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 220328 511718 220564 511954
rect 220328 511398 220564 511634
rect 356056 511718 356292 511954
rect 356056 511398 356292 511634
rect 221008 507218 221244 507454
rect 221008 506898 221244 507134
rect 355376 507218 355612 507454
rect 355376 506898 355612 507134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 208826 246218 209062 246454
rect 209146 246218 209382 246454
rect 208826 245898 209062 246134
rect 209146 245898 209382 246134
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 252010 439718 252246 439954
rect 252010 439398 252246 439634
rect 282730 439718 282966 439954
rect 282730 439398 282966 439634
rect 313450 439718 313686 439954
rect 313450 439398 313686 439634
rect 344170 439718 344406 439954
rect 344170 439398 344406 439634
rect 236650 435218 236886 435454
rect 236650 434898 236886 435134
rect 267370 435218 267606 435454
rect 267370 434898 267606 435134
rect 298090 435218 298326 435454
rect 298090 434898 298326 435134
rect 328810 435218 329046 435454
rect 328810 434898 329046 435134
rect 359530 435218 359766 435454
rect 359530 434898 359766 435134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 252010 403718 252246 403954
rect 252010 403398 252246 403634
rect 282730 403718 282966 403954
rect 282730 403398 282966 403634
rect 313450 403718 313686 403954
rect 313450 403398 313686 403634
rect 344170 403718 344406 403954
rect 344170 403398 344406 403634
rect 236650 399218 236886 399454
rect 236650 398898 236886 399134
rect 267370 399218 267606 399454
rect 267370 398898 267606 399134
rect 298090 399218 298326 399454
rect 298090 398898 298326 399134
rect 328810 399218 329046 399454
rect 328810 398898 329046 399134
rect 359530 399218 359766 399454
rect 359530 398898 359766 399134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 252010 367718 252246 367954
rect 252010 367398 252246 367634
rect 282730 367718 282966 367954
rect 282730 367398 282966 367634
rect 313450 367718 313686 367954
rect 313450 367398 313686 367634
rect 344170 367718 344406 367954
rect 344170 367398 344406 367634
rect 236650 363218 236886 363454
rect 236650 362898 236886 363134
rect 267370 363218 267606 363454
rect 267370 362898 267606 363134
rect 298090 363218 298326 363454
rect 298090 362898 298326 363134
rect 328810 363218 329046 363454
rect 328810 362898 329046 363134
rect 359530 363218 359766 363454
rect 359530 362898 359766 363134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 252010 331718 252246 331954
rect 252010 331398 252246 331634
rect 282730 331718 282966 331954
rect 282730 331398 282966 331634
rect 313450 331718 313686 331954
rect 313450 331398 313686 331634
rect 344170 331718 344406 331954
rect 344170 331398 344406 331634
rect 236650 327218 236886 327454
rect 236650 326898 236886 327134
rect 267370 327218 267606 327454
rect 267370 326898 267606 327134
rect 298090 327218 298326 327454
rect 298090 326898 298326 327134
rect 328810 327218 329046 327454
rect 328810 326898 329046 327134
rect 359530 327218 359766 327454
rect 359530 326898 359766 327134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 244826 246218 245062 246454
rect 245146 246218 245382 246454
rect 244826 245898 245062 246134
rect 245146 245898 245382 246134
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 280826 246218 281062 246454
rect 281146 246218 281382 246454
rect 280826 245898 281062 246134
rect 281146 245898 281382 246134
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 316826 246218 317062 246454
rect 317146 246218 317382 246454
rect 316826 245898 317062 246134
rect 317146 245898 317382 246134
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 220328 223718 220564 223954
rect 220328 223398 220564 223634
rect 356056 223718 356292 223954
rect 356056 223398 356292 223634
rect 221008 219218 221244 219454
rect 221008 218898 221244 219134
rect 355376 219218 355612 219454
rect 355376 218898 355612 219134
rect 220328 187718 220564 187954
rect 220328 187398 220564 187634
rect 356056 187718 356292 187954
rect 356056 187398 356292 187634
rect 221008 183218 221244 183454
rect 221008 182898 221244 183134
rect 355376 183218 355612 183454
rect 355376 182898 355612 183134
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 220328 547954
rect 220564 547718 356056 547954
rect 356292 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 220328 547634
rect 220564 547398 356056 547634
rect 356292 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 221008 543454
rect 221244 543218 355376 543454
rect 355612 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 221008 543134
rect 221244 542898 355376 543134
rect 355612 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 220328 511954
rect 220564 511718 356056 511954
rect 356292 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 220328 511634
rect 220564 511398 356056 511634
rect 356292 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 221008 507454
rect 221244 507218 355376 507454
rect 355612 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 221008 507134
rect 221244 506898 355376 507134
rect 355612 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 252010 439954
rect 252246 439718 282730 439954
rect 282966 439718 313450 439954
rect 313686 439718 344170 439954
rect 344406 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 252010 439634
rect 252246 439398 282730 439634
rect 282966 439398 313450 439634
rect 313686 439398 344170 439634
rect 344406 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 236650 435454
rect 236886 435218 267370 435454
rect 267606 435218 298090 435454
rect 298326 435218 328810 435454
rect 329046 435218 359530 435454
rect 359766 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 236650 435134
rect 236886 434898 267370 435134
rect 267606 434898 298090 435134
rect 298326 434898 328810 435134
rect 329046 434898 359530 435134
rect 359766 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 252010 403954
rect 252246 403718 282730 403954
rect 282966 403718 313450 403954
rect 313686 403718 344170 403954
rect 344406 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 252010 403634
rect 252246 403398 282730 403634
rect 282966 403398 313450 403634
rect 313686 403398 344170 403634
rect 344406 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 236650 399454
rect 236886 399218 267370 399454
rect 267606 399218 298090 399454
rect 298326 399218 328810 399454
rect 329046 399218 359530 399454
rect 359766 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 236650 399134
rect 236886 398898 267370 399134
rect 267606 398898 298090 399134
rect 298326 398898 328810 399134
rect 329046 398898 359530 399134
rect 359766 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 252010 367954
rect 252246 367718 282730 367954
rect 282966 367718 313450 367954
rect 313686 367718 344170 367954
rect 344406 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 252010 367634
rect 252246 367398 282730 367634
rect 282966 367398 313450 367634
rect 313686 367398 344170 367634
rect 344406 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 236650 363454
rect 236886 363218 267370 363454
rect 267606 363218 298090 363454
rect 298326 363218 328810 363454
rect 329046 363218 359530 363454
rect 359766 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 236650 363134
rect 236886 362898 267370 363134
rect 267606 362898 298090 363134
rect 298326 362898 328810 363134
rect 329046 362898 359530 363134
rect 359766 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 252010 331954
rect 252246 331718 282730 331954
rect 282966 331718 313450 331954
rect 313686 331718 344170 331954
rect 344406 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 252010 331634
rect 252246 331398 282730 331634
rect 282966 331398 313450 331634
rect 313686 331398 344170 331634
rect 344406 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 236650 327454
rect 236886 327218 267370 327454
rect 267606 327218 298090 327454
rect 298326 327218 328810 327454
rect 329046 327218 359530 327454
rect 359766 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 236650 327134
rect 236886 326898 267370 327134
rect 267606 326898 298090 327134
rect 298326 326898 328810 327134
rect 329046 326898 359530 327134
rect 359766 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 220328 223954
rect 220564 223718 356056 223954
rect 356292 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 220328 223634
rect 220564 223398 356056 223634
rect 356292 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 221008 219454
rect 221244 219218 355376 219454
rect 355612 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 221008 219134
rect 221244 218898 355376 219134
rect 355612 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 220328 187954
rect 220564 187718 356056 187954
rect 356292 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 220328 187634
rect 220564 187398 356056 187634
rect 356292 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 221008 183454
rect 221244 183218 355376 183454
rect 355612 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 221008 183134
rect 221244 182898 355376 183134
rect 355612 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 123326 124954
rect 123562 124718 123646 124954
rect 123882 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 123326 124634
rect 123562 124398 123646 124634
rect 123882 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sky130_sram_2kbyte_1rw1r_32x512_8  dram_inst
timestamp 0
transform 1 0 220000 0 1 480000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  iram_inst
timestamp 0
transform 1 0 220000 0 1 160000
box 0 0 136620 83308
use rvj1_caravel_soc  rvj1_soc
timestamp 0
transform 1 0 232400 0 1 310400
box 14 0 131362 133626
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 1794 -7654 2414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 37794 -7654 38414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 73794 -7654 74414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 109794 -7654 110414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 145794 -7654 146414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 181794 -7654 182414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 217794 -7654 218414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 217794 245308 218414 478000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 217794 565308 218414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 253794 -7654 254414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 253794 245308 254414 308400 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 253794 565308 254414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 289794 -7654 290414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 289794 245308 290414 308400 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 289794 565308 290414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 -7654 326414 158000 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 245308 326414 308400 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 565308 326414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 361794 -7654 362414 308400 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 361794 446026 362414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 397794 -7654 398414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 433794 -7654 434414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 469794 -7654 470414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 505794 -7654 506414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 541794 -7654 542414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 577794 -7654 578414 711590 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 2866 592650 3486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 38866 592650 39486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 74866 592650 75486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 110866 592650 111486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 146866 592650 147486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 182866 592650 183486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 218866 592650 219486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 254866 592650 255486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 290866 592650 291486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 326866 592650 327486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 362866 592650 363486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 398866 592650 399486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 434866 592650 435486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 470866 592650 471486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 506866 592650 507486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 542866 592650 543486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 578866 592650 579486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 614866 592650 615486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 650866 592650 651486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -8726 686866 592650 687486 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 10794 -7654 11414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 46794 -7654 47414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 82794 -7654 83414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 118794 -7654 119414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 154794 -7654 155414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 190794 -7654 191414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 226794 -7654 227414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 226794 245308 227414 478000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 226794 565308 227414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 262794 -7654 263414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 262794 245308 263414 308400 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 262794 565308 263414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 298794 -7654 299414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 298794 245308 299414 308400 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 298794 565308 299414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 334794 -7654 335414 158000 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 334794 245308 335414 308400 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 334794 565308 335414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 370794 -7654 371414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 406794 -7654 407414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 442794 -7654 443414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 478794 -7654 479414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 514794 -7654 515414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 550794 -7654 551414 711590 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 11866 592650 12486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 47866 592650 48486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 83866 592650 84486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 119866 592650 120486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 155866 592650 156486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 191866 592650 192486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 227866 592650 228486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 263866 592650 264486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 299866 592650 300486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 335866 592650 336486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 371866 592650 372486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 407866 592650 408486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 443866 592650 444486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 479866 592650 480486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 515866 592650 516486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 551866 592650 552486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 587866 592650 588486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 623866 592650 624486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 659866 592650 660486 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8726 695866 592650 696486 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 19794 -7654 20414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 55794 -7654 56414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 91794 -7654 92414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 127794 -7654 128414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 163794 -7654 164414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 199794 -7654 200414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 235794 -7654 236414 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 235794 565308 236414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 271794 -7654 272414 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 271794 565308 272414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 307794 -7654 308414 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 307794 565308 308414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 343794 -7654 344414 158000 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 343794 565308 344414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 379794 -7654 380414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 415794 -7654 416414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 451794 -7654 452414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 487794 -7654 488414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 523794 -7654 524414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 559794 -7654 560414 711590 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 20866 592650 21486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 56866 592650 57486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 92866 592650 93486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 128866 592650 129486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 164866 592650 165486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 200866 592650 201486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 236866 592650 237486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 272866 592650 273486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 308866 592650 309486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 344866 592650 345486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 380866 592650 381486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 416866 592650 417486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 452866 592650 453486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 488866 592650 489486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 524866 592650 525486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 560866 592650 561486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 596866 592650 597486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 632866 592650 633486 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -8726 668866 592650 669486 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 28794 -7654 29414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 64794 -7654 65414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 100794 -7654 101414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 136794 -7654 137414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 172794 -7654 173414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 208794 -7654 209414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 244794 -7654 245414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 244794 245308 245414 308400 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 244794 565308 245414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 280794 -7654 281414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 280794 245308 281414 308400 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 280794 565308 281414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 316794 -7654 317414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 316794 245308 317414 308400 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 316794 565308 317414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 352794 -7654 353414 158000 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 352794 245308 353414 308400 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 352794 565308 353414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 388794 -7654 389414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 424794 -7654 425414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 460794 -7654 461414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 496794 -7654 497414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 532794 -7654 533414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 568794 -7654 569414 711590 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 29866 592650 30486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 65866 592650 66486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 101866 592650 102486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 137866 592650 138486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 173866 592650 174486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 209866 592650 210486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 245866 592650 246486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 281866 592650 282486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 317866 592650 318486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 353866 592650 354486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 389866 592650 390486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 425866 592650 426486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 461866 592650 462486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 497866 592650 498486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 533866 592650 534486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 569866 592650 570486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 605866 592650 606486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 641866 592650 642486 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -8726 677866 592650 678486 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 24294 -7654 24914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 60294 -7654 60914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 96294 -7654 96914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 132294 -7654 132914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 168294 -7654 168914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 204294 -7654 204914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 240294 -7654 240914 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 240294 565308 240914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 276294 -7654 276914 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 276294 565308 276914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 312294 -7654 312914 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 312294 565308 312914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 348294 -7654 348914 158000 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 348294 565308 348914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 384294 -7654 384914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 420294 -7654 420914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 456294 -7654 456914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 492294 -7654 492914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 528294 -7654 528914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 564294 -7654 564914 711590 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 25366 592650 25986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 61366 592650 61986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 97366 592650 97986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 133366 592650 133986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 169366 592650 169986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 205366 592650 205986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 241366 592650 241986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 277366 592650 277986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 313366 592650 313986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 349366 592650 349986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 385366 592650 385986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 421366 592650 421986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 457366 592650 457986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 493366 592650 493986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 529366 592650 529986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 565366 592650 565986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 601366 592650 601986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 637366 592650 637986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -8726 673366 592650 673986 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 33294 -7654 33914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 69294 -7654 69914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 105294 -7654 105914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 141294 -7654 141914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 177294 -7654 177914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 213294 -7654 213914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 249294 -7654 249914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 249294 245308 249914 308400 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 249294 565308 249914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 285294 -7654 285914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 285294 245308 285914 308400 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 285294 565308 285914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 321294 -7654 321914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 321294 245308 321914 308400 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 321294 565308 321914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 357294 -7654 357914 158000 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 357294 245308 357914 308400 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 357294 565308 357914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 393294 -7654 393914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 429294 -7654 429914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 465294 -7654 465914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 501294 -7654 501914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 537294 -7654 537914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 573294 -7654 573914 711590 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 34366 592650 34986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 70366 592650 70986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 106366 592650 106986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 142366 592650 142986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 178366 592650 178986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 214366 592650 214986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 250366 592650 250986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 286366 592650 286986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 322366 592650 322986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 358366 592650 358986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 394366 592650 394986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 430366 592650 430986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 466366 592650 466986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 502366 592650 502986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 538366 592650 538986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 574366 592650 574986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 610366 592650 610986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 646366 592650 646986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -8726 682366 592650 682986 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 6294 -7654 6914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 42294 -7654 42914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 78294 -7654 78914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 114294 -7654 114914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 150294 -7654 150914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 186294 -7654 186914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 222294 -7654 222914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 222294 245308 222914 478000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 222294 565308 222914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 258294 -7654 258914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 258294 245308 258914 308400 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 258294 565308 258914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 294294 -7654 294914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 294294 245308 294914 308400 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 294294 565308 294914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 330294 -7654 330914 158000 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 330294 245308 330914 308400 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 330294 565308 330914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 366294 -7654 366914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 402294 -7654 402914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 438294 -7654 438914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 474294 -7654 474914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 510294 -7654 510914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 546294 -7654 546914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 582294 -7654 582914 711590 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 7366 592650 7986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 43366 592650 43986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 79366 592650 79986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 115366 592650 115986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 151366 592650 151986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 187366 592650 187986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 223366 592650 223986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 259366 592650 259986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 295366 592650 295986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 331366 592650 331986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 367366 592650 367986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 403366 592650 403986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 439366 592650 439986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 475366 592650 475986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 511366 592650 511986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 547366 592650 547986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 583366 592650 583986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 619366 592650 619986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 655366 592650 655986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -8726 691366 592650 691986 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 15294 -7654 15914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 51294 -7654 51914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 87294 -7654 87914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 123294 -7654 123914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 159294 -7654 159914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 195294 -7654 195914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 231294 -7654 231914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 231294 245308 231914 308400 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 231294 565308 231914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 267294 -7654 267914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 267294 245308 267914 308400 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 267294 565308 267914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 303294 -7654 303914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 303294 245308 303914 308400 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 303294 565308 303914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 339294 -7654 339914 158000 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 339294 245308 339914 308400 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 339294 565308 339914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 375294 -7654 375914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 411294 -7654 411914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 447294 -7654 447914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 483294 -7654 483914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 519294 -7654 519914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 555294 -7654 555914 711590 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 16366 592650 16986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 52366 592650 52986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 88366 592650 88986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 124366 592650 124986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 160366 592650 160986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 196366 592650 196986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 232366 592650 232986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 268366 592650 268986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 304366 592650 304986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 340366 592650 340986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 376366 592650 376986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 412366 592650 412986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 448366 592650 448986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 484366 592650 484986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 520366 592650 520986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 556366 592650 556986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 592366 592650 592986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 628366 592650 628986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 664366 592650 664986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -8726 700366 592650 700986 6 vssd2
port 538 nsew ground bidirectional
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
